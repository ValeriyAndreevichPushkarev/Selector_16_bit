module address_decode_2
(

    input wire[1:0] addr_src,

    output wire[3:0] addr_positional
);



assign addr_positional[3] = (addr_src==2'b11) ?1'b1:1'b0;

assign addr_positional[2] = (addr_src==2'b10) ?1'b1:1'b0;

assign addr_positional[1] = (addr_src==2'b01) ?1'b1:1'b0;

assign addr_positional[0] = (addr_src==2'b00) ?1'b1:1'b0;



endmodule

module address_decode_14
(

    input wire[13:0] addr_src,

    output wire[27:0] addr_positional
);



address_decode_2 enc0(addr_src[1:0], addr_positional[27:24]);

address_decode_2 enc1(addr_src[3:2], addr_positional[23:20]);

address_decode_2 enc2(addr_src[5:4], addr_positional[19:16]);

address_decode_2 enc3(addr_src[7:6], addr_positional[15:12]);

address_decode_2 enc4(addr_src[9:8], addr_positional[11:8]);

address_decode_2 enc5(addr_src[11:10], addr_positional[7:4]);

address_decode_2 enc6(addr_src[13:12], addr_positional[3:0]);



endmodule

module Selector_2
(

    input wire selector_enabled,

    input wire[27:0] addr_src,

    output wire[3:0] addr_positional,

    output wire[27:0] addr_remain
);




assign addr_remain =        (selector_enabled==1'b1)? {4'b0,addr_src[27:4]}:28'b0;
assign addr_positional =    (selector_enabled==1'b1)? addr_src[3:0] : 4'b0;

endmodule



module Selector_14
(

    input wire[13:0] addr,

    output wire[16383:0] addr_positional
);





 

   wire[27:0] addr_src;

   address_decode_14 sel_1 (addr, addr_src);wire[3:0] wires_0_0;

wire[27:0] addr_0_0;

Selector_2 s0_0(1'b1, addr_src, wires_0_0, addr_0_0);

wire[3:0] wires_0_1;

wire[27:0] addr_0_1;

Selector_2 s0_1(wires_0_0[0], addr_0_0, wires_0_1,addr_0_1);

wire[3:0] wires_1_1;

wire[27:0] addr_1_1;

Selector_2 s1_1(wires_0_0[1], addr_0_0, wires_1_1,addr_1_1);

wire[3:0] wires_2_1;

wire[27:0] addr_2_1;

Selector_2 s2_1(wires_0_0[2], addr_0_0, wires_2_1,addr_2_1);

wire[3:0] wires_3_1;

wire[27:0] addr_3_1;

Selector_2 s3_1(wires_0_0[3], addr_0_0, wires_3_1,addr_3_1);

wire[3:0] wires_0_2;

wire[27:0] addr_0_2;

Selector_2 s0_2(wires_0_1[0], addr_0_1, wires_0_2,addr_0_2);

wire[3:0] wires_1_2;

wire[27:0] addr_1_2;

Selector_2 s1_2(wires_0_1[1], addr_0_1, wires_1_2,addr_1_2);

wire[3:0] wires_2_2;

wire[27:0] addr_2_2;

Selector_2 s2_2(wires_0_1[2], addr_0_1, wires_2_2,addr_2_2);

wire[3:0] wires_3_2;

wire[27:0] addr_3_2;

Selector_2 s3_2(wires_0_1[3], addr_0_1, wires_3_2,addr_3_2);

wire[3:0] wires_4_2;

wire[27:0] addr_4_2;

Selector_2 s4_2(wires_1_1[0], addr_1_1, wires_4_2,addr_4_2);

wire[3:0] wires_5_2;

wire[27:0] addr_5_2;

Selector_2 s5_2(wires_1_1[1], addr_1_1, wires_5_2,addr_5_2);

wire[3:0] wires_6_2;

wire[27:0] addr_6_2;

Selector_2 s6_2(wires_1_1[2], addr_1_1, wires_6_2,addr_6_2);

wire[3:0] wires_7_2;

wire[27:0] addr_7_2;

Selector_2 s7_2(wires_1_1[3], addr_1_1, wires_7_2,addr_7_2);

wire[3:0] wires_8_2;

wire[27:0] addr_8_2;

Selector_2 s8_2(wires_2_1[0], addr_2_1, wires_8_2,addr_8_2);

wire[3:0] wires_9_2;

wire[27:0] addr_9_2;

Selector_2 s9_2(wires_2_1[1], addr_2_1, wires_9_2,addr_9_2);

wire[3:0] wires_10_2;

wire[27:0] addr_10_2;

Selector_2 s10_2(wires_2_1[2], addr_2_1, wires_10_2,addr_10_2);

wire[3:0] wires_11_2;

wire[27:0] addr_11_2;

Selector_2 s11_2(wires_2_1[3], addr_2_1, wires_11_2,addr_11_2);

wire[3:0] wires_12_2;

wire[27:0] addr_12_2;

Selector_2 s12_2(wires_3_1[0], addr_3_1, wires_12_2,addr_12_2);

wire[3:0] wires_13_2;

wire[27:0] addr_13_2;

Selector_2 s13_2(wires_3_1[1], addr_3_1, wires_13_2,addr_13_2);

wire[3:0] wires_14_2;

wire[27:0] addr_14_2;

Selector_2 s14_2(wires_3_1[2], addr_3_1, wires_14_2,addr_14_2);

wire[3:0] wires_15_2;

wire[27:0] addr_15_2;

Selector_2 s15_2(wires_3_1[3], addr_3_1, wires_15_2,addr_15_2);

wire[3:0] wires_0_3;

wire[27:0] addr_0_3;

Selector_2 s0_3(wires_0_2[0], addr_0_2, wires_0_3,addr_0_3);

wire[3:0] wires_1_3;

wire[27:0] addr_1_3;

Selector_2 s1_3(wires_0_2[1], addr_0_2, wires_1_3,addr_1_3);

wire[3:0] wires_2_3;

wire[27:0] addr_2_3;

Selector_2 s2_3(wires_0_2[2], addr_0_2, wires_2_3,addr_2_3);

wire[3:0] wires_3_3;

wire[27:0] addr_3_3;

Selector_2 s3_3(wires_0_2[3], addr_0_2, wires_3_3,addr_3_3);

wire[3:0] wires_4_3;

wire[27:0] addr_4_3;

Selector_2 s4_3(wires_1_2[0], addr_1_2, wires_4_3,addr_4_3);

wire[3:0] wires_5_3;

wire[27:0] addr_5_3;

Selector_2 s5_3(wires_1_2[1], addr_1_2, wires_5_3,addr_5_3);

wire[3:0] wires_6_3;

wire[27:0] addr_6_3;

Selector_2 s6_3(wires_1_2[2], addr_1_2, wires_6_3,addr_6_3);

wire[3:0] wires_7_3;

wire[27:0] addr_7_3;

Selector_2 s7_3(wires_1_2[3], addr_1_2, wires_7_3,addr_7_3);

wire[3:0] wires_8_3;

wire[27:0] addr_8_3;

Selector_2 s8_3(wires_2_2[0], addr_2_2, wires_8_3,addr_8_3);

wire[3:0] wires_9_3;

wire[27:0] addr_9_3;

Selector_2 s9_3(wires_2_2[1], addr_2_2, wires_9_3,addr_9_3);

wire[3:0] wires_10_3;

wire[27:0] addr_10_3;

Selector_2 s10_3(wires_2_2[2], addr_2_2, wires_10_3,addr_10_3);

wire[3:0] wires_11_3;

wire[27:0] addr_11_3;

Selector_2 s11_3(wires_2_2[3], addr_2_2, wires_11_3,addr_11_3);

wire[3:0] wires_12_3;

wire[27:0] addr_12_3;

Selector_2 s12_3(wires_3_2[0], addr_3_2, wires_12_3,addr_12_3);

wire[3:0] wires_13_3;

wire[27:0] addr_13_3;

Selector_2 s13_3(wires_3_2[1], addr_3_2, wires_13_3,addr_13_3);

wire[3:0] wires_14_3;

wire[27:0] addr_14_3;

Selector_2 s14_3(wires_3_2[2], addr_3_2, wires_14_3,addr_14_3);

wire[3:0] wires_15_3;

wire[27:0] addr_15_3;

Selector_2 s15_3(wires_3_2[3], addr_3_2, wires_15_3,addr_15_3);

wire[3:0] wires_16_3;

wire[27:0] addr_16_3;

Selector_2 s16_3(wires_4_2[0], addr_4_2, wires_16_3,addr_16_3);

wire[3:0] wires_17_3;

wire[27:0] addr_17_3;

Selector_2 s17_3(wires_4_2[1], addr_4_2, wires_17_3,addr_17_3);

wire[3:0] wires_18_3;

wire[27:0] addr_18_3;

Selector_2 s18_3(wires_4_2[2], addr_4_2, wires_18_3,addr_18_3);

wire[3:0] wires_19_3;

wire[27:0] addr_19_3;

Selector_2 s19_3(wires_4_2[3], addr_4_2, wires_19_3,addr_19_3);

wire[3:0] wires_20_3;

wire[27:0] addr_20_3;

Selector_2 s20_3(wires_5_2[0], addr_5_2, wires_20_3,addr_20_3);

wire[3:0] wires_21_3;

wire[27:0] addr_21_3;

Selector_2 s21_3(wires_5_2[1], addr_5_2, wires_21_3,addr_21_3);

wire[3:0] wires_22_3;

wire[27:0] addr_22_3;

Selector_2 s22_3(wires_5_2[2], addr_5_2, wires_22_3,addr_22_3);

wire[3:0] wires_23_3;

wire[27:0] addr_23_3;

Selector_2 s23_3(wires_5_2[3], addr_5_2, wires_23_3,addr_23_3);

wire[3:0] wires_24_3;

wire[27:0] addr_24_3;

Selector_2 s24_3(wires_6_2[0], addr_6_2, wires_24_3,addr_24_3);

wire[3:0] wires_25_3;

wire[27:0] addr_25_3;

Selector_2 s25_3(wires_6_2[1], addr_6_2, wires_25_3,addr_25_3);

wire[3:0] wires_26_3;

wire[27:0] addr_26_3;

Selector_2 s26_3(wires_6_2[2], addr_6_2, wires_26_3,addr_26_3);

wire[3:0] wires_27_3;

wire[27:0] addr_27_3;

Selector_2 s27_3(wires_6_2[3], addr_6_2, wires_27_3,addr_27_3);

wire[3:0] wires_28_3;

wire[27:0] addr_28_3;

Selector_2 s28_3(wires_7_2[0], addr_7_2, wires_28_3,addr_28_3);

wire[3:0] wires_29_3;

wire[27:0] addr_29_3;

Selector_2 s29_3(wires_7_2[1], addr_7_2, wires_29_3,addr_29_3);

wire[3:0] wires_30_3;

wire[27:0] addr_30_3;

Selector_2 s30_3(wires_7_2[2], addr_7_2, wires_30_3,addr_30_3);

wire[3:0] wires_31_3;

wire[27:0] addr_31_3;

Selector_2 s31_3(wires_7_2[3], addr_7_2, wires_31_3,addr_31_3);

wire[3:0] wires_32_3;

wire[27:0] addr_32_3;

Selector_2 s32_3(wires_8_2[0], addr_8_2, wires_32_3,addr_32_3);

wire[3:0] wires_33_3;

wire[27:0] addr_33_3;

Selector_2 s33_3(wires_8_2[1], addr_8_2, wires_33_3,addr_33_3);

wire[3:0] wires_34_3;

wire[27:0] addr_34_3;

Selector_2 s34_3(wires_8_2[2], addr_8_2, wires_34_3,addr_34_3);

wire[3:0] wires_35_3;

wire[27:0] addr_35_3;

Selector_2 s35_3(wires_8_2[3], addr_8_2, wires_35_3,addr_35_3);

wire[3:0] wires_36_3;

wire[27:0] addr_36_3;

Selector_2 s36_3(wires_9_2[0], addr_9_2, wires_36_3,addr_36_3);

wire[3:0] wires_37_3;

wire[27:0] addr_37_3;

Selector_2 s37_3(wires_9_2[1], addr_9_2, wires_37_3,addr_37_3);

wire[3:0] wires_38_3;

wire[27:0] addr_38_3;

Selector_2 s38_3(wires_9_2[2], addr_9_2, wires_38_3,addr_38_3);

wire[3:0] wires_39_3;

wire[27:0] addr_39_3;

Selector_2 s39_3(wires_9_2[3], addr_9_2, wires_39_3,addr_39_3);

wire[3:0] wires_40_3;

wire[27:0] addr_40_3;

Selector_2 s40_3(wires_10_2[0], addr_10_2, wires_40_3,addr_40_3);

wire[3:0] wires_41_3;

wire[27:0] addr_41_3;

Selector_2 s41_3(wires_10_2[1], addr_10_2, wires_41_3,addr_41_3);

wire[3:0] wires_42_3;

wire[27:0] addr_42_3;

Selector_2 s42_3(wires_10_2[2], addr_10_2, wires_42_3,addr_42_3);

wire[3:0] wires_43_3;

wire[27:0] addr_43_3;

Selector_2 s43_3(wires_10_2[3], addr_10_2, wires_43_3,addr_43_3);

wire[3:0] wires_44_3;

wire[27:0] addr_44_3;

Selector_2 s44_3(wires_11_2[0], addr_11_2, wires_44_3,addr_44_3);

wire[3:0] wires_45_3;

wire[27:0] addr_45_3;

Selector_2 s45_3(wires_11_2[1], addr_11_2, wires_45_3,addr_45_3);

wire[3:0] wires_46_3;

wire[27:0] addr_46_3;

Selector_2 s46_3(wires_11_2[2], addr_11_2, wires_46_3,addr_46_3);

wire[3:0] wires_47_3;

wire[27:0] addr_47_3;

Selector_2 s47_3(wires_11_2[3], addr_11_2, wires_47_3,addr_47_3);

wire[3:0] wires_48_3;

wire[27:0] addr_48_3;

Selector_2 s48_3(wires_12_2[0], addr_12_2, wires_48_3,addr_48_3);

wire[3:0] wires_49_3;

wire[27:0] addr_49_3;

Selector_2 s49_3(wires_12_2[1], addr_12_2, wires_49_3,addr_49_3);

wire[3:0] wires_50_3;

wire[27:0] addr_50_3;

Selector_2 s50_3(wires_12_2[2], addr_12_2, wires_50_3,addr_50_3);

wire[3:0] wires_51_3;

wire[27:0] addr_51_3;

Selector_2 s51_3(wires_12_2[3], addr_12_2, wires_51_3,addr_51_3);

wire[3:0] wires_52_3;

wire[27:0] addr_52_3;

Selector_2 s52_3(wires_13_2[0], addr_13_2, wires_52_3,addr_52_3);

wire[3:0] wires_53_3;

wire[27:0] addr_53_3;

Selector_2 s53_3(wires_13_2[1], addr_13_2, wires_53_3,addr_53_3);

wire[3:0] wires_54_3;

wire[27:0] addr_54_3;

Selector_2 s54_3(wires_13_2[2], addr_13_2, wires_54_3,addr_54_3);

wire[3:0] wires_55_3;

wire[27:0] addr_55_3;

Selector_2 s55_3(wires_13_2[3], addr_13_2, wires_55_3,addr_55_3);

wire[3:0] wires_56_3;

wire[27:0] addr_56_3;

Selector_2 s56_3(wires_14_2[0], addr_14_2, wires_56_3,addr_56_3);

wire[3:0] wires_57_3;

wire[27:0] addr_57_3;

Selector_2 s57_3(wires_14_2[1], addr_14_2, wires_57_3,addr_57_3);

wire[3:0] wires_58_3;

wire[27:0] addr_58_3;

Selector_2 s58_3(wires_14_2[2], addr_14_2, wires_58_3,addr_58_3);

wire[3:0] wires_59_3;

wire[27:0] addr_59_3;

Selector_2 s59_3(wires_14_2[3], addr_14_2, wires_59_3,addr_59_3);

wire[3:0] wires_60_3;

wire[27:0] addr_60_3;

Selector_2 s60_3(wires_15_2[0], addr_15_2, wires_60_3,addr_60_3);

wire[3:0] wires_61_3;

wire[27:0] addr_61_3;

Selector_2 s61_3(wires_15_2[1], addr_15_2, wires_61_3,addr_61_3);

wire[3:0] wires_62_3;

wire[27:0] addr_62_3;

Selector_2 s62_3(wires_15_2[2], addr_15_2, wires_62_3,addr_62_3);

wire[3:0] wires_63_3;

wire[27:0] addr_63_3;

Selector_2 s63_3(wires_15_2[3], addr_15_2, wires_63_3,addr_63_3);

wire[3:0] wires_0_4;

wire[27:0] addr_0_4;

Selector_2 s0_4(wires_0_3[0], addr_0_3, wires_0_4,addr_0_4);

wire[3:0] wires_1_4;

wire[27:0] addr_1_4;

Selector_2 s1_4(wires_0_3[1], addr_0_3, wires_1_4,addr_1_4);

wire[3:0] wires_2_4;

wire[27:0] addr_2_4;

Selector_2 s2_4(wires_0_3[2], addr_0_3, wires_2_4,addr_2_4);

wire[3:0] wires_3_4;

wire[27:0] addr_3_4;

Selector_2 s3_4(wires_0_3[3], addr_0_3, wires_3_4,addr_3_4);

wire[3:0] wires_4_4;

wire[27:0] addr_4_4;

Selector_2 s4_4(wires_1_3[0], addr_1_3, wires_4_4,addr_4_4);

wire[3:0] wires_5_4;

wire[27:0] addr_5_4;

Selector_2 s5_4(wires_1_3[1], addr_1_3, wires_5_4,addr_5_4);

wire[3:0] wires_6_4;

wire[27:0] addr_6_4;

Selector_2 s6_4(wires_1_3[2], addr_1_3, wires_6_4,addr_6_4);

wire[3:0] wires_7_4;

wire[27:0] addr_7_4;

Selector_2 s7_4(wires_1_3[3], addr_1_3, wires_7_4,addr_7_4);

wire[3:0] wires_8_4;

wire[27:0] addr_8_4;

Selector_2 s8_4(wires_2_3[0], addr_2_3, wires_8_4,addr_8_4);

wire[3:0] wires_9_4;

wire[27:0] addr_9_4;

Selector_2 s9_4(wires_2_3[1], addr_2_3, wires_9_4,addr_9_4);

wire[3:0] wires_10_4;

wire[27:0] addr_10_4;

Selector_2 s10_4(wires_2_3[2], addr_2_3, wires_10_4,addr_10_4);

wire[3:0] wires_11_4;

wire[27:0] addr_11_4;

Selector_2 s11_4(wires_2_3[3], addr_2_3, wires_11_4,addr_11_4);

wire[3:0] wires_12_4;

wire[27:0] addr_12_4;

Selector_2 s12_4(wires_3_3[0], addr_3_3, wires_12_4,addr_12_4);

wire[3:0] wires_13_4;

wire[27:0] addr_13_4;

Selector_2 s13_4(wires_3_3[1], addr_3_3, wires_13_4,addr_13_4);

wire[3:0] wires_14_4;

wire[27:0] addr_14_4;

Selector_2 s14_4(wires_3_3[2], addr_3_3, wires_14_4,addr_14_4);

wire[3:0] wires_15_4;

wire[27:0] addr_15_4;

Selector_2 s15_4(wires_3_3[3], addr_3_3, wires_15_4,addr_15_4);

wire[3:0] wires_16_4;

wire[27:0] addr_16_4;

Selector_2 s16_4(wires_4_3[0], addr_4_3, wires_16_4,addr_16_4);

wire[3:0] wires_17_4;

wire[27:0] addr_17_4;

Selector_2 s17_4(wires_4_3[1], addr_4_3, wires_17_4,addr_17_4);

wire[3:0] wires_18_4;

wire[27:0] addr_18_4;

Selector_2 s18_4(wires_4_3[2], addr_4_3, wires_18_4,addr_18_4);

wire[3:0] wires_19_4;

wire[27:0] addr_19_4;

Selector_2 s19_4(wires_4_3[3], addr_4_3, wires_19_4,addr_19_4);

wire[3:0] wires_20_4;

wire[27:0] addr_20_4;

Selector_2 s20_4(wires_5_3[0], addr_5_3, wires_20_4,addr_20_4);

wire[3:0] wires_21_4;

wire[27:0] addr_21_4;

Selector_2 s21_4(wires_5_3[1], addr_5_3, wires_21_4,addr_21_4);

wire[3:0] wires_22_4;

wire[27:0] addr_22_4;

Selector_2 s22_4(wires_5_3[2], addr_5_3, wires_22_4,addr_22_4);

wire[3:0] wires_23_4;

wire[27:0] addr_23_4;

Selector_2 s23_4(wires_5_3[3], addr_5_3, wires_23_4,addr_23_4);

wire[3:0] wires_24_4;

wire[27:0] addr_24_4;

Selector_2 s24_4(wires_6_3[0], addr_6_3, wires_24_4,addr_24_4);

wire[3:0] wires_25_4;

wire[27:0] addr_25_4;

Selector_2 s25_4(wires_6_3[1], addr_6_3, wires_25_4,addr_25_4);

wire[3:0] wires_26_4;

wire[27:0] addr_26_4;

Selector_2 s26_4(wires_6_3[2], addr_6_3, wires_26_4,addr_26_4);

wire[3:0] wires_27_4;

wire[27:0] addr_27_4;

Selector_2 s27_4(wires_6_3[3], addr_6_3, wires_27_4,addr_27_4);

wire[3:0] wires_28_4;

wire[27:0] addr_28_4;

Selector_2 s28_4(wires_7_3[0], addr_7_3, wires_28_4,addr_28_4);

wire[3:0] wires_29_4;

wire[27:0] addr_29_4;

Selector_2 s29_4(wires_7_3[1], addr_7_3, wires_29_4,addr_29_4);

wire[3:0] wires_30_4;

wire[27:0] addr_30_4;

Selector_2 s30_4(wires_7_3[2], addr_7_3, wires_30_4,addr_30_4);

wire[3:0] wires_31_4;

wire[27:0] addr_31_4;

Selector_2 s31_4(wires_7_3[3], addr_7_3, wires_31_4,addr_31_4);

wire[3:0] wires_32_4;

wire[27:0] addr_32_4;

Selector_2 s32_4(wires_8_3[0], addr_8_3, wires_32_4,addr_32_4);

wire[3:0] wires_33_4;

wire[27:0] addr_33_4;

Selector_2 s33_4(wires_8_3[1], addr_8_3, wires_33_4,addr_33_4);

wire[3:0] wires_34_4;

wire[27:0] addr_34_4;

Selector_2 s34_4(wires_8_3[2], addr_8_3, wires_34_4,addr_34_4);

wire[3:0] wires_35_4;

wire[27:0] addr_35_4;

Selector_2 s35_4(wires_8_3[3], addr_8_3, wires_35_4,addr_35_4);

wire[3:0] wires_36_4;

wire[27:0] addr_36_4;

Selector_2 s36_4(wires_9_3[0], addr_9_3, wires_36_4,addr_36_4);

wire[3:0] wires_37_4;

wire[27:0] addr_37_4;

Selector_2 s37_4(wires_9_3[1], addr_9_3, wires_37_4,addr_37_4);

wire[3:0] wires_38_4;

wire[27:0] addr_38_4;

Selector_2 s38_4(wires_9_3[2], addr_9_3, wires_38_4,addr_38_4);

wire[3:0] wires_39_4;

wire[27:0] addr_39_4;

Selector_2 s39_4(wires_9_3[3], addr_9_3, wires_39_4,addr_39_4);

wire[3:0] wires_40_4;

wire[27:0] addr_40_4;

Selector_2 s40_4(wires_10_3[0], addr_10_3, wires_40_4,addr_40_4);

wire[3:0] wires_41_4;

wire[27:0] addr_41_4;

Selector_2 s41_4(wires_10_3[1], addr_10_3, wires_41_4,addr_41_4);

wire[3:0] wires_42_4;

wire[27:0] addr_42_4;

Selector_2 s42_4(wires_10_3[2], addr_10_3, wires_42_4,addr_42_4);

wire[3:0] wires_43_4;

wire[27:0] addr_43_4;

Selector_2 s43_4(wires_10_3[3], addr_10_3, wires_43_4,addr_43_4);

wire[3:0] wires_44_4;

wire[27:0] addr_44_4;

Selector_2 s44_4(wires_11_3[0], addr_11_3, wires_44_4,addr_44_4);

wire[3:0] wires_45_4;

wire[27:0] addr_45_4;

Selector_2 s45_4(wires_11_3[1], addr_11_3, wires_45_4,addr_45_4);

wire[3:0] wires_46_4;

wire[27:0] addr_46_4;

Selector_2 s46_4(wires_11_3[2], addr_11_3, wires_46_4,addr_46_4);

wire[3:0] wires_47_4;

wire[27:0] addr_47_4;

Selector_2 s47_4(wires_11_3[3], addr_11_3, wires_47_4,addr_47_4);

wire[3:0] wires_48_4;

wire[27:0] addr_48_4;

Selector_2 s48_4(wires_12_3[0], addr_12_3, wires_48_4,addr_48_4);

wire[3:0] wires_49_4;

wire[27:0] addr_49_4;

Selector_2 s49_4(wires_12_3[1], addr_12_3, wires_49_4,addr_49_4);

wire[3:0] wires_50_4;

wire[27:0] addr_50_4;

Selector_2 s50_4(wires_12_3[2], addr_12_3, wires_50_4,addr_50_4);

wire[3:0] wires_51_4;

wire[27:0] addr_51_4;

Selector_2 s51_4(wires_12_3[3], addr_12_3, wires_51_4,addr_51_4);

wire[3:0] wires_52_4;

wire[27:0] addr_52_4;

Selector_2 s52_4(wires_13_3[0], addr_13_3, wires_52_4,addr_52_4);

wire[3:0] wires_53_4;

wire[27:0] addr_53_4;

Selector_2 s53_4(wires_13_3[1], addr_13_3, wires_53_4,addr_53_4);

wire[3:0] wires_54_4;

wire[27:0] addr_54_4;

Selector_2 s54_4(wires_13_3[2], addr_13_3, wires_54_4,addr_54_4);

wire[3:0] wires_55_4;

wire[27:0] addr_55_4;

Selector_2 s55_4(wires_13_3[3], addr_13_3, wires_55_4,addr_55_4);

wire[3:0] wires_56_4;

wire[27:0] addr_56_4;

Selector_2 s56_4(wires_14_3[0], addr_14_3, wires_56_4,addr_56_4);

wire[3:0] wires_57_4;

wire[27:0] addr_57_4;

Selector_2 s57_4(wires_14_3[1], addr_14_3, wires_57_4,addr_57_4);

wire[3:0] wires_58_4;

wire[27:0] addr_58_4;

Selector_2 s58_4(wires_14_3[2], addr_14_3, wires_58_4,addr_58_4);

wire[3:0] wires_59_4;

wire[27:0] addr_59_4;

Selector_2 s59_4(wires_14_3[3], addr_14_3, wires_59_4,addr_59_4);

wire[3:0] wires_60_4;

wire[27:0] addr_60_4;

Selector_2 s60_4(wires_15_3[0], addr_15_3, wires_60_4,addr_60_4);

wire[3:0] wires_61_4;

wire[27:0] addr_61_4;

Selector_2 s61_4(wires_15_3[1], addr_15_3, wires_61_4,addr_61_4);

wire[3:0] wires_62_4;

wire[27:0] addr_62_4;

Selector_2 s62_4(wires_15_3[2], addr_15_3, wires_62_4,addr_62_4);

wire[3:0] wires_63_4;

wire[27:0] addr_63_4;

Selector_2 s63_4(wires_15_3[3], addr_15_3, wires_63_4,addr_63_4);

wire[3:0] wires_64_4;

wire[27:0] addr_64_4;

Selector_2 s64_4(wires_16_3[0], addr_16_3, wires_64_4,addr_64_4);

wire[3:0] wires_65_4;

wire[27:0] addr_65_4;

Selector_2 s65_4(wires_16_3[1], addr_16_3, wires_65_4,addr_65_4);

wire[3:0] wires_66_4;

wire[27:0] addr_66_4;

Selector_2 s66_4(wires_16_3[2], addr_16_3, wires_66_4,addr_66_4);

wire[3:0] wires_67_4;

wire[27:0] addr_67_4;

Selector_2 s67_4(wires_16_3[3], addr_16_3, wires_67_4,addr_67_4);

wire[3:0] wires_68_4;

wire[27:0] addr_68_4;

Selector_2 s68_4(wires_17_3[0], addr_17_3, wires_68_4,addr_68_4);

wire[3:0] wires_69_4;

wire[27:0] addr_69_4;

Selector_2 s69_4(wires_17_3[1], addr_17_3, wires_69_4,addr_69_4);

wire[3:0] wires_70_4;

wire[27:0] addr_70_4;

Selector_2 s70_4(wires_17_3[2], addr_17_3, wires_70_4,addr_70_4);

wire[3:0] wires_71_4;

wire[27:0] addr_71_4;

Selector_2 s71_4(wires_17_3[3], addr_17_3, wires_71_4,addr_71_4);

wire[3:0] wires_72_4;

wire[27:0] addr_72_4;

Selector_2 s72_4(wires_18_3[0], addr_18_3, wires_72_4,addr_72_4);

wire[3:0] wires_73_4;

wire[27:0] addr_73_4;

Selector_2 s73_4(wires_18_3[1], addr_18_3, wires_73_4,addr_73_4);

wire[3:0] wires_74_4;

wire[27:0] addr_74_4;

Selector_2 s74_4(wires_18_3[2], addr_18_3, wires_74_4,addr_74_4);

wire[3:0] wires_75_4;

wire[27:0] addr_75_4;

Selector_2 s75_4(wires_18_3[3], addr_18_3, wires_75_4,addr_75_4);

wire[3:0] wires_76_4;

wire[27:0] addr_76_4;

Selector_2 s76_4(wires_19_3[0], addr_19_3, wires_76_4,addr_76_4);

wire[3:0] wires_77_4;

wire[27:0] addr_77_4;

Selector_2 s77_4(wires_19_3[1], addr_19_3, wires_77_4,addr_77_4);

wire[3:0] wires_78_4;

wire[27:0] addr_78_4;

Selector_2 s78_4(wires_19_3[2], addr_19_3, wires_78_4,addr_78_4);

wire[3:0] wires_79_4;

wire[27:0] addr_79_4;

Selector_2 s79_4(wires_19_3[3], addr_19_3, wires_79_4,addr_79_4);

wire[3:0] wires_80_4;

wire[27:0] addr_80_4;

Selector_2 s80_4(wires_20_3[0], addr_20_3, wires_80_4,addr_80_4);

wire[3:0] wires_81_4;

wire[27:0] addr_81_4;

Selector_2 s81_4(wires_20_3[1], addr_20_3, wires_81_4,addr_81_4);

wire[3:0] wires_82_4;

wire[27:0] addr_82_4;

Selector_2 s82_4(wires_20_3[2], addr_20_3, wires_82_4,addr_82_4);

wire[3:0] wires_83_4;

wire[27:0] addr_83_4;

Selector_2 s83_4(wires_20_3[3], addr_20_3, wires_83_4,addr_83_4);

wire[3:0] wires_84_4;

wire[27:0] addr_84_4;

Selector_2 s84_4(wires_21_3[0], addr_21_3, wires_84_4,addr_84_4);

wire[3:0] wires_85_4;

wire[27:0] addr_85_4;

Selector_2 s85_4(wires_21_3[1], addr_21_3, wires_85_4,addr_85_4);

wire[3:0] wires_86_4;

wire[27:0] addr_86_4;

Selector_2 s86_4(wires_21_3[2], addr_21_3, wires_86_4,addr_86_4);

wire[3:0] wires_87_4;

wire[27:0] addr_87_4;

Selector_2 s87_4(wires_21_3[3], addr_21_3, wires_87_4,addr_87_4);

wire[3:0] wires_88_4;

wire[27:0] addr_88_4;

Selector_2 s88_4(wires_22_3[0], addr_22_3, wires_88_4,addr_88_4);

wire[3:0] wires_89_4;

wire[27:0] addr_89_4;

Selector_2 s89_4(wires_22_3[1], addr_22_3, wires_89_4,addr_89_4);

wire[3:0] wires_90_4;

wire[27:0] addr_90_4;

Selector_2 s90_4(wires_22_3[2], addr_22_3, wires_90_4,addr_90_4);

wire[3:0] wires_91_4;

wire[27:0] addr_91_4;

Selector_2 s91_4(wires_22_3[3], addr_22_3, wires_91_4,addr_91_4);

wire[3:0] wires_92_4;

wire[27:0] addr_92_4;

Selector_2 s92_4(wires_23_3[0], addr_23_3, wires_92_4,addr_92_4);

wire[3:0] wires_93_4;

wire[27:0] addr_93_4;

Selector_2 s93_4(wires_23_3[1], addr_23_3, wires_93_4,addr_93_4);

wire[3:0] wires_94_4;

wire[27:0] addr_94_4;

Selector_2 s94_4(wires_23_3[2], addr_23_3, wires_94_4,addr_94_4);

wire[3:0] wires_95_4;

wire[27:0] addr_95_4;

Selector_2 s95_4(wires_23_3[3], addr_23_3, wires_95_4,addr_95_4);

wire[3:0] wires_96_4;

wire[27:0] addr_96_4;

Selector_2 s96_4(wires_24_3[0], addr_24_3, wires_96_4,addr_96_4);

wire[3:0] wires_97_4;

wire[27:0] addr_97_4;

Selector_2 s97_4(wires_24_3[1], addr_24_3, wires_97_4,addr_97_4);

wire[3:0] wires_98_4;

wire[27:0] addr_98_4;

Selector_2 s98_4(wires_24_3[2], addr_24_3, wires_98_4,addr_98_4);

wire[3:0] wires_99_4;

wire[27:0] addr_99_4;

Selector_2 s99_4(wires_24_3[3], addr_24_3, wires_99_4,addr_99_4);

wire[3:0] wires_100_4;

wire[27:0] addr_100_4;

Selector_2 s100_4(wires_25_3[0], addr_25_3, wires_100_4,addr_100_4);

wire[3:0] wires_101_4;

wire[27:0] addr_101_4;

Selector_2 s101_4(wires_25_3[1], addr_25_3, wires_101_4,addr_101_4);

wire[3:0] wires_102_4;

wire[27:0] addr_102_4;

Selector_2 s102_4(wires_25_3[2], addr_25_3, wires_102_4,addr_102_4);

wire[3:0] wires_103_4;

wire[27:0] addr_103_4;

Selector_2 s103_4(wires_25_3[3], addr_25_3, wires_103_4,addr_103_4);

wire[3:0] wires_104_4;

wire[27:0] addr_104_4;

Selector_2 s104_4(wires_26_3[0], addr_26_3, wires_104_4,addr_104_4);

wire[3:0] wires_105_4;

wire[27:0] addr_105_4;

Selector_2 s105_4(wires_26_3[1], addr_26_3, wires_105_4,addr_105_4);

wire[3:0] wires_106_4;

wire[27:0] addr_106_4;

Selector_2 s106_4(wires_26_3[2], addr_26_3, wires_106_4,addr_106_4);

wire[3:0] wires_107_4;

wire[27:0] addr_107_4;

Selector_2 s107_4(wires_26_3[3], addr_26_3, wires_107_4,addr_107_4);

wire[3:0] wires_108_4;

wire[27:0] addr_108_4;

Selector_2 s108_4(wires_27_3[0], addr_27_3, wires_108_4,addr_108_4);

wire[3:0] wires_109_4;

wire[27:0] addr_109_4;

Selector_2 s109_4(wires_27_3[1], addr_27_3, wires_109_4,addr_109_4);

wire[3:0] wires_110_4;

wire[27:0] addr_110_4;

Selector_2 s110_4(wires_27_3[2], addr_27_3, wires_110_4,addr_110_4);

wire[3:0] wires_111_4;

wire[27:0] addr_111_4;

Selector_2 s111_4(wires_27_3[3], addr_27_3, wires_111_4,addr_111_4);

wire[3:0] wires_112_4;

wire[27:0] addr_112_4;

Selector_2 s112_4(wires_28_3[0], addr_28_3, wires_112_4,addr_112_4);

wire[3:0] wires_113_4;

wire[27:0] addr_113_4;

Selector_2 s113_4(wires_28_3[1], addr_28_3, wires_113_4,addr_113_4);

wire[3:0] wires_114_4;

wire[27:0] addr_114_4;

Selector_2 s114_4(wires_28_3[2], addr_28_3, wires_114_4,addr_114_4);

wire[3:0] wires_115_4;

wire[27:0] addr_115_4;

Selector_2 s115_4(wires_28_3[3], addr_28_3, wires_115_4,addr_115_4);

wire[3:0] wires_116_4;

wire[27:0] addr_116_4;

Selector_2 s116_4(wires_29_3[0], addr_29_3, wires_116_4,addr_116_4);

wire[3:0] wires_117_4;

wire[27:0] addr_117_4;

Selector_2 s117_4(wires_29_3[1], addr_29_3, wires_117_4,addr_117_4);

wire[3:0] wires_118_4;

wire[27:0] addr_118_4;

Selector_2 s118_4(wires_29_3[2], addr_29_3, wires_118_4,addr_118_4);

wire[3:0] wires_119_4;

wire[27:0] addr_119_4;

Selector_2 s119_4(wires_29_3[3], addr_29_3, wires_119_4,addr_119_4);

wire[3:0] wires_120_4;

wire[27:0] addr_120_4;

Selector_2 s120_4(wires_30_3[0], addr_30_3, wires_120_4,addr_120_4);

wire[3:0] wires_121_4;

wire[27:0] addr_121_4;

Selector_2 s121_4(wires_30_3[1], addr_30_3, wires_121_4,addr_121_4);

wire[3:0] wires_122_4;

wire[27:0] addr_122_4;

Selector_2 s122_4(wires_30_3[2], addr_30_3, wires_122_4,addr_122_4);

wire[3:0] wires_123_4;

wire[27:0] addr_123_4;

Selector_2 s123_4(wires_30_3[3], addr_30_3, wires_123_4,addr_123_4);

wire[3:0] wires_124_4;

wire[27:0] addr_124_4;

Selector_2 s124_4(wires_31_3[0], addr_31_3, wires_124_4,addr_124_4);

wire[3:0] wires_125_4;

wire[27:0] addr_125_4;

Selector_2 s125_4(wires_31_3[1], addr_31_3, wires_125_4,addr_125_4);

wire[3:0] wires_126_4;

wire[27:0] addr_126_4;

Selector_2 s126_4(wires_31_3[2], addr_31_3, wires_126_4,addr_126_4);

wire[3:0] wires_127_4;

wire[27:0] addr_127_4;

Selector_2 s127_4(wires_31_3[3], addr_31_3, wires_127_4,addr_127_4);

wire[3:0] wires_128_4;

wire[27:0] addr_128_4;

Selector_2 s128_4(wires_32_3[0], addr_32_3, wires_128_4,addr_128_4);

wire[3:0] wires_129_4;

wire[27:0] addr_129_4;

Selector_2 s129_4(wires_32_3[1], addr_32_3, wires_129_4,addr_129_4);

wire[3:0] wires_130_4;

wire[27:0] addr_130_4;

Selector_2 s130_4(wires_32_3[2], addr_32_3, wires_130_4,addr_130_4);

wire[3:0] wires_131_4;

wire[27:0] addr_131_4;

Selector_2 s131_4(wires_32_3[3], addr_32_3, wires_131_4,addr_131_4);

wire[3:0] wires_132_4;

wire[27:0] addr_132_4;

Selector_2 s132_4(wires_33_3[0], addr_33_3, wires_132_4,addr_132_4);

wire[3:0] wires_133_4;

wire[27:0] addr_133_4;

Selector_2 s133_4(wires_33_3[1], addr_33_3, wires_133_4,addr_133_4);

wire[3:0] wires_134_4;

wire[27:0] addr_134_4;

Selector_2 s134_4(wires_33_3[2], addr_33_3, wires_134_4,addr_134_4);

wire[3:0] wires_135_4;

wire[27:0] addr_135_4;

Selector_2 s135_4(wires_33_3[3], addr_33_3, wires_135_4,addr_135_4);

wire[3:0] wires_136_4;

wire[27:0] addr_136_4;

Selector_2 s136_4(wires_34_3[0], addr_34_3, wires_136_4,addr_136_4);

wire[3:0] wires_137_4;

wire[27:0] addr_137_4;

Selector_2 s137_4(wires_34_3[1], addr_34_3, wires_137_4,addr_137_4);

wire[3:0] wires_138_4;

wire[27:0] addr_138_4;

Selector_2 s138_4(wires_34_3[2], addr_34_3, wires_138_4,addr_138_4);

wire[3:0] wires_139_4;

wire[27:0] addr_139_4;

Selector_2 s139_4(wires_34_3[3], addr_34_3, wires_139_4,addr_139_4);

wire[3:0] wires_140_4;

wire[27:0] addr_140_4;

Selector_2 s140_4(wires_35_3[0], addr_35_3, wires_140_4,addr_140_4);

wire[3:0] wires_141_4;

wire[27:0] addr_141_4;

Selector_2 s141_4(wires_35_3[1], addr_35_3, wires_141_4,addr_141_4);

wire[3:0] wires_142_4;

wire[27:0] addr_142_4;

Selector_2 s142_4(wires_35_3[2], addr_35_3, wires_142_4,addr_142_4);

wire[3:0] wires_143_4;

wire[27:0] addr_143_4;

Selector_2 s143_4(wires_35_3[3], addr_35_3, wires_143_4,addr_143_4);

wire[3:0] wires_144_4;

wire[27:0] addr_144_4;

Selector_2 s144_4(wires_36_3[0], addr_36_3, wires_144_4,addr_144_4);

wire[3:0] wires_145_4;

wire[27:0] addr_145_4;

Selector_2 s145_4(wires_36_3[1], addr_36_3, wires_145_4,addr_145_4);

wire[3:0] wires_146_4;

wire[27:0] addr_146_4;

Selector_2 s146_4(wires_36_3[2], addr_36_3, wires_146_4,addr_146_4);

wire[3:0] wires_147_4;

wire[27:0] addr_147_4;

Selector_2 s147_4(wires_36_3[3], addr_36_3, wires_147_4,addr_147_4);

wire[3:0] wires_148_4;

wire[27:0] addr_148_4;

Selector_2 s148_4(wires_37_3[0], addr_37_3, wires_148_4,addr_148_4);

wire[3:0] wires_149_4;

wire[27:0] addr_149_4;

Selector_2 s149_4(wires_37_3[1], addr_37_3, wires_149_4,addr_149_4);

wire[3:0] wires_150_4;

wire[27:0] addr_150_4;

Selector_2 s150_4(wires_37_3[2], addr_37_3, wires_150_4,addr_150_4);

wire[3:0] wires_151_4;

wire[27:0] addr_151_4;

Selector_2 s151_4(wires_37_3[3], addr_37_3, wires_151_4,addr_151_4);

wire[3:0] wires_152_4;

wire[27:0] addr_152_4;

Selector_2 s152_4(wires_38_3[0], addr_38_3, wires_152_4,addr_152_4);

wire[3:0] wires_153_4;

wire[27:0] addr_153_4;

Selector_2 s153_4(wires_38_3[1], addr_38_3, wires_153_4,addr_153_4);

wire[3:0] wires_154_4;

wire[27:0] addr_154_4;

Selector_2 s154_4(wires_38_3[2], addr_38_3, wires_154_4,addr_154_4);

wire[3:0] wires_155_4;

wire[27:0] addr_155_4;

Selector_2 s155_4(wires_38_3[3], addr_38_3, wires_155_4,addr_155_4);

wire[3:0] wires_156_4;

wire[27:0] addr_156_4;

Selector_2 s156_4(wires_39_3[0], addr_39_3, wires_156_4,addr_156_4);

wire[3:0] wires_157_4;

wire[27:0] addr_157_4;

Selector_2 s157_4(wires_39_3[1], addr_39_3, wires_157_4,addr_157_4);

wire[3:0] wires_158_4;

wire[27:0] addr_158_4;

Selector_2 s158_4(wires_39_3[2], addr_39_3, wires_158_4,addr_158_4);

wire[3:0] wires_159_4;

wire[27:0] addr_159_4;

Selector_2 s159_4(wires_39_3[3], addr_39_3, wires_159_4,addr_159_4);

wire[3:0] wires_160_4;

wire[27:0] addr_160_4;

Selector_2 s160_4(wires_40_3[0], addr_40_3, wires_160_4,addr_160_4);

wire[3:0] wires_161_4;

wire[27:0] addr_161_4;

Selector_2 s161_4(wires_40_3[1], addr_40_3, wires_161_4,addr_161_4);

wire[3:0] wires_162_4;

wire[27:0] addr_162_4;

Selector_2 s162_4(wires_40_3[2], addr_40_3, wires_162_4,addr_162_4);

wire[3:0] wires_163_4;

wire[27:0] addr_163_4;

Selector_2 s163_4(wires_40_3[3], addr_40_3, wires_163_4,addr_163_4);

wire[3:0] wires_164_4;

wire[27:0] addr_164_4;

Selector_2 s164_4(wires_41_3[0], addr_41_3, wires_164_4,addr_164_4);

wire[3:0] wires_165_4;

wire[27:0] addr_165_4;

Selector_2 s165_4(wires_41_3[1], addr_41_3, wires_165_4,addr_165_4);

wire[3:0] wires_166_4;

wire[27:0] addr_166_4;

Selector_2 s166_4(wires_41_3[2], addr_41_3, wires_166_4,addr_166_4);

wire[3:0] wires_167_4;

wire[27:0] addr_167_4;

Selector_2 s167_4(wires_41_3[3], addr_41_3, wires_167_4,addr_167_4);

wire[3:0] wires_168_4;

wire[27:0] addr_168_4;

Selector_2 s168_4(wires_42_3[0], addr_42_3, wires_168_4,addr_168_4);

wire[3:0] wires_169_4;

wire[27:0] addr_169_4;

Selector_2 s169_4(wires_42_3[1], addr_42_3, wires_169_4,addr_169_4);

wire[3:0] wires_170_4;

wire[27:0] addr_170_4;

Selector_2 s170_4(wires_42_3[2], addr_42_3, wires_170_4,addr_170_4);

wire[3:0] wires_171_4;

wire[27:0] addr_171_4;

Selector_2 s171_4(wires_42_3[3], addr_42_3, wires_171_4,addr_171_4);

wire[3:0] wires_172_4;

wire[27:0] addr_172_4;

Selector_2 s172_4(wires_43_3[0], addr_43_3, wires_172_4,addr_172_4);

wire[3:0] wires_173_4;

wire[27:0] addr_173_4;

Selector_2 s173_4(wires_43_3[1], addr_43_3, wires_173_4,addr_173_4);

wire[3:0] wires_174_4;

wire[27:0] addr_174_4;

Selector_2 s174_4(wires_43_3[2], addr_43_3, wires_174_4,addr_174_4);

wire[3:0] wires_175_4;

wire[27:0] addr_175_4;

Selector_2 s175_4(wires_43_3[3], addr_43_3, wires_175_4,addr_175_4);

wire[3:0] wires_176_4;

wire[27:0] addr_176_4;

Selector_2 s176_4(wires_44_3[0], addr_44_3, wires_176_4,addr_176_4);

wire[3:0] wires_177_4;

wire[27:0] addr_177_4;

Selector_2 s177_4(wires_44_3[1], addr_44_3, wires_177_4,addr_177_4);

wire[3:0] wires_178_4;

wire[27:0] addr_178_4;

Selector_2 s178_4(wires_44_3[2], addr_44_3, wires_178_4,addr_178_4);

wire[3:0] wires_179_4;

wire[27:0] addr_179_4;

Selector_2 s179_4(wires_44_3[3], addr_44_3, wires_179_4,addr_179_4);

wire[3:0] wires_180_4;

wire[27:0] addr_180_4;

Selector_2 s180_4(wires_45_3[0], addr_45_3, wires_180_4,addr_180_4);

wire[3:0] wires_181_4;

wire[27:0] addr_181_4;

Selector_2 s181_4(wires_45_3[1], addr_45_3, wires_181_4,addr_181_4);

wire[3:0] wires_182_4;

wire[27:0] addr_182_4;

Selector_2 s182_4(wires_45_3[2], addr_45_3, wires_182_4,addr_182_4);

wire[3:0] wires_183_4;

wire[27:0] addr_183_4;

Selector_2 s183_4(wires_45_3[3], addr_45_3, wires_183_4,addr_183_4);

wire[3:0] wires_184_4;

wire[27:0] addr_184_4;

Selector_2 s184_4(wires_46_3[0], addr_46_3, wires_184_4,addr_184_4);

wire[3:0] wires_185_4;

wire[27:0] addr_185_4;

Selector_2 s185_4(wires_46_3[1], addr_46_3, wires_185_4,addr_185_4);

wire[3:0] wires_186_4;

wire[27:0] addr_186_4;

Selector_2 s186_4(wires_46_3[2], addr_46_3, wires_186_4,addr_186_4);

wire[3:0] wires_187_4;

wire[27:0] addr_187_4;

Selector_2 s187_4(wires_46_3[3], addr_46_3, wires_187_4,addr_187_4);

wire[3:0] wires_188_4;

wire[27:0] addr_188_4;

Selector_2 s188_4(wires_47_3[0], addr_47_3, wires_188_4,addr_188_4);

wire[3:0] wires_189_4;

wire[27:0] addr_189_4;

Selector_2 s189_4(wires_47_3[1], addr_47_3, wires_189_4,addr_189_4);

wire[3:0] wires_190_4;

wire[27:0] addr_190_4;

Selector_2 s190_4(wires_47_3[2], addr_47_3, wires_190_4,addr_190_4);

wire[3:0] wires_191_4;

wire[27:0] addr_191_4;

Selector_2 s191_4(wires_47_3[3], addr_47_3, wires_191_4,addr_191_4);

wire[3:0] wires_192_4;

wire[27:0] addr_192_4;

Selector_2 s192_4(wires_48_3[0], addr_48_3, wires_192_4,addr_192_4);

wire[3:0] wires_193_4;

wire[27:0] addr_193_4;

Selector_2 s193_4(wires_48_3[1], addr_48_3, wires_193_4,addr_193_4);

wire[3:0] wires_194_4;

wire[27:0] addr_194_4;

Selector_2 s194_4(wires_48_3[2], addr_48_3, wires_194_4,addr_194_4);

wire[3:0] wires_195_4;

wire[27:0] addr_195_4;

Selector_2 s195_4(wires_48_3[3], addr_48_3, wires_195_4,addr_195_4);

wire[3:0] wires_196_4;

wire[27:0] addr_196_4;

Selector_2 s196_4(wires_49_3[0], addr_49_3, wires_196_4,addr_196_4);

wire[3:0] wires_197_4;

wire[27:0] addr_197_4;

Selector_2 s197_4(wires_49_3[1], addr_49_3, wires_197_4,addr_197_4);

wire[3:0] wires_198_4;

wire[27:0] addr_198_4;

Selector_2 s198_4(wires_49_3[2], addr_49_3, wires_198_4,addr_198_4);

wire[3:0] wires_199_4;

wire[27:0] addr_199_4;

Selector_2 s199_4(wires_49_3[3], addr_49_3, wires_199_4,addr_199_4);

wire[3:0] wires_200_4;

wire[27:0] addr_200_4;

Selector_2 s200_4(wires_50_3[0], addr_50_3, wires_200_4,addr_200_4);

wire[3:0] wires_201_4;

wire[27:0] addr_201_4;

Selector_2 s201_4(wires_50_3[1], addr_50_3, wires_201_4,addr_201_4);

wire[3:0] wires_202_4;

wire[27:0] addr_202_4;

Selector_2 s202_4(wires_50_3[2], addr_50_3, wires_202_4,addr_202_4);

wire[3:0] wires_203_4;

wire[27:0] addr_203_4;

Selector_2 s203_4(wires_50_3[3], addr_50_3, wires_203_4,addr_203_4);

wire[3:0] wires_204_4;

wire[27:0] addr_204_4;

Selector_2 s204_4(wires_51_3[0], addr_51_3, wires_204_4,addr_204_4);

wire[3:0] wires_205_4;

wire[27:0] addr_205_4;

Selector_2 s205_4(wires_51_3[1], addr_51_3, wires_205_4,addr_205_4);

wire[3:0] wires_206_4;

wire[27:0] addr_206_4;

Selector_2 s206_4(wires_51_3[2], addr_51_3, wires_206_4,addr_206_4);

wire[3:0] wires_207_4;

wire[27:0] addr_207_4;

Selector_2 s207_4(wires_51_3[3], addr_51_3, wires_207_4,addr_207_4);

wire[3:0] wires_208_4;

wire[27:0] addr_208_4;

Selector_2 s208_4(wires_52_3[0], addr_52_3, wires_208_4,addr_208_4);

wire[3:0] wires_209_4;

wire[27:0] addr_209_4;

Selector_2 s209_4(wires_52_3[1], addr_52_3, wires_209_4,addr_209_4);

wire[3:0] wires_210_4;

wire[27:0] addr_210_4;

Selector_2 s210_4(wires_52_3[2], addr_52_3, wires_210_4,addr_210_4);

wire[3:0] wires_211_4;

wire[27:0] addr_211_4;

Selector_2 s211_4(wires_52_3[3], addr_52_3, wires_211_4,addr_211_4);

wire[3:0] wires_212_4;

wire[27:0] addr_212_4;

Selector_2 s212_4(wires_53_3[0], addr_53_3, wires_212_4,addr_212_4);

wire[3:0] wires_213_4;

wire[27:0] addr_213_4;

Selector_2 s213_4(wires_53_3[1], addr_53_3, wires_213_4,addr_213_4);

wire[3:0] wires_214_4;

wire[27:0] addr_214_4;

Selector_2 s214_4(wires_53_3[2], addr_53_3, wires_214_4,addr_214_4);

wire[3:0] wires_215_4;

wire[27:0] addr_215_4;

Selector_2 s215_4(wires_53_3[3], addr_53_3, wires_215_4,addr_215_4);

wire[3:0] wires_216_4;

wire[27:0] addr_216_4;

Selector_2 s216_4(wires_54_3[0], addr_54_3, wires_216_4,addr_216_4);

wire[3:0] wires_217_4;

wire[27:0] addr_217_4;

Selector_2 s217_4(wires_54_3[1], addr_54_3, wires_217_4,addr_217_4);

wire[3:0] wires_218_4;

wire[27:0] addr_218_4;

Selector_2 s218_4(wires_54_3[2], addr_54_3, wires_218_4,addr_218_4);

wire[3:0] wires_219_4;

wire[27:0] addr_219_4;

Selector_2 s219_4(wires_54_3[3], addr_54_3, wires_219_4,addr_219_4);

wire[3:0] wires_220_4;

wire[27:0] addr_220_4;

Selector_2 s220_4(wires_55_3[0], addr_55_3, wires_220_4,addr_220_4);

wire[3:0] wires_221_4;

wire[27:0] addr_221_4;

Selector_2 s221_4(wires_55_3[1], addr_55_3, wires_221_4,addr_221_4);

wire[3:0] wires_222_4;

wire[27:0] addr_222_4;

Selector_2 s222_4(wires_55_3[2], addr_55_3, wires_222_4,addr_222_4);

wire[3:0] wires_223_4;

wire[27:0] addr_223_4;

Selector_2 s223_4(wires_55_3[3], addr_55_3, wires_223_4,addr_223_4);

wire[3:0] wires_224_4;

wire[27:0] addr_224_4;

Selector_2 s224_4(wires_56_3[0], addr_56_3, wires_224_4,addr_224_4);

wire[3:0] wires_225_4;

wire[27:0] addr_225_4;

Selector_2 s225_4(wires_56_3[1], addr_56_3, wires_225_4,addr_225_4);

wire[3:0] wires_226_4;

wire[27:0] addr_226_4;

Selector_2 s226_4(wires_56_3[2], addr_56_3, wires_226_4,addr_226_4);

wire[3:0] wires_227_4;

wire[27:0] addr_227_4;

Selector_2 s227_4(wires_56_3[3], addr_56_3, wires_227_4,addr_227_4);

wire[3:0] wires_228_4;

wire[27:0] addr_228_4;

Selector_2 s228_4(wires_57_3[0], addr_57_3, wires_228_4,addr_228_4);

wire[3:0] wires_229_4;

wire[27:0] addr_229_4;

Selector_2 s229_4(wires_57_3[1], addr_57_3, wires_229_4,addr_229_4);

wire[3:0] wires_230_4;

wire[27:0] addr_230_4;

Selector_2 s230_4(wires_57_3[2], addr_57_3, wires_230_4,addr_230_4);

wire[3:0] wires_231_4;

wire[27:0] addr_231_4;

Selector_2 s231_4(wires_57_3[3], addr_57_3, wires_231_4,addr_231_4);

wire[3:0] wires_232_4;

wire[27:0] addr_232_4;

Selector_2 s232_4(wires_58_3[0], addr_58_3, wires_232_4,addr_232_4);

wire[3:0] wires_233_4;

wire[27:0] addr_233_4;

Selector_2 s233_4(wires_58_3[1], addr_58_3, wires_233_4,addr_233_4);

wire[3:0] wires_234_4;

wire[27:0] addr_234_4;

Selector_2 s234_4(wires_58_3[2], addr_58_3, wires_234_4,addr_234_4);

wire[3:0] wires_235_4;

wire[27:0] addr_235_4;

Selector_2 s235_4(wires_58_3[3], addr_58_3, wires_235_4,addr_235_4);

wire[3:0] wires_236_4;

wire[27:0] addr_236_4;

Selector_2 s236_4(wires_59_3[0], addr_59_3, wires_236_4,addr_236_4);

wire[3:0] wires_237_4;

wire[27:0] addr_237_4;

Selector_2 s237_4(wires_59_3[1], addr_59_3, wires_237_4,addr_237_4);

wire[3:0] wires_238_4;

wire[27:0] addr_238_4;

Selector_2 s238_4(wires_59_3[2], addr_59_3, wires_238_4,addr_238_4);

wire[3:0] wires_239_4;

wire[27:0] addr_239_4;

Selector_2 s239_4(wires_59_3[3], addr_59_3, wires_239_4,addr_239_4);

wire[3:0] wires_240_4;

wire[27:0] addr_240_4;

Selector_2 s240_4(wires_60_3[0], addr_60_3, wires_240_4,addr_240_4);

wire[3:0] wires_241_4;

wire[27:0] addr_241_4;

Selector_2 s241_4(wires_60_3[1], addr_60_3, wires_241_4,addr_241_4);

wire[3:0] wires_242_4;

wire[27:0] addr_242_4;

Selector_2 s242_4(wires_60_3[2], addr_60_3, wires_242_4,addr_242_4);

wire[3:0] wires_243_4;

wire[27:0] addr_243_4;

Selector_2 s243_4(wires_60_3[3], addr_60_3, wires_243_4,addr_243_4);

wire[3:0] wires_244_4;

wire[27:0] addr_244_4;

Selector_2 s244_4(wires_61_3[0], addr_61_3, wires_244_4,addr_244_4);

wire[3:0] wires_245_4;

wire[27:0] addr_245_4;

Selector_2 s245_4(wires_61_3[1], addr_61_3, wires_245_4,addr_245_4);

wire[3:0] wires_246_4;

wire[27:0] addr_246_4;

Selector_2 s246_4(wires_61_3[2], addr_61_3, wires_246_4,addr_246_4);

wire[3:0] wires_247_4;

wire[27:0] addr_247_4;

Selector_2 s247_4(wires_61_3[3], addr_61_3, wires_247_4,addr_247_4);

wire[3:0] wires_248_4;

wire[27:0] addr_248_4;

Selector_2 s248_4(wires_62_3[0], addr_62_3, wires_248_4,addr_248_4);

wire[3:0] wires_249_4;

wire[27:0] addr_249_4;

Selector_2 s249_4(wires_62_3[1], addr_62_3, wires_249_4,addr_249_4);

wire[3:0] wires_250_4;

wire[27:0] addr_250_4;

Selector_2 s250_4(wires_62_3[2], addr_62_3, wires_250_4,addr_250_4);

wire[3:0] wires_251_4;

wire[27:0] addr_251_4;

Selector_2 s251_4(wires_62_3[3], addr_62_3, wires_251_4,addr_251_4);

wire[3:0] wires_252_4;

wire[27:0] addr_252_4;

Selector_2 s252_4(wires_63_3[0], addr_63_3, wires_252_4,addr_252_4);

wire[3:0] wires_253_4;

wire[27:0] addr_253_4;

Selector_2 s253_4(wires_63_3[1], addr_63_3, wires_253_4,addr_253_4);

wire[3:0] wires_254_4;

wire[27:0] addr_254_4;

Selector_2 s254_4(wires_63_3[2], addr_63_3, wires_254_4,addr_254_4);

wire[3:0] wires_255_4;

wire[27:0] addr_255_4;

Selector_2 s255_4(wires_63_3[3], addr_63_3, wires_255_4,addr_255_4);

wire[3:0] wires_0_5;

wire[27:0] addr_0_5;

Selector_2 s0_5(wires_0_4[0], addr_0_4, wires_0_5,addr_0_5);

wire[3:0] wires_1_5;

wire[27:0] addr_1_5;

Selector_2 s1_5(wires_0_4[1], addr_0_4, wires_1_5,addr_1_5);

wire[3:0] wires_2_5;

wire[27:0] addr_2_5;

Selector_2 s2_5(wires_0_4[2], addr_0_4, wires_2_5,addr_2_5);

wire[3:0] wires_3_5;

wire[27:0] addr_3_5;

Selector_2 s3_5(wires_0_4[3], addr_0_4, wires_3_5,addr_3_5);

wire[3:0] wires_4_5;

wire[27:0] addr_4_5;

Selector_2 s4_5(wires_1_4[0], addr_1_4, wires_4_5,addr_4_5);

wire[3:0] wires_5_5;

wire[27:0] addr_5_5;

Selector_2 s5_5(wires_1_4[1], addr_1_4, wires_5_5,addr_5_5);

wire[3:0] wires_6_5;

wire[27:0] addr_6_5;

Selector_2 s6_5(wires_1_4[2], addr_1_4, wires_6_5,addr_6_5);

wire[3:0] wires_7_5;

wire[27:0] addr_7_5;

Selector_2 s7_5(wires_1_4[3], addr_1_4, wires_7_5,addr_7_5);

wire[3:0] wires_8_5;

wire[27:0] addr_8_5;

Selector_2 s8_5(wires_2_4[0], addr_2_4, wires_8_5,addr_8_5);

wire[3:0] wires_9_5;

wire[27:0] addr_9_5;

Selector_2 s9_5(wires_2_4[1], addr_2_4, wires_9_5,addr_9_5);

wire[3:0] wires_10_5;

wire[27:0] addr_10_5;

Selector_2 s10_5(wires_2_4[2], addr_2_4, wires_10_5,addr_10_5);

wire[3:0] wires_11_5;

wire[27:0] addr_11_5;

Selector_2 s11_5(wires_2_4[3], addr_2_4, wires_11_5,addr_11_5);

wire[3:0] wires_12_5;

wire[27:0] addr_12_5;

Selector_2 s12_5(wires_3_4[0], addr_3_4, wires_12_5,addr_12_5);

wire[3:0] wires_13_5;

wire[27:0] addr_13_5;

Selector_2 s13_5(wires_3_4[1], addr_3_4, wires_13_5,addr_13_5);

wire[3:0] wires_14_5;

wire[27:0] addr_14_5;

Selector_2 s14_5(wires_3_4[2], addr_3_4, wires_14_5,addr_14_5);

wire[3:0] wires_15_5;

wire[27:0] addr_15_5;

Selector_2 s15_5(wires_3_4[3], addr_3_4, wires_15_5,addr_15_5);

wire[3:0] wires_16_5;

wire[27:0] addr_16_5;

Selector_2 s16_5(wires_4_4[0], addr_4_4, wires_16_5,addr_16_5);

wire[3:0] wires_17_5;

wire[27:0] addr_17_5;

Selector_2 s17_5(wires_4_4[1], addr_4_4, wires_17_5,addr_17_5);

wire[3:0] wires_18_5;

wire[27:0] addr_18_5;

Selector_2 s18_5(wires_4_4[2], addr_4_4, wires_18_5,addr_18_5);

wire[3:0] wires_19_5;

wire[27:0] addr_19_5;

Selector_2 s19_5(wires_4_4[3], addr_4_4, wires_19_5,addr_19_5);

wire[3:0] wires_20_5;

wire[27:0] addr_20_5;

Selector_2 s20_5(wires_5_4[0], addr_5_4, wires_20_5,addr_20_5);

wire[3:0] wires_21_5;

wire[27:0] addr_21_5;

Selector_2 s21_5(wires_5_4[1], addr_5_4, wires_21_5,addr_21_5);

wire[3:0] wires_22_5;

wire[27:0] addr_22_5;

Selector_2 s22_5(wires_5_4[2], addr_5_4, wires_22_5,addr_22_5);

wire[3:0] wires_23_5;

wire[27:0] addr_23_5;

Selector_2 s23_5(wires_5_4[3], addr_5_4, wires_23_5,addr_23_5);

wire[3:0] wires_24_5;

wire[27:0] addr_24_5;

Selector_2 s24_5(wires_6_4[0], addr_6_4, wires_24_5,addr_24_5);

wire[3:0] wires_25_5;

wire[27:0] addr_25_5;

Selector_2 s25_5(wires_6_4[1], addr_6_4, wires_25_5,addr_25_5);

wire[3:0] wires_26_5;

wire[27:0] addr_26_5;

Selector_2 s26_5(wires_6_4[2], addr_6_4, wires_26_5,addr_26_5);

wire[3:0] wires_27_5;

wire[27:0] addr_27_5;

Selector_2 s27_5(wires_6_4[3], addr_6_4, wires_27_5,addr_27_5);

wire[3:0] wires_28_5;

wire[27:0] addr_28_5;

Selector_2 s28_5(wires_7_4[0], addr_7_4, wires_28_5,addr_28_5);

wire[3:0] wires_29_5;

wire[27:0] addr_29_5;

Selector_2 s29_5(wires_7_4[1], addr_7_4, wires_29_5,addr_29_5);

wire[3:0] wires_30_5;

wire[27:0] addr_30_5;

Selector_2 s30_5(wires_7_4[2], addr_7_4, wires_30_5,addr_30_5);

wire[3:0] wires_31_5;

wire[27:0] addr_31_5;

Selector_2 s31_5(wires_7_4[3], addr_7_4, wires_31_5,addr_31_5);

wire[3:0] wires_32_5;

wire[27:0] addr_32_5;

Selector_2 s32_5(wires_8_4[0], addr_8_4, wires_32_5,addr_32_5);

wire[3:0] wires_33_5;

wire[27:0] addr_33_5;

Selector_2 s33_5(wires_8_4[1], addr_8_4, wires_33_5,addr_33_5);

wire[3:0] wires_34_5;

wire[27:0] addr_34_5;

Selector_2 s34_5(wires_8_4[2], addr_8_4, wires_34_5,addr_34_5);

wire[3:0] wires_35_5;

wire[27:0] addr_35_5;

Selector_2 s35_5(wires_8_4[3], addr_8_4, wires_35_5,addr_35_5);

wire[3:0] wires_36_5;

wire[27:0] addr_36_5;

Selector_2 s36_5(wires_9_4[0], addr_9_4, wires_36_5,addr_36_5);

wire[3:0] wires_37_5;

wire[27:0] addr_37_5;

Selector_2 s37_5(wires_9_4[1], addr_9_4, wires_37_5,addr_37_5);

wire[3:0] wires_38_5;

wire[27:0] addr_38_5;

Selector_2 s38_5(wires_9_4[2], addr_9_4, wires_38_5,addr_38_5);

wire[3:0] wires_39_5;

wire[27:0] addr_39_5;

Selector_2 s39_5(wires_9_4[3], addr_9_4, wires_39_5,addr_39_5);

wire[3:0] wires_40_5;

wire[27:0] addr_40_5;

Selector_2 s40_5(wires_10_4[0], addr_10_4, wires_40_5,addr_40_5);

wire[3:0] wires_41_5;

wire[27:0] addr_41_5;

Selector_2 s41_5(wires_10_4[1], addr_10_4, wires_41_5,addr_41_5);

wire[3:0] wires_42_5;

wire[27:0] addr_42_5;

Selector_2 s42_5(wires_10_4[2], addr_10_4, wires_42_5,addr_42_5);

wire[3:0] wires_43_5;

wire[27:0] addr_43_5;

Selector_2 s43_5(wires_10_4[3], addr_10_4, wires_43_5,addr_43_5);

wire[3:0] wires_44_5;

wire[27:0] addr_44_5;

Selector_2 s44_5(wires_11_4[0], addr_11_4, wires_44_5,addr_44_5);

wire[3:0] wires_45_5;

wire[27:0] addr_45_5;

Selector_2 s45_5(wires_11_4[1], addr_11_4, wires_45_5,addr_45_5);

wire[3:0] wires_46_5;

wire[27:0] addr_46_5;

Selector_2 s46_5(wires_11_4[2], addr_11_4, wires_46_5,addr_46_5);

wire[3:0] wires_47_5;

wire[27:0] addr_47_5;

Selector_2 s47_5(wires_11_4[3], addr_11_4, wires_47_5,addr_47_5);

wire[3:0] wires_48_5;

wire[27:0] addr_48_5;

Selector_2 s48_5(wires_12_4[0], addr_12_4, wires_48_5,addr_48_5);

wire[3:0] wires_49_5;

wire[27:0] addr_49_5;

Selector_2 s49_5(wires_12_4[1], addr_12_4, wires_49_5,addr_49_5);

wire[3:0] wires_50_5;

wire[27:0] addr_50_5;

Selector_2 s50_5(wires_12_4[2], addr_12_4, wires_50_5,addr_50_5);

wire[3:0] wires_51_5;

wire[27:0] addr_51_5;

Selector_2 s51_5(wires_12_4[3], addr_12_4, wires_51_5,addr_51_5);

wire[3:0] wires_52_5;

wire[27:0] addr_52_5;

Selector_2 s52_5(wires_13_4[0], addr_13_4, wires_52_5,addr_52_5);

wire[3:0] wires_53_5;

wire[27:0] addr_53_5;

Selector_2 s53_5(wires_13_4[1], addr_13_4, wires_53_5,addr_53_5);

wire[3:0] wires_54_5;

wire[27:0] addr_54_5;

Selector_2 s54_5(wires_13_4[2], addr_13_4, wires_54_5,addr_54_5);

wire[3:0] wires_55_5;

wire[27:0] addr_55_5;

Selector_2 s55_5(wires_13_4[3], addr_13_4, wires_55_5,addr_55_5);

wire[3:0] wires_56_5;

wire[27:0] addr_56_5;

Selector_2 s56_5(wires_14_4[0], addr_14_4, wires_56_5,addr_56_5);

wire[3:0] wires_57_5;

wire[27:0] addr_57_5;

Selector_2 s57_5(wires_14_4[1], addr_14_4, wires_57_5,addr_57_5);

wire[3:0] wires_58_5;

wire[27:0] addr_58_5;

Selector_2 s58_5(wires_14_4[2], addr_14_4, wires_58_5,addr_58_5);

wire[3:0] wires_59_5;

wire[27:0] addr_59_5;

Selector_2 s59_5(wires_14_4[3], addr_14_4, wires_59_5,addr_59_5);

wire[3:0] wires_60_5;

wire[27:0] addr_60_5;

Selector_2 s60_5(wires_15_4[0], addr_15_4, wires_60_5,addr_60_5);

wire[3:0] wires_61_5;

wire[27:0] addr_61_5;

Selector_2 s61_5(wires_15_4[1], addr_15_4, wires_61_5,addr_61_5);

wire[3:0] wires_62_5;

wire[27:0] addr_62_5;

Selector_2 s62_5(wires_15_4[2], addr_15_4, wires_62_5,addr_62_5);

wire[3:0] wires_63_5;

wire[27:0] addr_63_5;

Selector_2 s63_5(wires_15_4[3], addr_15_4, wires_63_5,addr_63_5);

wire[3:0] wires_64_5;

wire[27:0] addr_64_5;

Selector_2 s64_5(wires_16_4[0], addr_16_4, wires_64_5,addr_64_5);

wire[3:0] wires_65_5;

wire[27:0] addr_65_5;

Selector_2 s65_5(wires_16_4[1], addr_16_4, wires_65_5,addr_65_5);

wire[3:0] wires_66_5;

wire[27:0] addr_66_5;

Selector_2 s66_5(wires_16_4[2], addr_16_4, wires_66_5,addr_66_5);

wire[3:0] wires_67_5;

wire[27:0] addr_67_5;

Selector_2 s67_5(wires_16_4[3], addr_16_4, wires_67_5,addr_67_5);

wire[3:0] wires_68_5;

wire[27:0] addr_68_5;

Selector_2 s68_5(wires_17_4[0], addr_17_4, wires_68_5,addr_68_5);

wire[3:0] wires_69_5;

wire[27:0] addr_69_5;

Selector_2 s69_5(wires_17_4[1], addr_17_4, wires_69_5,addr_69_5);

wire[3:0] wires_70_5;

wire[27:0] addr_70_5;

Selector_2 s70_5(wires_17_4[2], addr_17_4, wires_70_5,addr_70_5);

wire[3:0] wires_71_5;

wire[27:0] addr_71_5;

Selector_2 s71_5(wires_17_4[3], addr_17_4, wires_71_5,addr_71_5);

wire[3:0] wires_72_5;

wire[27:0] addr_72_5;

Selector_2 s72_5(wires_18_4[0], addr_18_4, wires_72_5,addr_72_5);

wire[3:0] wires_73_5;

wire[27:0] addr_73_5;

Selector_2 s73_5(wires_18_4[1], addr_18_4, wires_73_5,addr_73_5);

wire[3:0] wires_74_5;

wire[27:0] addr_74_5;

Selector_2 s74_5(wires_18_4[2], addr_18_4, wires_74_5,addr_74_5);

wire[3:0] wires_75_5;

wire[27:0] addr_75_5;

Selector_2 s75_5(wires_18_4[3], addr_18_4, wires_75_5,addr_75_5);

wire[3:0] wires_76_5;

wire[27:0] addr_76_5;

Selector_2 s76_5(wires_19_4[0], addr_19_4, wires_76_5,addr_76_5);

wire[3:0] wires_77_5;

wire[27:0] addr_77_5;

Selector_2 s77_5(wires_19_4[1], addr_19_4, wires_77_5,addr_77_5);

wire[3:0] wires_78_5;

wire[27:0] addr_78_5;

Selector_2 s78_5(wires_19_4[2], addr_19_4, wires_78_5,addr_78_5);

wire[3:0] wires_79_5;

wire[27:0] addr_79_5;

Selector_2 s79_5(wires_19_4[3], addr_19_4, wires_79_5,addr_79_5);

wire[3:0] wires_80_5;

wire[27:0] addr_80_5;

Selector_2 s80_5(wires_20_4[0], addr_20_4, wires_80_5,addr_80_5);

wire[3:0] wires_81_5;

wire[27:0] addr_81_5;

Selector_2 s81_5(wires_20_4[1], addr_20_4, wires_81_5,addr_81_5);

wire[3:0] wires_82_5;

wire[27:0] addr_82_5;

Selector_2 s82_5(wires_20_4[2], addr_20_4, wires_82_5,addr_82_5);

wire[3:0] wires_83_5;

wire[27:0] addr_83_5;

Selector_2 s83_5(wires_20_4[3], addr_20_4, wires_83_5,addr_83_5);

wire[3:0] wires_84_5;

wire[27:0] addr_84_5;

Selector_2 s84_5(wires_21_4[0], addr_21_4, wires_84_5,addr_84_5);

wire[3:0] wires_85_5;

wire[27:0] addr_85_5;

Selector_2 s85_5(wires_21_4[1], addr_21_4, wires_85_5,addr_85_5);

wire[3:0] wires_86_5;

wire[27:0] addr_86_5;

Selector_2 s86_5(wires_21_4[2], addr_21_4, wires_86_5,addr_86_5);

wire[3:0] wires_87_5;

wire[27:0] addr_87_5;

Selector_2 s87_5(wires_21_4[3], addr_21_4, wires_87_5,addr_87_5);

wire[3:0] wires_88_5;

wire[27:0] addr_88_5;

Selector_2 s88_5(wires_22_4[0], addr_22_4, wires_88_5,addr_88_5);

wire[3:0] wires_89_5;

wire[27:0] addr_89_5;

Selector_2 s89_5(wires_22_4[1], addr_22_4, wires_89_5,addr_89_5);

wire[3:0] wires_90_5;

wire[27:0] addr_90_5;

Selector_2 s90_5(wires_22_4[2], addr_22_4, wires_90_5,addr_90_5);

wire[3:0] wires_91_5;

wire[27:0] addr_91_5;

Selector_2 s91_5(wires_22_4[3], addr_22_4, wires_91_5,addr_91_5);

wire[3:0] wires_92_5;

wire[27:0] addr_92_5;

Selector_2 s92_5(wires_23_4[0], addr_23_4, wires_92_5,addr_92_5);

wire[3:0] wires_93_5;

wire[27:0] addr_93_5;

Selector_2 s93_5(wires_23_4[1], addr_23_4, wires_93_5,addr_93_5);

wire[3:0] wires_94_5;

wire[27:0] addr_94_5;

Selector_2 s94_5(wires_23_4[2], addr_23_4, wires_94_5,addr_94_5);

wire[3:0] wires_95_5;

wire[27:0] addr_95_5;

Selector_2 s95_5(wires_23_4[3], addr_23_4, wires_95_5,addr_95_5);

wire[3:0] wires_96_5;

wire[27:0] addr_96_5;

Selector_2 s96_5(wires_24_4[0], addr_24_4, wires_96_5,addr_96_5);

wire[3:0] wires_97_5;

wire[27:0] addr_97_5;

Selector_2 s97_5(wires_24_4[1], addr_24_4, wires_97_5,addr_97_5);

wire[3:0] wires_98_5;

wire[27:0] addr_98_5;

Selector_2 s98_5(wires_24_4[2], addr_24_4, wires_98_5,addr_98_5);

wire[3:0] wires_99_5;

wire[27:0] addr_99_5;

Selector_2 s99_5(wires_24_4[3], addr_24_4, wires_99_5,addr_99_5);

wire[3:0] wires_100_5;

wire[27:0] addr_100_5;

Selector_2 s100_5(wires_25_4[0], addr_25_4, wires_100_5,addr_100_5);

wire[3:0] wires_101_5;

wire[27:0] addr_101_5;

Selector_2 s101_5(wires_25_4[1], addr_25_4, wires_101_5,addr_101_5);

wire[3:0] wires_102_5;

wire[27:0] addr_102_5;

Selector_2 s102_5(wires_25_4[2], addr_25_4, wires_102_5,addr_102_5);

wire[3:0] wires_103_5;

wire[27:0] addr_103_5;

Selector_2 s103_5(wires_25_4[3], addr_25_4, wires_103_5,addr_103_5);

wire[3:0] wires_104_5;

wire[27:0] addr_104_5;

Selector_2 s104_5(wires_26_4[0], addr_26_4, wires_104_5,addr_104_5);

wire[3:0] wires_105_5;

wire[27:0] addr_105_5;

Selector_2 s105_5(wires_26_4[1], addr_26_4, wires_105_5,addr_105_5);

wire[3:0] wires_106_5;

wire[27:0] addr_106_5;

Selector_2 s106_5(wires_26_4[2], addr_26_4, wires_106_5,addr_106_5);

wire[3:0] wires_107_5;

wire[27:0] addr_107_5;

Selector_2 s107_5(wires_26_4[3], addr_26_4, wires_107_5,addr_107_5);

wire[3:0] wires_108_5;

wire[27:0] addr_108_5;

Selector_2 s108_5(wires_27_4[0], addr_27_4, wires_108_5,addr_108_5);

wire[3:0] wires_109_5;

wire[27:0] addr_109_5;

Selector_2 s109_5(wires_27_4[1], addr_27_4, wires_109_5,addr_109_5);

wire[3:0] wires_110_5;

wire[27:0] addr_110_5;

Selector_2 s110_5(wires_27_4[2], addr_27_4, wires_110_5,addr_110_5);

wire[3:0] wires_111_5;

wire[27:0] addr_111_5;

Selector_2 s111_5(wires_27_4[3], addr_27_4, wires_111_5,addr_111_5);

wire[3:0] wires_112_5;

wire[27:0] addr_112_5;

Selector_2 s112_5(wires_28_4[0], addr_28_4, wires_112_5,addr_112_5);

wire[3:0] wires_113_5;

wire[27:0] addr_113_5;

Selector_2 s113_5(wires_28_4[1], addr_28_4, wires_113_5,addr_113_5);

wire[3:0] wires_114_5;

wire[27:0] addr_114_5;

Selector_2 s114_5(wires_28_4[2], addr_28_4, wires_114_5,addr_114_5);

wire[3:0] wires_115_5;

wire[27:0] addr_115_5;

Selector_2 s115_5(wires_28_4[3], addr_28_4, wires_115_5,addr_115_5);

wire[3:0] wires_116_5;

wire[27:0] addr_116_5;

Selector_2 s116_5(wires_29_4[0], addr_29_4, wires_116_5,addr_116_5);

wire[3:0] wires_117_5;

wire[27:0] addr_117_5;

Selector_2 s117_5(wires_29_4[1], addr_29_4, wires_117_5,addr_117_5);

wire[3:0] wires_118_5;

wire[27:0] addr_118_5;

Selector_2 s118_5(wires_29_4[2], addr_29_4, wires_118_5,addr_118_5);

wire[3:0] wires_119_5;

wire[27:0] addr_119_5;

Selector_2 s119_5(wires_29_4[3], addr_29_4, wires_119_5,addr_119_5);

wire[3:0] wires_120_5;

wire[27:0] addr_120_5;

Selector_2 s120_5(wires_30_4[0], addr_30_4, wires_120_5,addr_120_5);

wire[3:0] wires_121_5;

wire[27:0] addr_121_5;

Selector_2 s121_5(wires_30_4[1], addr_30_4, wires_121_5,addr_121_5);

wire[3:0] wires_122_5;

wire[27:0] addr_122_5;

Selector_2 s122_5(wires_30_4[2], addr_30_4, wires_122_5,addr_122_5);

wire[3:0] wires_123_5;

wire[27:0] addr_123_5;

Selector_2 s123_5(wires_30_4[3], addr_30_4, wires_123_5,addr_123_5);

wire[3:0] wires_124_5;

wire[27:0] addr_124_5;

Selector_2 s124_5(wires_31_4[0], addr_31_4, wires_124_5,addr_124_5);

wire[3:0] wires_125_5;

wire[27:0] addr_125_5;

Selector_2 s125_5(wires_31_4[1], addr_31_4, wires_125_5,addr_125_5);

wire[3:0] wires_126_5;

wire[27:0] addr_126_5;

Selector_2 s126_5(wires_31_4[2], addr_31_4, wires_126_5,addr_126_5);

wire[3:0] wires_127_5;

wire[27:0] addr_127_5;

Selector_2 s127_5(wires_31_4[3], addr_31_4, wires_127_5,addr_127_5);

wire[3:0] wires_128_5;

wire[27:0] addr_128_5;

Selector_2 s128_5(wires_32_4[0], addr_32_4, wires_128_5,addr_128_5);

wire[3:0] wires_129_5;

wire[27:0] addr_129_5;

Selector_2 s129_5(wires_32_4[1], addr_32_4, wires_129_5,addr_129_5);

wire[3:0] wires_130_5;

wire[27:0] addr_130_5;

Selector_2 s130_5(wires_32_4[2], addr_32_4, wires_130_5,addr_130_5);

wire[3:0] wires_131_5;

wire[27:0] addr_131_5;

Selector_2 s131_5(wires_32_4[3], addr_32_4, wires_131_5,addr_131_5);

wire[3:0] wires_132_5;

wire[27:0] addr_132_5;

Selector_2 s132_5(wires_33_4[0], addr_33_4, wires_132_5,addr_132_5);

wire[3:0] wires_133_5;

wire[27:0] addr_133_5;

Selector_2 s133_5(wires_33_4[1], addr_33_4, wires_133_5,addr_133_5);

wire[3:0] wires_134_5;

wire[27:0] addr_134_5;

Selector_2 s134_5(wires_33_4[2], addr_33_4, wires_134_5,addr_134_5);

wire[3:0] wires_135_5;

wire[27:0] addr_135_5;

Selector_2 s135_5(wires_33_4[3], addr_33_4, wires_135_5,addr_135_5);

wire[3:0] wires_136_5;

wire[27:0] addr_136_5;

Selector_2 s136_5(wires_34_4[0], addr_34_4, wires_136_5,addr_136_5);

wire[3:0] wires_137_5;

wire[27:0] addr_137_5;

Selector_2 s137_5(wires_34_4[1], addr_34_4, wires_137_5,addr_137_5);

wire[3:0] wires_138_5;

wire[27:0] addr_138_5;

Selector_2 s138_5(wires_34_4[2], addr_34_4, wires_138_5,addr_138_5);

wire[3:0] wires_139_5;

wire[27:0] addr_139_5;

Selector_2 s139_5(wires_34_4[3], addr_34_4, wires_139_5,addr_139_5);

wire[3:0] wires_140_5;

wire[27:0] addr_140_5;

Selector_2 s140_5(wires_35_4[0], addr_35_4, wires_140_5,addr_140_5);

wire[3:0] wires_141_5;

wire[27:0] addr_141_5;

Selector_2 s141_5(wires_35_4[1], addr_35_4, wires_141_5,addr_141_5);

wire[3:0] wires_142_5;

wire[27:0] addr_142_5;

Selector_2 s142_5(wires_35_4[2], addr_35_4, wires_142_5,addr_142_5);

wire[3:0] wires_143_5;

wire[27:0] addr_143_5;

Selector_2 s143_5(wires_35_4[3], addr_35_4, wires_143_5,addr_143_5);

wire[3:0] wires_144_5;

wire[27:0] addr_144_5;

Selector_2 s144_5(wires_36_4[0], addr_36_4, wires_144_5,addr_144_5);

wire[3:0] wires_145_5;

wire[27:0] addr_145_5;

Selector_2 s145_5(wires_36_4[1], addr_36_4, wires_145_5,addr_145_5);

wire[3:0] wires_146_5;

wire[27:0] addr_146_5;

Selector_2 s146_5(wires_36_4[2], addr_36_4, wires_146_5,addr_146_5);

wire[3:0] wires_147_5;

wire[27:0] addr_147_5;

Selector_2 s147_5(wires_36_4[3], addr_36_4, wires_147_5,addr_147_5);

wire[3:0] wires_148_5;

wire[27:0] addr_148_5;

Selector_2 s148_5(wires_37_4[0], addr_37_4, wires_148_5,addr_148_5);

wire[3:0] wires_149_5;

wire[27:0] addr_149_5;

Selector_2 s149_5(wires_37_4[1], addr_37_4, wires_149_5,addr_149_5);

wire[3:0] wires_150_5;

wire[27:0] addr_150_5;

Selector_2 s150_5(wires_37_4[2], addr_37_4, wires_150_5,addr_150_5);

wire[3:0] wires_151_5;

wire[27:0] addr_151_5;

Selector_2 s151_5(wires_37_4[3], addr_37_4, wires_151_5,addr_151_5);

wire[3:0] wires_152_5;

wire[27:0] addr_152_5;

Selector_2 s152_5(wires_38_4[0], addr_38_4, wires_152_5,addr_152_5);

wire[3:0] wires_153_5;

wire[27:0] addr_153_5;

Selector_2 s153_5(wires_38_4[1], addr_38_4, wires_153_5,addr_153_5);

wire[3:0] wires_154_5;

wire[27:0] addr_154_5;

Selector_2 s154_5(wires_38_4[2], addr_38_4, wires_154_5,addr_154_5);

wire[3:0] wires_155_5;

wire[27:0] addr_155_5;

Selector_2 s155_5(wires_38_4[3], addr_38_4, wires_155_5,addr_155_5);

wire[3:0] wires_156_5;

wire[27:0] addr_156_5;

Selector_2 s156_5(wires_39_4[0], addr_39_4, wires_156_5,addr_156_5);

wire[3:0] wires_157_5;

wire[27:0] addr_157_5;

Selector_2 s157_5(wires_39_4[1], addr_39_4, wires_157_5,addr_157_5);

wire[3:0] wires_158_5;

wire[27:0] addr_158_5;

Selector_2 s158_5(wires_39_4[2], addr_39_4, wires_158_5,addr_158_5);

wire[3:0] wires_159_5;

wire[27:0] addr_159_5;

Selector_2 s159_5(wires_39_4[3], addr_39_4, wires_159_5,addr_159_5);

wire[3:0] wires_160_5;

wire[27:0] addr_160_5;

Selector_2 s160_5(wires_40_4[0], addr_40_4, wires_160_5,addr_160_5);

wire[3:0] wires_161_5;

wire[27:0] addr_161_5;

Selector_2 s161_5(wires_40_4[1], addr_40_4, wires_161_5,addr_161_5);

wire[3:0] wires_162_5;

wire[27:0] addr_162_5;

Selector_2 s162_5(wires_40_4[2], addr_40_4, wires_162_5,addr_162_5);

wire[3:0] wires_163_5;

wire[27:0] addr_163_5;

Selector_2 s163_5(wires_40_4[3], addr_40_4, wires_163_5,addr_163_5);

wire[3:0] wires_164_5;

wire[27:0] addr_164_5;

Selector_2 s164_5(wires_41_4[0], addr_41_4, wires_164_5,addr_164_5);

wire[3:0] wires_165_5;

wire[27:0] addr_165_5;

Selector_2 s165_5(wires_41_4[1], addr_41_4, wires_165_5,addr_165_5);

wire[3:0] wires_166_5;

wire[27:0] addr_166_5;

Selector_2 s166_5(wires_41_4[2], addr_41_4, wires_166_5,addr_166_5);

wire[3:0] wires_167_5;

wire[27:0] addr_167_5;

Selector_2 s167_5(wires_41_4[3], addr_41_4, wires_167_5,addr_167_5);

wire[3:0] wires_168_5;

wire[27:0] addr_168_5;

Selector_2 s168_5(wires_42_4[0], addr_42_4, wires_168_5,addr_168_5);

wire[3:0] wires_169_5;

wire[27:0] addr_169_5;

Selector_2 s169_5(wires_42_4[1], addr_42_4, wires_169_5,addr_169_5);

wire[3:0] wires_170_5;

wire[27:0] addr_170_5;

Selector_2 s170_5(wires_42_4[2], addr_42_4, wires_170_5,addr_170_5);

wire[3:0] wires_171_5;

wire[27:0] addr_171_5;

Selector_2 s171_5(wires_42_4[3], addr_42_4, wires_171_5,addr_171_5);

wire[3:0] wires_172_5;

wire[27:0] addr_172_5;

Selector_2 s172_5(wires_43_4[0], addr_43_4, wires_172_5,addr_172_5);

wire[3:0] wires_173_5;

wire[27:0] addr_173_5;

Selector_2 s173_5(wires_43_4[1], addr_43_4, wires_173_5,addr_173_5);

wire[3:0] wires_174_5;

wire[27:0] addr_174_5;

Selector_2 s174_5(wires_43_4[2], addr_43_4, wires_174_5,addr_174_5);

wire[3:0] wires_175_5;

wire[27:0] addr_175_5;

Selector_2 s175_5(wires_43_4[3], addr_43_4, wires_175_5,addr_175_5);

wire[3:0] wires_176_5;

wire[27:0] addr_176_5;

Selector_2 s176_5(wires_44_4[0], addr_44_4, wires_176_5,addr_176_5);

wire[3:0] wires_177_5;

wire[27:0] addr_177_5;

Selector_2 s177_5(wires_44_4[1], addr_44_4, wires_177_5,addr_177_5);

wire[3:0] wires_178_5;

wire[27:0] addr_178_5;

Selector_2 s178_5(wires_44_4[2], addr_44_4, wires_178_5,addr_178_5);

wire[3:0] wires_179_5;

wire[27:0] addr_179_5;

Selector_2 s179_5(wires_44_4[3], addr_44_4, wires_179_5,addr_179_5);

wire[3:0] wires_180_5;

wire[27:0] addr_180_5;

Selector_2 s180_5(wires_45_4[0], addr_45_4, wires_180_5,addr_180_5);

wire[3:0] wires_181_5;

wire[27:0] addr_181_5;

Selector_2 s181_5(wires_45_4[1], addr_45_4, wires_181_5,addr_181_5);

wire[3:0] wires_182_5;

wire[27:0] addr_182_5;

Selector_2 s182_5(wires_45_4[2], addr_45_4, wires_182_5,addr_182_5);

wire[3:0] wires_183_5;

wire[27:0] addr_183_5;

Selector_2 s183_5(wires_45_4[3], addr_45_4, wires_183_5,addr_183_5);

wire[3:0] wires_184_5;

wire[27:0] addr_184_5;

Selector_2 s184_5(wires_46_4[0], addr_46_4, wires_184_5,addr_184_5);

wire[3:0] wires_185_5;

wire[27:0] addr_185_5;

Selector_2 s185_5(wires_46_4[1], addr_46_4, wires_185_5,addr_185_5);

wire[3:0] wires_186_5;

wire[27:0] addr_186_5;

Selector_2 s186_5(wires_46_4[2], addr_46_4, wires_186_5,addr_186_5);

wire[3:0] wires_187_5;

wire[27:0] addr_187_5;

Selector_2 s187_5(wires_46_4[3], addr_46_4, wires_187_5,addr_187_5);

wire[3:0] wires_188_5;

wire[27:0] addr_188_5;

Selector_2 s188_5(wires_47_4[0], addr_47_4, wires_188_5,addr_188_5);

wire[3:0] wires_189_5;

wire[27:0] addr_189_5;

Selector_2 s189_5(wires_47_4[1], addr_47_4, wires_189_5,addr_189_5);

wire[3:0] wires_190_5;

wire[27:0] addr_190_5;

Selector_2 s190_5(wires_47_4[2], addr_47_4, wires_190_5,addr_190_5);

wire[3:0] wires_191_5;

wire[27:0] addr_191_5;

Selector_2 s191_5(wires_47_4[3], addr_47_4, wires_191_5,addr_191_5);

wire[3:0] wires_192_5;

wire[27:0] addr_192_5;

Selector_2 s192_5(wires_48_4[0], addr_48_4, wires_192_5,addr_192_5);

wire[3:0] wires_193_5;

wire[27:0] addr_193_5;

Selector_2 s193_5(wires_48_4[1], addr_48_4, wires_193_5,addr_193_5);

wire[3:0] wires_194_5;

wire[27:0] addr_194_5;

Selector_2 s194_5(wires_48_4[2], addr_48_4, wires_194_5,addr_194_5);

wire[3:0] wires_195_5;

wire[27:0] addr_195_5;

Selector_2 s195_5(wires_48_4[3], addr_48_4, wires_195_5,addr_195_5);

wire[3:0] wires_196_5;

wire[27:0] addr_196_5;

Selector_2 s196_5(wires_49_4[0], addr_49_4, wires_196_5,addr_196_5);

wire[3:0] wires_197_5;

wire[27:0] addr_197_5;

Selector_2 s197_5(wires_49_4[1], addr_49_4, wires_197_5,addr_197_5);

wire[3:0] wires_198_5;

wire[27:0] addr_198_5;

Selector_2 s198_5(wires_49_4[2], addr_49_4, wires_198_5,addr_198_5);

wire[3:0] wires_199_5;

wire[27:0] addr_199_5;

Selector_2 s199_5(wires_49_4[3], addr_49_4, wires_199_5,addr_199_5);

wire[3:0] wires_200_5;

wire[27:0] addr_200_5;

Selector_2 s200_5(wires_50_4[0], addr_50_4, wires_200_5,addr_200_5);

wire[3:0] wires_201_5;

wire[27:0] addr_201_5;

Selector_2 s201_5(wires_50_4[1], addr_50_4, wires_201_5,addr_201_5);

wire[3:0] wires_202_5;

wire[27:0] addr_202_5;

Selector_2 s202_5(wires_50_4[2], addr_50_4, wires_202_5,addr_202_5);

wire[3:0] wires_203_5;

wire[27:0] addr_203_5;

Selector_2 s203_5(wires_50_4[3], addr_50_4, wires_203_5,addr_203_5);

wire[3:0] wires_204_5;

wire[27:0] addr_204_5;

Selector_2 s204_5(wires_51_4[0], addr_51_4, wires_204_5,addr_204_5);

wire[3:0] wires_205_5;

wire[27:0] addr_205_5;

Selector_2 s205_5(wires_51_4[1], addr_51_4, wires_205_5,addr_205_5);

wire[3:0] wires_206_5;

wire[27:0] addr_206_5;

Selector_2 s206_5(wires_51_4[2], addr_51_4, wires_206_5,addr_206_5);

wire[3:0] wires_207_5;

wire[27:0] addr_207_5;

Selector_2 s207_5(wires_51_4[3], addr_51_4, wires_207_5,addr_207_5);

wire[3:0] wires_208_5;

wire[27:0] addr_208_5;

Selector_2 s208_5(wires_52_4[0], addr_52_4, wires_208_5,addr_208_5);

wire[3:0] wires_209_5;

wire[27:0] addr_209_5;

Selector_2 s209_5(wires_52_4[1], addr_52_4, wires_209_5,addr_209_5);

wire[3:0] wires_210_5;

wire[27:0] addr_210_5;

Selector_2 s210_5(wires_52_4[2], addr_52_4, wires_210_5,addr_210_5);

wire[3:0] wires_211_5;

wire[27:0] addr_211_5;

Selector_2 s211_5(wires_52_4[3], addr_52_4, wires_211_5,addr_211_5);

wire[3:0] wires_212_5;

wire[27:0] addr_212_5;

Selector_2 s212_5(wires_53_4[0], addr_53_4, wires_212_5,addr_212_5);

wire[3:0] wires_213_5;

wire[27:0] addr_213_5;

Selector_2 s213_5(wires_53_4[1], addr_53_4, wires_213_5,addr_213_5);

wire[3:0] wires_214_5;

wire[27:0] addr_214_5;

Selector_2 s214_5(wires_53_4[2], addr_53_4, wires_214_5,addr_214_5);

wire[3:0] wires_215_5;

wire[27:0] addr_215_5;

Selector_2 s215_5(wires_53_4[3], addr_53_4, wires_215_5,addr_215_5);

wire[3:0] wires_216_5;

wire[27:0] addr_216_5;

Selector_2 s216_5(wires_54_4[0], addr_54_4, wires_216_5,addr_216_5);

wire[3:0] wires_217_5;

wire[27:0] addr_217_5;

Selector_2 s217_5(wires_54_4[1], addr_54_4, wires_217_5,addr_217_5);

wire[3:0] wires_218_5;

wire[27:0] addr_218_5;

Selector_2 s218_5(wires_54_4[2], addr_54_4, wires_218_5,addr_218_5);

wire[3:0] wires_219_5;

wire[27:0] addr_219_5;

Selector_2 s219_5(wires_54_4[3], addr_54_4, wires_219_5,addr_219_5);

wire[3:0] wires_220_5;

wire[27:0] addr_220_5;

Selector_2 s220_5(wires_55_4[0], addr_55_4, wires_220_5,addr_220_5);

wire[3:0] wires_221_5;

wire[27:0] addr_221_5;

Selector_2 s221_5(wires_55_4[1], addr_55_4, wires_221_5,addr_221_5);

wire[3:0] wires_222_5;

wire[27:0] addr_222_5;

Selector_2 s222_5(wires_55_4[2], addr_55_4, wires_222_5,addr_222_5);

wire[3:0] wires_223_5;

wire[27:0] addr_223_5;

Selector_2 s223_5(wires_55_4[3], addr_55_4, wires_223_5,addr_223_5);

wire[3:0] wires_224_5;

wire[27:0] addr_224_5;

Selector_2 s224_5(wires_56_4[0], addr_56_4, wires_224_5,addr_224_5);

wire[3:0] wires_225_5;

wire[27:0] addr_225_5;

Selector_2 s225_5(wires_56_4[1], addr_56_4, wires_225_5,addr_225_5);

wire[3:0] wires_226_5;

wire[27:0] addr_226_5;

Selector_2 s226_5(wires_56_4[2], addr_56_4, wires_226_5,addr_226_5);

wire[3:0] wires_227_5;

wire[27:0] addr_227_5;

Selector_2 s227_5(wires_56_4[3], addr_56_4, wires_227_5,addr_227_5);

wire[3:0] wires_228_5;

wire[27:0] addr_228_5;

Selector_2 s228_5(wires_57_4[0], addr_57_4, wires_228_5,addr_228_5);

wire[3:0] wires_229_5;

wire[27:0] addr_229_5;

Selector_2 s229_5(wires_57_4[1], addr_57_4, wires_229_5,addr_229_5);

wire[3:0] wires_230_5;

wire[27:0] addr_230_5;

Selector_2 s230_5(wires_57_4[2], addr_57_4, wires_230_5,addr_230_5);

wire[3:0] wires_231_5;

wire[27:0] addr_231_5;

Selector_2 s231_5(wires_57_4[3], addr_57_4, wires_231_5,addr_231_5);

wire[3:0] wires_232_5;

wire[27:0] addr_232_5;

Selector_2 s232_5(wires_58_4[0], addr_58_4, wires_232_5,addr_232_5);

wire[3:0] wires_233_5;

wire[27:0] addr_233_5;

Selector_2 s233_5(wires_58_4[1], addr_58_4, wires_233_5,addr_233_5);

wire[3:0] wires_234_5;

wire[27:0] addr_234_5;

Selector_2 s234_5(wires_58_4[2], addr_58_4, wires_234_5,addr_234_5);

wire[3:0] wires_235_5;

wire[27:0] addr_235_5;

Selector_2 s235_5(wires_58_4[3], addr_58_4, wires_235_5,addr_235_5);

wire[3:0] wires_236_5;

wire[27:0] addr_236_5;

Selector_2 s236_5(wires_59_4[0], addr_59_4, wires_236_5,addr_236_5);

wire[3:0] wires_237_5;

wire[27:0] addr_237_5;

Selector_2 s237_5(wires_59_4[1], addr_59_4, wires_237_5,addr_237_5);

wire[3:0] wires_238_5;

wire[27:0] addr_238_5;

Selector_2 s238_5(wires_59_4[2], addr_59_4, wires_238_5,addr_238_5);

wire[3:0] wires_239_5;

wire[27:0] addr_239_5;

Selector_2 s239_5(wires_59_4[3], addr_59_4, wires_239_5,addr_239_5);

wire[3:0] wires_240_5;

wire[27:0] addr_240_5;

Selector_2 s240_5(wires_60_4[0], addr_60_4, wires_240_5,addr_240_5);

wire[3:0] wires_241_5;

wire[27:0] addr_241_5;

Selector_2 s241_5(wires_60_4[1], addr_60_4, wires_241_5,addr_241_5);

wire[3:0] wires_242_5;

wire[27:0] addr_242_5;

Selector_2 s242_5(wires_60_4[2], addr_60_4, wires_242_5,addr_242_5);

wire[3:0] wires_243_5;

wire[27:0] addr_243_5;

Selector_2 s243_5(wires_60_4[3], addr_60_4, wires_243_5,addr_243_5);

wire[3:0] wires_244_5;

wire[27:0] addr_244_5;

Selector_2 s244_5(wires_61_4[0], addr_61_4, wires_244_5,addr_244_5);

wire[3:0] wires_245_5;

wire[27:0] addr_245_5;

Selector_2 s245_5(wires_61_4[1], addr_61_4, wires_245_5,addr_245_5);

wire[3:0] wires_246_5;

wire[27:0] addr_246_5;

Selector_2 s246_5(wires_61_4[2], addr_61_4, wires_246_5,addr_246_5);

wire[3:0] wires_247_5;

wire[27:0] addr_247_5;

Selector_2 s247_5(wires_61_4[3], addr_61_4, wires_247_5,addr_247_5);

wire[3:0] wires_248_5;

wire[27:0] addr_248_5;

Selector_2 s248_5(wires_62_4[0], addr_62_4, wires_248_5,addr_248_5);

wire[3:0] wires_249_5;

wire[27:0] addr_249_5;

Selector_2 s249_5(wires_62_4[1], addr_62_4, wires_249_5,addr_249_5);

wire[3:0] wires_250_5;

wire[27:0] addr_250_5;

Selector_2 s250_5(wires_62_4[2], addr_62_4, wires_250_5,addr_250_5);

wire[3:0] wires_251_5;

wire[27:0] addr_251_5;

Selector_2 s251_5(wires_62_4[3], addr_62_4, wires_251_5,addr_251_5);

wire[3:0] wires_252_5;

wire[27:0] addr_252_5;

Selector_2 s252_5(wires_63_4[0], addr_63_4, wires_252_5,addr_252_5);

wire[3:0] wires_253_5;

wire[27:0] addr_253_5;

Selector_2 s253_5(wires_63_4[1], addr_63_4, wires_253_5,addr_253_5);

wire[3:0] wires_254_5;

wire[27:0] addr_254_5;

Selector_2 s254_5(wires_63_4[2], addr_63_4, wires_254_5,addr_254_5);

wire[3:0] wires_255_5;

wire[27:0] addr_255_5;

Selector_2 s255_5(wires_63_4[3], addr_63_4, wires_255_5,addr_255_5);

wire[3:0] wires_256_5;

wire[27:0] addr_256_5;

Selector_2 s256_5(wires_64_4[0], addr_64_4, wires_256_5,addr_256_5);

wire[3:0] wires_257_5;

wire[27:0] addr_257_5;

Selector_2 s257_5(wires_64_4[1], addr_64_4, wires_257_5,addr_257_5);

wire[3:0] wires_258_5;

wire[27:0] addr_258_5;

Selector_2 s258_5(wires_64_4[2], addr_64_4, wires_258_5,addr_258_5);

wire[3:0] wires_259_5;

wire[27:0] addr_259_5;

Selector_2 s259_5(wires_64_4[3], addr_64_4, wires_259_5,addr_259_5);

wire[3:0] wires_260_5;

wire[27:0] addr_260_5;

Selector_2 s260_5(wires_65_4[0], addr_65_4, wires_260_5,addr_260_5);

wire[3:0] wires_261_5;

wire[27:0] addr_261_5;

Selector_2 s261_5(wires_65_4[1], addr_65_4, wires_261_5,addr_261_5);

wire[3:0] wires_262_5;

wire[27:0] addr_262_5;

Selector_2 s262_5(wires_65_4[2], addr_65_4, wires_262_5,addr_262_5);

wire[3:0] wires_263_5;

wire[27:0] addr_263_5;

Selector_2 s263_5(wires_65_4[3], addr_65_4, wires_263_5,addr_263_5);

wire[3:0] wires_264_5;

wire[27:0] addr_264_5;

Selector_2 s264_5(wires_66_4[0], addr_66_4, wires_264_5,addr_264_5);

wire[3:0] wires_265_5;

wire[27:0] addr_265_5;

Selector_2 s265_5(wires_66_4[1], addr_66_4, wires_265_5,addr_265_5);

wire[3:0] wires_266_5;

wire[27:0] addr_266_5;

Selector_2 s266_5(wires_66_4[2], addr_66_4, wires_266_5,addr_266_5);

wire[3:0] wires_267_5;

wire[27:0] addr_267_5;

Selector_2 s267_5(wires_66_4[3], addr_66_4, wires_267_5,addr_267_5);

wire[3:0] wires_268_5;

wire[27:0] addr_268_5;

Selector_2 s268_5(wires_67_4[0], addr_67_4, wires_268_5,addr_268_5);

wire[3:0] wires_269_5;

wire[27:0] addr_269_5;

Selector_2 s269_5(wires_67_4[1], addr_67_4, wires_269_5,addr_269_5);

wire[3:0] wires_270_5;

wire[27:0] addr_270_5;

Selector_2 s270_5(wires_67_4[2], addr_67_4, wires_270_5,addr_270_5);

wire[3:0] wires_271_5;

wire[27:0] addr_271_5;

Selector_2 s271_5(wires_67_4[3], addr_67_4, wires_271_5,addr_271_5);

wire[3:0] wires_272_5;

wire[27:0] addr_272_5;

Selector_2 s272_5(wires_68_4[0], addr_68_4, wires_272_5,addr_272_5);

wire[3:0] wires_273_5;

wire[27:0] addr_273_5;

Selector_2 s273_5(wires_68_4[1], addr_68_4, wires_273_5,addr_273_5);

wire[3:0] wires_274_5;

wire[27:0] addr_274_5;

Selector_2 s274_5(wires_68_4[2], addr_68_4, wires_274_5,addr_274_5);

wire[3:0] wires_275_5;

wire[27:0] addr_275_5;

Selector_2 s275_5(wires_68_4[3], addr_68_4, wires_275_5,addr_275_5);

wire[3:0] wires_276_5;

wire[27:0] addr_276_5;

Selector_2 s276_5(wires_69_4[0], addr_69_4, wires_276_5,addr_276_5);

wire[3:0] wires_277_5;

wire[27:0] addr_277_5;

Selector_2 s277_5(wires_69_4[1], addr_69_4, wires_277_5,addr_277_5);

wire[3:0] wires_278_5;

wire[27:0] addr_278_5;

Selector_2 s278_5(wires_69_4[2], addr_69_4, wires_278_5,addr_278_5);

wire[3:0] wires_279_5;

wire[27:0] addr_279_5;

Selector_2 s279_5(wires_69_4[3], addr_69_4, wires_279_5,addr_279_5);

wire[3:0] wires_280_5;

wire[27:0] addr_280_5;

Selector_2 s280_5(wires_70_4[0], addr_70_4, wires_280_5,addr_280_5);

wire[3:0] wires_281_5;

wire[27:0] addr_281_5;

Selector_2 s281_5(wires_70_4[1], addr_70_4, wires_281_5,addr_281_5);

wire[3:0] wires_282_5;

wire[27:0] addr_282_5;

Selector_2 s282_5(wires_70_4[2], addr_70_4, wires_282_5,addr_282_5);

wire[3:0] wires_283_5;

wire[27:0] addr_283_5;

Selector_2 s283_5(wires_70_4[3], addr_70_4, wires_283_5,addr_283_5);

wire[3:0] wires_284_5;

wire[27:0] addr_284_5;

Selector_2 s284_5(wires_71_4[0], addr_71_4, wires_284_5,addr_284_5);

wire[3:0] wires_285_5;

wire[27:0] addr_285_5;

Selector_2 s285_5(wires_71_4[1], addr_71_4, wires_285_5,addr_285_5);

wire[3:0] wires_286_5;

wire[27:0] addr_286_5;

Selector_2 s286_5(wires_71_4[2], addr_71_4, wires_286_5,addr_286_5);

wire[3:0] wires_287_5;

wire[27:0] addr_287_5;

Selector_2 s287_5(wires_71_4[3], addr_71_4, wires_287_5,addr_287_5);

wire[3:0] wires_288_5;

wire[27:0] addr_288_5;

Selector_2 s288_5(wires_72_4[0], addr_72_4, wires_288_5,addr_288_5);

wire[3:0] wires_289_5;

wire[27:0] addr_289_5;

Selector_2 s289_5(wires_72_4[1], addr_72_4, wires_289_5,addr_289_5);

wire[3:0] wires_290_5;

wire[27:0] addr_290_5;

Selector_2 s290_5(wires_72_4[2], addr_72_4, wires_290_5,addr_290_5);

wire[3:0] wires_291_5;

wire[27:0] addr_291_5;

Selector_2 s291_5(wires_72_4[3], addr_72_4, wires_291_5,addr_291_5);

wire[3:0] wires_292_5;

wire[27:0] addr_292_5;

Selector_2 s292_5(wires_73_4[0], addr_73_4, wires_292_5,addr_292_5);

wire[3:0] wires_293_5;

wire[27:0] addr_293_5;

Selector_2 s293_5(wires_73_4[1], addr_73_4, wires_293_5,addr_293_5);

wire[3:0] wires_294_5;

wire[27:0] addr_294_5;

Selector_2 s294_5(wires_73_4[2], addr_73_4, wires_294_5,addr_294_5);

wire[3:0] wires_295_5;

wire[27:0] addr_295_5;

Selector_2 s295_5(wires_73_4[3], addr_73_4, wires_295_5,addr_295_5);

wire[3:0] wires_296_5;

wire[27:0] addr_296_5;

Selector_2 s296_5(wires_74_4[0], addr_74_4, wires_296_5,addr_296_5);

wire[3:0] wires_297_5;

wire[27:0] addr_297_5;

Selector_2 s297_5(wires_74_4[1], addr_74_4, wires_297_5,addr_297_5);

wire[3:0] wires_298_5;

wire[27:0] addr_298_5;

Selector_2 s298_5(wires_74_4[2], addr_74_4, wires_298_5,addr_298_5);

wire[3:0] wires_299_5;

wire[27:0] addr_299_5;

Selector_2 s299_5(wires_74_4[3], addr_74_4, wires_299_5,addr_299_5);

wire[3:0] wires_300_5;

wire[27:0] addr_300_5;

Selector_2 s300_5(wires_75_4[0], addr_75_4, wires_300_5,addr_300_5);

wire[3:0] wires_301_5;

wire[27:0] addr_301_5;

Selector_2 s301_5(wires_75_4[1], addr_75_4, wires_301_5,addr_301_5);

wire[3:0] wires_302_5;

wire[27:0] addr_302_5;

Selector_2 s302_5(wires_75_4[2], addr_75_4, wires_302_5,addr_302_5);

wire[3:0] wires_303_5;

wire[27:0] addr_303_5;

Selector_2 s303_5(wires_75_4[3], addr_75_4, wires_303_5,addr_303_5);

wire[3:0] wires_304_5;

wire[27:0] addr_304_5;

Selector_2 s304_5(wires_76_4[0], addr_76_4, wires_304_5,addr_304_5);

wire[3:0] wires_305_5;

wire[27:0] addr_305_5;

Selector_2 s305_5(wires_76_4[1], addr_76_4, wires_305_5,addr_305_5);

wire[3:0] wires_306_5;

wire[27:0] addr_306_5;

Selector_2 s306_5(wires_76_4[2], addr_76_4, wires_306_5,addr_306_5);

wire[3:0] wires_307_5;

wire[27:0] addr_307_5;

Selector_2 s307_5(wires_76_4[3], addr_76_4, wires_307_5,addr_307_5);

wire[3:0] wires_308_5;

wire[27:0] addr_308_5;

Selector_2 s308_5(wires_77_4[0], addr_77_4, wires_308_5,addr_308_5);

wire[3:0] wires_309_5;

wire[27:0] addr_309_5;

Selector_2 s309_5(wires_77_4[1], addr_77_4, wires_309_5,addr_309_5);

wire[3:0] wires_310_5;

wire[27:0] addr_310_5;

Selector_2 s310_5(wires_77_4[2], addr_77_4, wires_310_5,addr_310_5);

wire[3:0] wires_311_5;

wire[27:0] addr_311_5;

Selector_2 s311_5(wires_77_4[3], addr_77_4, wires_311_5,addr_311_5);

wire[3:0] wires_312_5;

wire[27:0] addr_312_5;

Selector_2 s312_5(wires_78_4[0], addr_78_4, wires_312_5,addr_312_5);

wire[3:0] wires_313_5;

wire[27:0] addr_313_5;

Selector_2 s313_5(wires_78_4[1], addr_78_4, wires_313_5,addr_313_5);

wire[3:0] wires_314_5;

wire[27:0] addr_314_5;

Selector_2 s314_5(wires_78_4[2], addr_78_4, wires_314_5,addr_314_5);

wire[3:0] wires_315_5;

wire[27:0] addr_315_5;

Selector_2 s315_5(wires_78_4[3], addr_78_4, wires_315_5,addr_315_5);

wire[3:0] wires_316_5;

wire[27:0] addr_316_5;

Selector_2 s316_5(wires_79_4[0], addr_79_4, wires_316_5,addr_316_5);

wire[3:0] wires_317_5;

wire[27:0] addr_317_5;

Selector_2 s317_5(wires_79_4[1], addr_79_4, wires_317_5,addr_317_5);

wire[3:0] wires_318_5;

wire[27:0] addr_318_5;

Selector_2 s318_5(wires_79_4[2], addr_79_4, wires_318_5,addr_318_5);

wire[3:0] wires_319_5;

wire[27:0] addr_319_5;

Selector_2 s319_5(wires_79_4[3], addr_79_4, wires_319_5,addr_319_5);

wire[3:0] wires_320_5;

wire[27:0] addr_320_5;

Selector_2 s320_5(wires_80_4[0], addr_80_4, wires_320_5,addr_320_5);

wire[3:0] wires_321_5;

wire[27:0] addr_321_5;

Selector_2 s321_5(wires_80_4[1], addr_80_4, wires_321_5,addr_321_5);

wire[3:0] wires_322_5;

wire[27:0] addr_322_5;

Selector_2 s322_5(wires_80_4[2], addr_80_4, wires_322_5,addr_322_5);

wire[3:0] wires_323_5;

wire[27:0] addr_323_5;

Selector_2 s323_5(wires_80_4[3], addr_80_4, wires_323_5,addr_323_5);

wire[3:0] wires_324_5;

wire[27:0] addr_324_5;

Selector_2 s324_5(wires_81_4[0], addr_81_4, wires_324_5,addr_324_5);

wire[3:0] wires_325_5;

wire[27:0] addr_325_5;

Selector_2 s325_5(wires_81_4[1], addr_81_4, wires_325_5,addr_325_5);

wire[3:0] wires_326_5;

wire[27:0] addr_326_5;

Selector_2 s326_5(wires_81_4[2], addr_81_4, wires_326_5,addr_326_5);

wire[3:0] wires_327_5;

wire[27:0] addr_327_5;

Selector_2 s327_5(wires_81_4[3], addr_81_4, wires_327_5,addr_327_5);

wire[3:0] wires_328_5;

wire[27:0] addr_328_5;

Selector_2 s328_5(wires_82_4[0], addr_82_4, wires_328_5,addr_328_5);

wire[3:0] wires_329_5;

wire[27:0] addr_329_5;

Selector_2 s329_5(wires_82_4[1], addr_82_4, wires_329_5,addr_329_5);

wire[3:0] wires_330_5;

wire[27:0] addr_330_5;

Selector_2 s330_5(wires_82_4[2], addr_82_4, wires_330_5,addr_330_5);

wire[3:0] wires_331_5;

wire[27:0] addr_331_5;

Selector_2 s331_5(wires_82_4[3], addr_82_4, wires_331_5,addr_331_5);

wire[3:0] wires_332_5;

wire[27:0] addr_332_5;

Selector_2 s332_5(wires_83_4[0], addr_83_4, wires_332_5,addr_332_5);

wire[3:0] wires_333_5;

wire[27:0] addr_333_5;

Selector_2 s333_5(wires_83_4[1], addr_83_4, wires_333_5,addr_333_5);

wire[3:0] wires_334_5;

wire[27:0] addr_334_5;

Selector_2 s334_5(wires_83_4[2], addr_83_4, wires_334_5,addr_334_5);

wire[3:0] wires_335_5;

wire[27:0] addr_335_5;

Selector_2 s335_5(wires_83_4[3], addr_83_4, wires_335_5,addr_335_5);

wire[3:0] wires_336_5;

wire[27:0] addr_336_5;

Selector_2 s336_5(wires_84_4[0], addr_84_4, wires_336_5,addr_336_5);

wire[3:0] wires_337_5;

wire[27:0] addr_337_5;

Selector_2 s337_5(wires_84_4[1], addr_84_4, wires_337_5,addr_337_5);

wire[3:0] wires_338_5;

wire[27:0] addr_338_5;

Selector_2 s338_5(wires_84_4[2], addr_84_4, wires_338_5,addr_338_5);

wire[3:0] wires_339_5;

wire[27:0] addr_339_5;

Selector_2 s339_5(wires_84_4[3], addr_84_4, wires_339_5,addr_339_5);

wire[3:0] wires_340_5;

wire[27:0] addr_340_5;

Selector_2 s340_5(wires_85_4[0], addr_85_4, wires_340_5,addr_340_5);

wire[3:0] wires_341_5;

wire[27:0] addr_341_5;

Selector_2 s341_5(wires_85_4[1], addr_85_4, wires_341_5,addr_341_5);

wire[3:0] wires_342_5;

wire[27:0] addr_342_5;

Selector_2 s342_5(wires_85_4[2], addr_85_4, wires_342_5,addr_342_5);

wire[3:0] wires_343_5;

wire[27:0] addr_343_5;

Selector_2 s343_5(wires_85_4[3], addr_85_4, wires_343_5,addr_343_5);

wire[3:0] wires_344_5;

wire[27:0] addr_344_5;

Selector_2 s344_5(wires_86_4[0], addr_86_4, wires_344_5,addr_344_5);

wire[3:0] wires_345_5;

wire[27:0] addr_345_5;

Selector_2 s345_5(wires_86_4[1], addr_86_4, wires_345_5,addr_345_5);

wire[3:0] wires_346_5;

wire[27:0] addr_346_5;

Selector_2 s346_5(wires_86_4[2], addr_86_4, wires_346_5,addr_346_5);

wire[3:0] wires_347_5;

wire[27:0] addr_347_5;

Selector_2 s347_5(wires_86_4[3], addr_86_4, wires_347_5,addr_347_5);

wire[3:0] wires_348_5;

wire[27:0] addr_348_5;

Selector_2 s348_5(wires_87_4[0], addr_87_4, wires_348_5,addr_348_5);

wire[3:0] wires_349_5;

wire[27:0] addr_349_5;

Selector_2 s349_5(wires_87_4[1], addr_87_4, wires_349_5,addr_349_5);

wire[3:0] wires_350_5;

wire[27:0] addr_350_5;

Selector_2 s350_5(wires_87_4[2], addr_87_4, wires_350_5,addr_350_5);

wire[3:0] wires_351_5;

wire[27:0] addr_351_5;

Selector_2 s351_5(wires_87_4[3], addr_87_4, wires_351_5,addr_351_5);

wire[3:0] wires_352_5;

wire[27:0] addr_352_5;

Selector_2 s352_5(wires_88_4[0], addr_88_4, wires_352_5,addr_352_5);

wire[3:0] wires_353_5;

wire[27:0] addr_353_5;

Selector_2 s353_5(wires_88_4[1], addr_88_4, wires_353_5,addr_353_5);

wire[3:0] wires_354_5;

wire[27:0] addr_354_5;

Selector_2 s354_5(wires_88_4[2], addr_88_4, wires_354_5,addr_354_5);

wire[3:0] wires_355_5;

wire[27:0] addr_355_5;

Selector_2 s355_5(wires_88_4[3], addr_88_4, wires_355_5,addr_355_5);

wire[3:0] wires_356_5;

wire[27:0] addr_356_5;

Selector_2 s356_5(wires_89_4[0], addr_89_4, wires_356_5,addr_356_5);

wire[3:0] wires_357_5;

wire[27:0] addr_357_5;

Selector_2 s357_5(wires_89_4[1], addr_89_4, wires_357_5,addr_357_5);

wire[3:0] wires_358_5;

wire[27:0] addr_358_5;

Selector_2 s358_5(wires_89_4[2], addr_89_4, wires_358_5,addr_358_5);

wire[3:0] wires_359_5;

wire[27:0] addr_359_5;

Selector_2 s359_5(wires_89_4[3], addr_89_4, wires_359_5,addr_359_5);

wire[3:0] wires_360_5;

wire[27:0] addr_360_5;

Selector_2 s360_5(wires_90_4[0], addr_90_4, wires_360_5,addr_360_5);

wire[3:0] wires_361_5;

wire[27:0] addr_361_5;

Selector_2 s361_5(wires_90_4[1], addr_90_4, wires_361_5,addr_361_5);

wire[3:0] wires_362_5;

wire[27:0] addr_362_5;

Selector_2 s362_5(wires_90_4[2], addr_90_4, wires_362_5,addr_362_5);

wire[3:0] wires_363_5;

wire[27:0] addr_363_5;

Selector_2 s363_5(wires_90_4[3], addr_90_4, wires_363_5,addr_363_5);

wire[3:0] wires_364_5;

wire[27:0] addr_364_5;

Selector_2 s364_5(wires_91_4[0], addr_91_4, wires_364_5,addr_364_5);

wire[3:0] wires_365_5;

wire[27:0] addr_365_5;

Selector_2 s365_5(wires_91_4[1], addr_91_4, wires_365_5,addr_365_5);

wire[3:0] wires_366_5;

wire[27:0] addr_366_5;

Selector_2 s366_5(wires_91_4[2], addr_91_4, wires_366_5,addr_366_5);

wire[3:0] wires_367_5;

wire[27:0] addr_367_5;

Selector_2 s367_5(wires_91_4[3], addr_91_4, wires_367_5,addr_367_5);

wire[3:0] wires_368_5;

wire[27:0] addr_368_5;

Selector_2 s368_5(wires_92_4[0], addr_92_4, wires_368_5,addr_368_5);

wire[3:0] wires_369_5;

wire[27:0] addr_369_5;

Selector_2 s369_5(wires_92_4[1], addr_92_4, wires_369_5,addr_369_5);

wire[3:0] wires_370_5;

wire[27:0] addr_370_5;

Selector_2 s370_5(wires_92_4[2], addr_92_4, wires_370_5,addr_370_5);

wire[3:0] wires_371_5;

wire[27:0] addr_371_5;

Selector_2 s371_5(wires_92_4[3], addr_92_4, wires_371_5,addr_371_5);

wire[3:0] wires_372_5;

wire[27:0] addr_372_5;

Selector_2 s372_5(wires_93_4[0], addr_93_4, wires_372_5,addr_372_5);

wire[3:0] wires_373_5;

wire[27:0] addr_373_5;

Selector_2 s373_5(wires_93_4[1], addr_93_4, wires_373_5,addr_373_5);

wire[3:0] wires_374_5;

wire[27:0] addr_374_5;

Selector_2 s374_5(wires_93_4[2], addr_93_4, wires_374_5,addr_374_5);

wire[3:0] wires_375_5;

wire[27:0] addr_375_5;

Selector_2 s375_5(wires_93_4[3], addr_93_4, wires_375_5,addr_375_5);

wire[3:0] wires_376_5;

wire[27:0] addr_376_5;

Selector_2 s376_5(wires_94_4[0], addr_94_4, wires_376_5,addr_376_5);

wire[3:0] wires_377_5;

wire[27:0] addr_377_5;

Selector_2 s377_5(wires_94_4[1], addr_94_4, wires_377_5,addr_377_5);

wire[3:0] wires_378_5;

wire[27:0] addr_378_5;

Selector_2 s378_5(wires_94_4[2], addr_94_4, wires_378_5,addr_378_5);

wire[3:0] wires_379_5;

wire[27:0] addr_379_5;

Selector_2 s379_5(wires_94_4[3], addr_94_4, wires_379_5,addr_379_5);

wire[3:0] wires_380_5;

wire[27:0] addr_380_5;

Selector_2 s380_5(wires_95_4[0], addr_95_4, wires_380_5,addr_380_5);

wire[3:0] wires_381_5;

wire[27:0] addr_381_5;

Selector_2 s381_5(wires_95_4[1], addr_95_4, wires_381_5,addr_381_5);

wire[3:0] wires_382_5;

wire[27:0] addr_382_5;

Selector_2 s382_5(wires_95_4[2], addr_95_4, wires_382_5,addr_382_5);

wire[3:0] wires_383_5;

wire[27:0] addr_383_5;

Selector_2 s383_5(wires_95_4[3], addr_95_4, wires_383_5,addr_383_5);

wire[3:0] wires_384_5;

wire[27:0] addr_384_5;

Selector_2 s384_5(wires_96_4[0], addr_96_4, wires_384_5,addr_384_5);

wire[3:0] wires_385_5;

wire[27:0] addr_385_5;

Selector_2 s385_5(wires_96_4[1], addr_96_4, wires_385_5,addr_385_5);

wire[3:0] wires_386_5;

wire[27:0] addr_386_5;

Selector_2 s386_5(wires_96_4[2], addr_96_4, wires_386_5,addr_386_5);

wire[3:0] wires_387_5;

wire[27:0] addr_387_5;

Selector_2 s387_5(wires_96_4[3], addr_96_4, wires_387_5,addr_387_5);

wire[3:0] wires_388_5;

wire[27:0] addr_388_5;

Selector_2 s388_5(wires_97_4[0], addr_97_4, wires_388_5,addr_388_5);

wire[3:0] wires_389_5;

wire[27:0] addr_389_5;

Selector_2 s389_5(wires_97_4[1], addr_97_4, wires_389_5,addr_389_5);

wire[3:0] wires_390_5;

wire[27:0] addr_390_5;

Selector_2 s390_5(wires_97_4[2], addr_97_4, wires_390_5,addr_390_5);

wire[3:0] wires_391_5;

wire[27:0] addr_391_5;

Selector_2 s391_5(wires_97_4[3], addr_97_4, wires_391_5,addr_391_5);

wire[3:0] wires_392_5;

wire[27:0] addr_392_5;

Selector_2 s392_5(wires_98_4[0], addr_98_4, wires_392_5,addr_392_5);

wire[3:0] wires_393_5;

wire[27:0] addr_393_5;

Selector_2 s393_5(wires_98_4[1], addr_98_4, wires_393_5,addr_393_5);

wire[3:0] wires_394_5;

wire[27:0] addr_394_5;

Selector_2 s394_5(wires_98_4[2], addr_98_4, wires_394_5,addr_394_5);

wire[3:0] wires_395_5;

wire[27:0] addr_395_5;

Selector_2 s395_5(wires_98_4[3], addr_98_4, wires_395_5,addr_395_5);

wire[3:0] wires_396_5;

wire[27:0] addr_396_5;

Selector_2 s396_5(wires_99_4[0], addr_99_4, wires_396_5,addr_396_5);

wire[3:0] wires_397_5;

wire[27:0] addr_397_5;

Selector_2 s397_5(wires_99_4[1], addr_99_4, wires_397_5,addr_397_5);

wire[3:0] wires_398_5;

wire[27:0] addr_398_5;

Selector_2 s398_5(wires_99_4[2], addr_99_4, wires_398_5,addr_398_5);

wire[3:0] wires_399_5;

wire[27:0] addr_399_5;

Selector_2 s399_5(wires_99_4[3], addr_99_4, wires_399_5,addr_399_5);

wire[3:0] wires_400_5;

wire[27:0] addr_400_5;

Selector_2 s400_5(wires_100_4[0], addr_100_4, wires_400_5,addr_400_5);

wire[3:0] wires_401_5;

wire[27:0] addr_401_5;

Selector_2 s401_5(wires_100_4[1], addr_100_4, wires_401_5,addr_401_5);

wire[3:0] wires_402_5;

wire[27:0] addr_402_5;

Selector_2 s402_5(wires_100_4[2], addr_100_4, wires_402_5,addr_402_5);

wire[3:0] wires_403_5;

wire[27:0] addr_403_5;

Selector_2 s403_5(wires_100_4[3], addr_100_4, wires_403_5,addr_403_5);

wire[3:0] wires_404_5;

wire[27:0] addr_404_5;

Selector_2 s404_5(wires_101_4[0], addr_101_4, wires_404_5,addr_404_5);

wire[3:0] wires_405_5;

wire[27:0] addr_405_5;

Selector_2 s405_5(wires_101_4[1], addr_101_4, wires_405_5,addr_405_5);

wire[3:0] wires_406_5;

wire[27:0] addr_406_5;

Selector_2 s406_5(wires_101_4[2], addr_101_4, wires_406_5,addr_406_5);

wire[3:0] wires_407_5;

wire[27:0] addr_407_5;

Selector_2 s407_5(wires_101_4[3], addr_101_4, wires_407_5,addr_407_5);

wire[3:0] wires_408_5;

wire[27:0] addr_408_5;

Selector_2 s408_5(wires_102_4[0], addr_102_4, wires_408_5,addr_408_5);

wire[3:0] wires_409_5;

wire[27:0] addr_409_5;

Selector_2 s409_5(wires_102_4[1], addr_102_4, wires_409_5,addr_409_5);

wire[3:0] wires_410_5;

wire[27:0] addr_410_5;

Selector_2 s410_5(wires_102_4[2], addr_102_4, wires_410_5,addr_410_5);

wire[3:0] wires_411_5;

wire[27:0] addr_411_5;

Selector_2 s411_5(wires_102_4[3], addr_102_4, wires_411_5,addr_411_5);

wire[3:0] wires_412_5;

wire[27:0] addr_412_5;

Selector_2 s412_5(wires_103_4[0], addr_103_4, wires_412_5,addr_412_5);

wire[3:0] wires_413_5;

wire[27:0] addr_413_5;

Selector_2 s413_5(wires_103_4[1], addr_103_4, wires_413_5,addr_413_5);

wire[3:0] wires_414_5;

wire[27:0] addr_414_5;

Selector_2 s414_5(wires_103_4[2], addr_103_4, wires_414_5,addr_414_5);

wire[3:0] wires_415_5;

wire[27:0] addr_415_5;

Selector_2 s415_5(wires_103_4[3], addr_103_4, wires_415_5,addr_415_5);

wire[3:0] wires_416_5;

wire[27:0] addr_416_5;

Selector_2 s416_5(wires_104_4[0], addr_104_4, wires_416_5,addr_416_5);

wire[3:0] wires_417_5;

wire[27:0] addr_417_5;

Selector_2 s417_5(wires_104_4[1], addr_104_4, wires_417_5,addr_417_5);

wire[3:0] wires_418_5;

wire[27:0] addr_418_5;

Selector_2 s418_5(wires_104_4[2], addr_104_4, wires_418_5,addr_418_5);

wire[3:0] wires_419_5;

wire[27:0] addr_419_5;

Selector_2 s419_5(wires_104_4[3], addr_104_4, wires_419_5,addr_419_5);

wire[3:0] wires_420_5;

wire[27:0] addr_420_5;

Selector_2 s420_5(wires_105_4[0], addr_105_4, wires_420_5,addr_420_5);

wire[3:0] wires_421_5;

wire[27:0] addr_421_5;

Selector_2 s421_5(wires_105_4[1], addr_105_4, wires_421_5,addr_421_5);

wire[3:0] wires_422_5;

wire[27:0] addr_422_5;

Selector_2 s422_5(wires_105_4[2], addr_105_4, wires_422_5,addr_422_5);

wire[3:0] wires_423_5;

wire[27:0] addr_423_5;

Selector_2 s423_5(wires_105_4[3], addr_105_4, wires_423_5,addr_423_5);

wire[3:0] wires_424_5;

wire[27:0] addr_424_5;

Selector_2 s424_5(wires_106_4[0], addr_106_4, wires_424_5,addr_424_5);

wire[3:0] wires_425_5;

wire[27:0] addr_425_5;

Selector_2 s425_5(wires_106_4[1], addr_106_4, wires_425_5,addr_425_5);

wire[3:0] wires_426_5;

wire[27:0] addr_426_5;

Selector_2 s426_5(wires_106_4[2], addr_106_4, wires_426_5,addr_426_5);

wire[3:0] wires_427_5;

wire[27:0] addr_427_5;

Selector_2 s427_5(wires_106_4[3], addr_106_4, wires_427_5,addr_427_5);

wire[3:0] wires_428_5;

wire[27:0] addr_428_5;

Selector_2 s428_5(wires_107_4[0], addr_107_4, wires_428_5,addr_428_5);

wire[3:0] wires_429_5;

wire[27:0] addr_429_5;

Selector_2 s429_5(wires_107_4[1], addr_107_4, wires_429_5,addr_429_5);

wire[3:0] wires_430_5;

wire[27:0] addr_430_5;

Selector_2 s430_5(wires_107_4[2], addr_107_4, wires_430_5,addr_430_5);

wire[3:0] wires_431_5;

wire[27:0] addr_431_5;

Selector_2 s431_5(wires_107_4[3], addr_107_4, wires_431_5,addr_431_5);

wire[3:0] wires_432_5;

wire[27:0] addr_432_5;

Selector_2 s432_5(wires_108_4[0], addr_108_4, wires_432_5,addr_432_5);

wire[3:0] wires_433_5;

wire[27:0] addr_433_5;

Selector_2 s433_5(wires_108_4[1], addr_108_4, wires_433_5,addr_433_5);

wire[3:0] wires_434_5;

wire[27:0] addr_434_5;

Selector_2 s434_5(wires_108_4[2], addr_108_4, wires_434_5,addr_434_5);

wire[3:0] wires_435_5;

wire[27:0] addr_435_5;

Selector_2 s435_5(wires_108_4[3], addr_108_4, wires_435_5,addr_435_5);

wire[3:0] wires_436_5;

wire[27:0] addr_436_5;

Selector_2 s436_5(wires_109_4[0], addr_109_4, wires_436_5,addr_436_5);

wire[3:0] wires_437_5;

wire[27:0] addr_437_5;

Selector_2 s437_5(wires_109_4[1], addr_109_4, wires_437_5,addr_437_5);

wire[3:0] wires_438_5;

wire[27:0] addr_438_5;

Selector_2 s438_5(wires_109_4[2], addr_109_4, wires_438_5,addr_438_5);

wire[3:0] wires_439_5;

wire[27:0] addr_439_5;

Selector_2 s439_5(wires_109_4[3], addr_109_4, wires_439_5,addr_439_5);

wire[3:0] wires_440_5;

wire[27:0] addr_440_5;

Selector_2 s440_5(wires_110_4[0], addr_110_4, wires_440_5,addr_440_5);

wire[3:0] wires_441_5;

wire[27:0] addr_441_5;

Selector_2 s441_5(wires_110_4[1], addr_110_4, wires_441_5,addr_441_5);

wire[3:0] wires_442_5;

wire[27:0] addr_442_5;

Selector_2 s442_5(wires_110_4[2], addr_110_4, wires_442_5,addr_442_5);

wire[3:0] wires_443_5;

wire[27:0] addr_443_5;

Selector_2 s443_5(wires_110_4[3], addr_110_4, wires_443_5,addr_443_5);

wire[3:0] wires_444_5;

wire[27:0] addr_444_5;

Selector_2 s444_5(wires_111_4[0], addr_111_4, wires_444_5,addr_444_5);

wire[3:0] wires_445_5;

wire[27:0] addr_445_5;

Selector_2 s445_5(wires_111_4[1], addr_111_4, wires_445_5,addr_445_5);

wire[3:0] wires_446_5;

wire[27:0] addr_446_5;

Selector_2 s446_5(wires_111_4[2], addr_111_4, wires_446_5,addr_446_5);

wire[3:0] wires_447_5;

wire[27:0] addr_447_5;

Selector_2 s447_5(wires_111_4[3], addr_111_4, wires_447_5,addr_447_5);

wire[3:0] wires_448_5;

wire[27:0] addr_448_5;

Selector_2 s448_5(wires_112_4[0], addr_112_4, wires_448_5,addr_448_5);

wire[3:0] wires_449_5;

wire[27:0] addr_449_5;

Selector_2 s449_5(wires_112_4[1], addr_112_4, wires_449_5,addr_449_5);

wire[3:0] wires_450_5;

wire[27:0] addr_450_5;

Selector_2 s450_5(wires_112_4[2], addr_112_4, wires_450_5,addr_450_5);

wire[3:0] wires_451_5;

wire[27:0] addr_451_5;

Selector_2 s451_5(wires_112_4[3], addr_112_4, wires_451_5,addr_451_5);

wire[3:0] wires_452_5;

wire[27:0] addr_452_5;

Selector_2 s452_5(wires_113_4[0], addr_113_4, wires_452_5,addr_452_5);

wire[3:0] wires_453_5;

wire[27:0] addr_453_5;

Selector_2 s453_5(wires_113_4[1], addr_113_4, wires_453_5,addr_453_5);

wire[3:0] wires_454_5;

wire[27:0] addr_454_5;

Selector_2 s454_5(wires_113_4[2], addr_113_4, wires_454_5,addr_454_5);

wire[3:0] wires_455_5;

wire[27:0] addr_455_5;

Selector_2 s455_5(wires_113_4[3], addr_113_4, wires_455_5,addr_455_5);

wire[3:0] wires_456_5;

wire[27:0] addr_456_5;

Selector_2 s456_5(wires_114_4[0], addr_114_4, wires_456_5,addr_456_5);

wire[3:0] wires_457_5;

wire[27:0] addr_457_5;

Selector_2 s457_5(wires_114_4[1], addr_114_4, wires_457_5,addr_457_5);

wire[3:0] wires_458_5;

wire[27:0] addr_458_5;

Selector_2 s458_5(wires_114_4[2], addr_114_4, wires_458_5,addr_458_5);

wire[3:0] wires_459_5;

wire[27:0] addr_459_5;

Selector_2 s459_5(wires_114_4[3], addr_114_4, wires_459_5,addr_459_5);

wire[3:0] wires_460_5;

wire[27:0] addr_460_5;

Selector_2 s460_5(wires_115_4[0], addr_115_4, wires_460_5,addr_460_5);

wire[3:0] wires_461_5;

wire[27:0] addr_461_5;

Selector_2 s461_5(wires_115_4[1], addr_115_4, wires_461_5,addr_461_5);

wire[3:0] wires_462_5;

wire[27:0] addr_462_5;

Selector_2 s462_5(wires_115_4[2], addr_115_4, wires_462_5,addr_462_5);

wire[3:0] wires_463_5;

wire[27:0] addr_463_5;

Selector_2 s463_5(wires_115_4[3], addr_115_4, wires_463_5,addr_463_5);

wire[3:0] wires_464_5;

wire[27:0] addr_464_5;

Selector_2 s464_5(wires_116_4[0], addr_116_4, wires_464_5,addr_464_5);

wire[3:0] wires_465_5;

wire[27:0] addr_465_5;

Selector_2 s465_5(wires_116_4[1], addr_116_4, wires_465_5,addr_465_5);

wire[3:0] wires_466_5;

wire[27:0] addr_466_5;

Selector_2 s466_5(wires_116_4[2], addr_116_4, wires_466_5,addr_466_5);

wire[3:0] wires_467_5;

wire[27:0] addr_467_5;

Selector_2 s467_5(wires_116_4[3], addr_116_4, wires_467_5,addr_467_5);

wire[3:0] wires_468_5;

wire[27:0] addr_468_5;

Selector_2 s468_5(wires_117_4[0], addr_117_4, wires_468_5,addr_468_5);

wire[3:0] wires_469_5;

wire[27:0] addr_469_5;

Selector_2 s469_5(wires_117_4[1], addr_117_4, wires_469_5,addr_469_5);

wire[3:0] wires_470_5;

wire[27:0] addr_470_5;

Selector_2 s470_5(wires_117_4[2], addr_117_4, wires_470_5,addr_470_5);

wire[3:0] wires_471_5;

wire[27:0] addr_471_5;

Selector_2 s471_5(wires_117_4[3], addr_117_4, wires_471_5,addr_471_5);

wire[3:0] wires_472_5;

wire[27:0] addr_472_5;

Selector_2 s472_5(wires_118_4[0], addr_118_4, wires_472_5,addr_472_5);

wire[3:0] wires_473_5;

wire[27:0] addr_473_5;

Selector_2 s473_5(wires_118_4[1], addr_118_4, wires_473_5,addr_473_5);

wire[3:0] wires_474_5;

wire[27:0] addr_474_5;

Selector_2 s474_5(wires_118_4[2], addr_118_4, wires_474_5,addr_474_5);

wire[3:0] wires_475_5;

wire[27:0] addr_475_5;

Selector_2 s475_5(wires_118_4[3], addr_118_4, wires_475_5,addr_475_5);

wire[3:0] wires_476_5;

wire[27:0] addr_476_5;

Selector_2 s476_5(wires_119_4[0], addr_119_4, wires_476_5,addr_476_5);

wire[3:0] wires_477_5;

wire[27:0] addr_477_5;

Selector_2 s477_5(wires_119_4[1], addr_119_4, wires_477_5,addr_477_5);

wire[3:0] wires_478_5;

wire[27:0] addr_478_5;

Selector_2 s478_5(wires_119_4[2], addr_119_4, wires_478_5,addr_478_5);

wire[3:0] wires_479_5;

wire[27:0] addr_479_5;

Selector_2 s479_5(wires_119_4[3], addr_119_4, wires_479_5,addr_479_5);

wire[3:0] wires_480_5;

wire[27:0] addr_480_5;

Selector_2 s480_5(wires_120_4[0], addr_120_4, wires_480_5,addr_480_5);

wire[3:0] wires_481_5;

wire[27:0] addr_481_5;

Selector_2 s481_5(wires_120_4[1], addr_120_4, wires_481_5,addr_481_5);

wire[3:0] wires_482_5;

wire[27:0] addr_482_5;

Selector_2 s482_5(wires_120_4[2], addr_120_4, wires_482_5,addr_482_5);

wire[3:0] wires_483_5;

wire[27:0] addr_483_5;

Selector_2 s483_5(wires_120_4[3], addr_120_4, wires_483_5,addr_483_5);

wire[3:0] wires_484_5;

wire[27:0] addr_484_5;

Selector_2 s484_5(wires_121_4[0], addr_121_4, wires_484_5,addr_484_5);

wire[3:0] wires_485_5;

wire[27:0] addr_485_5;

Selector_2 s485_5(wires_121_4[1], addr_121_4, wires_485_5,addr_485_5);

wire[3:0] wires_486_5;

wire[27:0] addr_486_5;

Selector_2 s486_5(wires_121_4[2], addr_121_4, wires_486_5,addr_486_5);

wire[3:0] wires_487_5;

wire[27:0] addr_487_5;

Selector_2 s487_5(wires_121_4[3], addr_121_4, wires_487_5,addr_487_5);

wire[3:0] wires_488_5;

wire[27:0] addr_488_5;

Selector_2 s488_5(wires_122_4[0], addr_122_4, wires_488_5,addr_488_5);

wire[3:0] wires_489_5;

wire[27:0] addr_489_5;

Selector_2 s489_5(wires_122_4[1], addr_122_4, wires_489_5,addr_489_5);

wire[3:0] wires_490_5;

wire[27:0] addr_490_5;

Selector_2 s490_5(wires_122_4[2], addr_122_4, wires_490_5,addr_490_5);

wire[3:0] wires_491_5;

wire[27:0] addr_491_5;

Selector_2 s491_5(wires_122_4[3], addr_122_4, wires_491_5,addr_491_5);

wire[3:0] wires_492_5;

wire[27:0] addr_492_5;

Selector_2 s492_5(wires_123_4[0], addr_123_4, wires_492_5,addr_492_5);

wire[3:0] wires_493_5;

wire[27:0] addr_493_5;

Selector_2 s493_5(wires_123_4[1], addr_123_4, wires_493_5,addr_493_5);

wire[3:0] wires_494_5;

wire[27:0] addr_494_5;

Selector_2 s494_5(wires_123_4[2], addr_123_4, wires_494_5,addr_494_5);

wire[3:0] wires_495_5;

wire[27:0] addr_495_5;

Selector_2 s495_5(wires_123_4[3], addr_123_4, wires_495_5,addr_495_5);

wire[3:0] wires_496_5;

wire[27:0] addr_496_5;

Selector_2 s496_5(wires_124_4[0], addr_124_4, wires_496_5,addr_496_5);

wire[3:0] wires_497_5;

wire[27:0] addr_497_5;

Selector_2 s497_5(wires_124_4[1], addr_124_4, wires_497_5,addr_497_5);

wire[3:0] wires_498_5;

wire[27:0] addr_498_5;

Selector_2 s498_5(wires_124_4[2], addr_124_4, wires_498_5,addr_498_5);

wire[3:0] wires_499_5;

wire[27:0] addr_499_5;

Selector_2 s499_5(wires_124_4[3], addr_124_4, wires_499_5,addr_499_5);

wire[3:0] wires_500_5;

wire[27:0] addr_500_5;

Selector_2 s500_5(wires_125_4[0], addr_125_4, wires_500_5,addr_500_5);

wire[3:0] wires_501_5;

wire[27:0] addr_501_5;

Selector_2 s501_5(wires_125_4[1], addr_125_4, wires_501_5,addr_501_5);

wire[3:0] wires_502_5;

wire[27:0] addr_502_5;

Selector_2 s502_5(wires_125_4[2], addr_125_4, wires_502_5,addr_502_5);

wire[3:0] wires_503_5;

wire[27:0] addr_503_5;

Selector_2 s503_5(wires_125_4[3], addr_125_4, wires_503_5,addr_503_5);

wire[3:0] wires_504_5;

wire[27:0] addr_504_5;

Selector_2 s504_5(wires_126_4[0], addr_126_4, wires_504_5,addr_504_5);

wire[3:0] wires_505_5;

wire[27:0] addr_505_5;

Selector_2 s505_5(wires_126_4[1], addr_126_4, wires_505_5,addr_505_5);

wire[3:0] wires_506_5;

wire[27:0] addr_506_5;

Selector_2 s506_5(wires_126_4[2], addr_126_4, wires_506_5,addr_506_5);

wire[3:0] wires_507_5;

wire[27:0] addr_507_5;

Selector_2 s507_5(wires_126_4[3], addr_126_4, wires_507_5,addr_507_5);

wire[3:0] wires_508_5;

wire[27:0] addr_508_5;

Selector_2 s508_5(wires_127_4[0], addr_127_4, wires_508_5,addr_508_5);

wire[3:0] wires_509_5;

wire[27:0] addr_509_5;

Selector_2 s509_5(wires_127_4[1], addr_127_4, wires_509_5,addr_509_5);

wire[3:0] wires_510_5;

wire[27:0] addr_510_5;

Selector_2 s510_5(wires_127_4[2], addr_127_4, wires_510_5,addr_510_5);

wire[3:0] wires_511_5;

wire[27:0] addr_511_5;

Selector_2 s511_5(wires_127_4[3], addr_127_4, wires_511_5,addr_511_5);

wire[3:0] wires_512_5;

wire[27:0] addr_512_5;

Selector_2 s512_5(wires_128_4[0], addr_128_4, wires_512_5,addr_512_5);

wire[3:0] wires_513_5;

wire[27:0] addr_513_5;

Selector_2 s513_5(wires_128_4[1], addr_128_4, wires_513_5,addr_513_5);

wire[3:0] wires_514_5;

wire[27:0] addr_514_5;

Selector_2 s514_5(wires_128_4[2], addr_128_4, wires_514_5,addr_514_5);

wire[3:0] wires_515_5;

wire[27:0] addr_515_5;

Selector_2 s515_5(wires_128_4[3], addr_128_4, wires_515_5,addr_515_5);

wire[3:0] wires_516_5;

wire[27:0] addr_516_5;

Selector_2 s516_5(wires_129_4[0], addr_129_4, wires_516_5,addr_516_5);

wire[3:0] wires_517_5;

wire[27:0] addr_517_5;

Selector_2 s517_5(wires_129_4[1], addr_129_4, wires_517_5,addr_517_5);

wire[3:0] wires_518_5;

wire[27:0] addr_518_5;

Selector_2 s518_5(wires_129_4[2], addr_129_4, wires_518_5,addr_518_5);

wire[3:0] wires_519_5;

wire[27:0] addr_519_5;

Selector_2 s519_5(wires_129_4[3], addr_129_4, wires_519_5,addr_519_5);

wire[3:0] wires_520_5;

wire[27:0] addr_520_5;

Selector_2 s520_5(wires_130_4[0], addr_130_4, wires_520_5,addr_520_5);

wire[3:0] wires_521_5;

wire[27:0] addr_521_5;

Selector_2 s521_5(wires_130_4[1], addr_130_4, wires_521_5,addr_521_5);

wire[3:0] wires_522_5;

wire[27:0] addr_522_5;

Selector_2 s522_5(wires_130_4[2], addr_130_4, wires_522_5,addr_522_5);

wire[3:0] wires_523_5;

wire[27:0] addr_523_5;

Selector_2 s523_5(wires_130_4[3], addr_130_4, wires_523_5,addr_523_5);

wire[3:0] wires_524_5;

wire[27:0] addr_524_5;

Selector_2 s524_5(wires_131_4[0], addr_131_4, wires_524_5,addr_524_5);

wire[3:0] wires_525_5;

wire[27:0] addr_525_5;

Selector_2 s525_5(wires_131_4[1], addr_131_4, wires_525_5,addr_525_5);

wire[3:0] wires_526_5;

wire[27:0] addr_526_5;

Selector_2 s526_5(wires_131_4[2], addr_131_4, wires_526_5,addr_526_5);

wire[3:0] wires_527_5;

wire[27:0] addr_527_5;

Selector_2 s527_5(wires_131_4[3], addr_131_4, wires_527_5,addr_527_5);

wire[3:0] wires_528_5;

wire[27:0] addr_528_5;

Selector_2 s528_5(wires_132_4[0], addr_132_4, wires_528_5,addr_528_5);

wire[3:0] wires_529_5;

wire[27:0] addr_529_5;

Selector_2 s529_5(wires_132_4[1], addr_132_4, wires_529_5,addr_529_5);

wire[3:0] wires_530_5;

wire[27:0] addr_530_5;

Selector_2 s530_5(wires_132_4[2], addr_132_4, wires_530_5,addr_530_5);

wire[3:0] wires_531_5;

wire[27:0] addr_531_5;

Selector_2 s531_5(wires_132_4[3], addr_132_4, wires_531_5,addr_531_5);

wire[3:0] wires_532_5;

wire[27:0] addr_532_5;

Selector_2 s532_5(wires_133_4[0], addr_133_4, wires_532_5,addr_532_5);

wire[3:0] wires_533_5;

wire[27:0] addr_533_5;

Selector_2 s533_5(wires_133_4[1], addr_133_4, wires_533_5,addr_533_5);

wire[3:0] wires_534_5;

wire[27:0] addr_534_5;

Selector_2 s534_5(wires_133_4[2], addr_133_4, wires_534_5,addr_534_5);

wire[3:0] wires_535_5;

wire[27:0] addr_535_5;

Selector_2 s535_5(wires_133_4[3], addr_133_4, wires_535_5,addr_535_5);

wire[3:0] wires_536_5;

wire[27:0] addr_536_5;

Selector_2 s536_5(wires_134_4[0], addr_134_4, wires_536_5,addr_536_5);

wire[3:0] wires_537_5;

wire[27:0] addr_537_5;

Selector_2 s537_5(wires_134_4[1], addr_134_4, wires_537_5,addr_537_5);

wire[3:0] wires_538_5;

wire[27:0] addr_538_5;

Selector_2 s538_5(wires_134_4[2], addr_134_4, wires_538_5,addr_538_5);

wire[3:0] wires_539_5;

wire[27:0] addr_539_5;

Selector_2 s539_5(wires_134_4[3], addr_134_4, wires_539_5,addr_539_5);

wire[3:0] wires_540_5;

wire[27:0] addr_540_5;

Selector_2 s540_5(wires_135_4[0], addr_135_4, wires_540_5,addr_540_5);

wire[3:0] wires_541_5;

wire[27:0] addr_541_5;

Selector_2 s541_5(wires_135_4[1], addr_135_4, wires_541_5,addr_541_5);

wire[3:0] wires_542_5;

wire[27:0] addr_542_5;

Selector_2 s542_5(wires_135_4[2], addr_135_4, wires_542_5,addr_542_5);

wire[3:0] wires_543_5;

wire[27:0] addr_543_5;

Selector_2 s543_5(wires_135_4[3], addr_135_4, wires_543_5,addr_543_5);

wire[3:0] wires_544_5;

wire[27:0] addr_544_5;

Selector_2 s544_5(wires_136_4[0], addr_136_4, wires_544_5,addr_544_5);

wire[3:0] wires_545_5;

wire[27:0] addr_545_5;

Selector_2 s545_5(wires_136_4[1], addr_136_4, wires_545_5,addr_545_5);

wire[3:0] wires_546_5;

wire[27:0] addr_546_5;

Selector_2 s546_5(wires_136_4[2], addr_136_4, wires_546_5,addr_546_5);

wire[3:0] wires_547_5;

wire[27:0] addr_547_5;

Selector_2 s547_5(wires_136_4[3], addr_136_4, wires_547_5,addr_547_5);

wire[3:0] wires_548_5;

wire[27:0] addr_548_5;

Selector_2 s548_5(wires_137_4[0], addr_137_4, wires_548_5,addr_548_5);

wire[3:0] wires_549_5;

wire[27:0] addr_549_5;

Selector_2 s549_5(wires_137_4[1], addr_137_4, wires_549_5,addr_549_5);

wire[3:0] wires_550_5;

wire[27:0] addr_550_5;

Selector_2 s550_5(wires_137_4[2], addr_137_4, wires_550_5,addr_550_5);

wire[3:0] wires_551_5;

wire[27:0] addr_551_5;

Selector_2 s551_5(wires_137_4[3], addr_137_4, wires_551_5,addr_551_5);

wire[3:0] wires_552_5;

wire[27:0] addr_552_5;

Selector_2 s552_5(wires_138_4[0], addr_138_4, wires_552_5,addr_552_5);

wire[3:0] wires_553_5;

wire[27:0] addr_553_5;

Selector_2 s553_5(wires_138_4[1], addr_138_4, wires_553_5,addr_553_5);

wire[3:0] wires_554_5;

wire[27:0] addr_554_5;

Selector_2 s554_5(wires_138_4[2], addr_138_4, wires_554_5,addr_554_5);

wire[3:0] wires_555_5;

wire[27:0] addr_555_5;

Selector_2 s555_5(wires_138_4[3], addr_138_4, wires_555_5,addr_555_5);

wire[3:0] wires_556_5;

wire[27:0] addr_556_5;

Selector_2 s556_5(wires_139_4[0], addr_139_4, wires_556_5,addr_556_5);

wire[3:0] wires_557_5;

wire[27:0] addr_557_5;

Selector_2 s557_5(wires_139_4[1], addr_139_4, wires_557_5,addr_557_5);

wire[3:0] wires_558_5;

wire[27:0] addr_558_5;

Selector_2 s558_5(wires_139_4[2], addr_139_4, wires_558_5,addr_558_5);

wire[3:0] wires_559_5;

wire[27:0] addr_559_5;

Selector_2 s559_5(wires_139_4[3], addr_139_4, wires_559_5,addr_559_5);

wire[3:0] wires_560_5;

wire[27:0] addr_560_5;

Selector_2 s560_5(wires_140_4[0], addr_140_4, wires_560_5,addr_560_5);

wire[3:0] wires_561_5;

wire[27:0] addr_561_5;

Selector_2 s561_5(wires_140_4[1], addr_140_4, wires_561_5,addr_561_5);

wire[3:0] wires_562_5;

wire[27:0] addr_562_5;

Selector_2 s562_5(wires_140_4[2], addr_140_4, wires_562_5,addr_562_5);

wire[3:0] wires_563_5;

wire[27:0] addr_563_5;

Selector_2 s563_5(wires_140_4[3], addr_140_4, wires_563_5,addr_563_5);

wire[3:0] wires_564_5;

wire[27:0] addr_564_5;

Selector_2 s564_5(wires_141_4[0], addr_141_4, wires_564_5,addr_564_5);

wire[3:0] wires_565_5;

wire[27:0] addr_565_5;

Selector_2 s565_5(wires_141_4[1], addr_141_4, wires_565_5,addr_565_5);

wire[3:0] wires_566_5;

wire[27:0] addr_566_5;

Selector_2 s566_5(wires_141_4[2], addr_141_4, wires_566_5,addr_566_5);

wire[3:0] wires_567_5;

wire[27:0] addr_567_5;

Selector_2 s567_5(wires_141_4[3], addr_141_4, wires_567_5,addr_567_5);

wire[3:0] wires_568_5;

wire[27:0] addr_568_5;

Selector_2 s568_5(wires_142_4[0], addr_142_4, wires_568_5,addr_568_5);

wire[3:0] wires_569_5;

wire[27:0] addr_569_5;

Selector_2 s569_5(wires_142_4[1], addr_142_4, wires_569_5,addr_569_5);

wire[3:0] wires_570_5;

wire[27:0] addr_570_5;

Selector_2 s570_5(wires_142_4[2], addr_142_4, wires_570_5,addr_570_5);

wire[3:0] wires_571_5;

wire[27:0] addr_571_5;

Selector_2 s571_5(wires_142_4[3], addr_142_4, wires_571_5,addr_571_5);

wire[3:0] wires_572_5;

wire[27:0] addr_572_5;

Selector_2 s572_5(wires_143_4[0], addr_143_4, wires_572_5,addr_572_5);

wire[3:0] wires_573_5;

wire[27:0] addr_573_5;

Selector_2 s573_5(wires_143_4[1], addr_143_4, wires_573_5,addr_573_5);

wire[3:0] wires_574_5;

wire[27:0] addr_574_5;

Selector_2 s574_5(wires_143_4[2], addr_143_4, wires_574_5,addr_574_5);

wire[3:0] wires_575_5;

wire[27:0] addr_575_5;

Selector_2 s575_5(wires_143_4[3], addr_143_4, wires_575_5,addr_575_5);

wire[3:0] wires_576_5;

wire[27:0] addr_576_5;

Selector_2 s576_5(wires_144_4[0], addr_144_4, wires_576_5,addr_576_5);

wire[3:0] wires_577_5;

wire[27:0] addr_577_5;

Selector_2 s577_5(wires_144_4[1], addr_144_4, wires_577_5,addr_577_5);

wire[3:0] wires_578_5;

wire[27:0] addr_578_5;

Selector_2 s578_5(wires_144_4[2], addr_144_4, wires_578_5,addr_578_5);

wire[3:0] wires_579_5;

wire[27:0] addr_579_5;

Selector_2 s579_5(wires_144_4[3], addr_144_4, wires_579_5,addr_579_5);

wire[3:0] wires_580_5;

wire[27:0] addr_580_5;

Selector_2 s580_5(wires_145_4[0], addr_145_4, wires_580_5,addr_580_5);

wire[3:0] wires_581_5;

wire[27:0] addr_581_5;

Selector_2 s581_5(wires_145_4[1], addr_145_4, wires_581_5,addr_581_5);

wire[3:0] wires_582_5;

wire[27:0] addr_582_5;

Selector_2 s582_5(wires_145_4[2], addr_145_4, wires_582_5,addr_582_5);

wire[3:0] wires_583_5;

wire[27:0] addr_583_5;

Selector_2 s583_5(wires_145_4[3], addr_145_4, wires_583_5,addr_583_5);

wire[3:0] wires_584_5;

wire[27:0] addr_584_5;

Selector_2 s584_5(wires_146_4[0], addr_146_4, wires_584_5,addr_584_5);

wire[3:0] wires_585_5;

wire[27:0] addr_585_5;

Selector_2 s585_5(wires_146_4[1], addr_146_4, wires_585_5,addr_585_5);

wire[3:0] wires_586_5;

wire[27:0] addr_586_5;

Selector_2 s586_5(wires_146_4[2], addr_146_4, wires_586_5,addr_586_5);

wire[3:0] wires_587_5;

wire[27:0] addr_587_5;

Selector_2 s587_5(wires_146_4[3], addr_146_4, wires_587_5,addr_587_5);

wire[3:0] wires_588_5;

wire[27:0] addr_588_5;

Selector_2 s588_5(wires_147_4[0], addr_147_4, wires_588_5,addr_588_5);

wire[3:0] wires_589_5;

wire[27:0] addr_589_5;

Selector_2 s589_5(wires_147_4[1], addr_147_4, wires_589_5,addr_589_5);

wire[3:0] wires_590_5;

wire[27:0] addr_590_5;

Selector_2 s590_5(wires_147_4[2], addr_147_4, wires_590_5,addr_590_5);

wire[3:0] wires_591_5;

wire[27:0] addr_591_5;

Selector_2 s591_5(wires_147_4[3], addr_147_4, wires_591_5,addr_591_5);

wire[3:0] wires_592_5;

wire[27:0] addr_592_5;

Selector_2 s592_5(wires_148_4[0], addr_148_4, wires_592_5,addr_592_5);

wire[3:0] wires_593_5;

wire[27:0] addr_593_5;

Selector_2 s593_5(wires_148_4[1], addr_148_4, wires_593_5,addr_593_5);

wire[3:0] wires_594_5;

wire[27:0] addr_594_5;

Selector_2 s594_5(wires_148_4[2], addr_148_4, wires_594_5,addr_594_5);

wire[3:0] wires_595_5;

wire[27:0] addr_595_5;

Selector_2 s595_5(wires_148_4[3], addr_148_4, wires_595_5,addr_595_5);

wire[3:0] wires_596_5;

wire[27:0] addr_596_5;

Selector_2 s596_5(wires_149_4[0], addr_149_4, wires_596_5,addr_596_5);

wire[3:0] wires_597_5;

wire[27:0] addr_597_5;

Selector_2 s597_5(wires_149_4[1], addr_149_4, wires_597_5,addr_597_5);

wire[3:0] wires_598_5;

wire[27:0] addr_598_5;

Selector_2 s598_5(wires_149_4[2], addr_149_4, wires_598_5,addr_598_5);

wire[3:0] wires_599_5;

wire[27:0] addr_599_5;

Selector_2 s599_5(wires_149_4[3], addr_149_4, wires_599_5,addr_599_5);

wire[3:0] wires_600_5;

wire[27:0] addr_600_5;

Selector_2 s600_5(wires_150_4[0], addr_150_4, wires_600_5,addr_600_5);

wire[3:0] wires_601_5;

wire[27:0] addr_601_5;

Selector_2 s601_5(wires_150_4[1], addr_150_4, wires_601_5,addr_601_5);

wire[3:0] wires_602_5;

wire[27:0] addr_602_5;

Selector_2 s602_5(wires_150_4[2], addr_150_4, wires_602_5,addr_602_5);

wire[3:0] wires_603_5;

wire[27:0] addr_603_5;

Selector_2 s603_5(wires_150_4[3], addr_150_4, wires_603_5,addr_603_5);

wire[3:0] wires_604_5;

wire[27:0] addr_604_5;

Selector_2 s604_5(wires_151_4[0], addr_151_4, wires_604_5,addr_604_5);

wire[3:0] wires_605_5;

wire[27:0] addr_605_5;

Selector_2 s605_5(wires_151_4[1], addr_151_4, wires_605_5,addr_605_5);

wire[3:0] wires_606_5;

wire[27:0] addr_606_5;

Selector_2 s606_5(wires_151_4[2], addr_151_4, wires_606_5,addr_606_5);

wire[3:0] wires_607_5;

wire[27:0] addr_607_5;

Selector_2 s607_5(wires_151_4[3], addr_151_4, wires_607_5,addr_607_5);

wire[3:0] wires_608_5;

wire[27:0] addr_608_5;

Selector_2 s608_5(wires_152_4[0], addr_152_4, wires_608_5,addr_608_5);

wire[3:0] wires_609_5;

wire[27:0] addr_609_5;

Selector_2 s609_5(wires_152_4[1], addr_152_4, wires_609_5,addr_609_5);

wire[3:0] wires_610_5;

wire[27:0] addr_610_5;

Selector_2 s610_5(wires_152_4[2], addr_152_4, wires_610_5,addr_610_5);

wire[3:0] wires_611_5;

wire[27:0] addr_611_5;

Selector_2 s611_5(wires_152_4[3], addr_152_4, wires_611_5,addr_611_5);

wire[3:0] wires_612_5;

wire[27:0] addr_612_5;

Selector_2 s612_5(wires_153_4[0], addr_153_4, wires_612_5,addr_612_5);

wire[3:0] wires_613_5;

wire[27:0] addr_613_5;

Selector_2 s613_5(wires_153_4[1], addr_153_4, wires_613_5,addr_613_5);

wire[3:0] wires_614_5;

wire[27:0] addr_614_5;

Selector_2 s614_5(wires_153_4[2], addr_153_4, wires_614_5,addr_614_5);

wire[3:0] wires_615_5;

wire[27:0] addr_615_5;

Selector_2 s615_5(wires_153_4[3], addr_153_4, wires_615_5,addr_615_5);

wire[3:0] wires_616_5;

wire[27:0] addr_616_5;

Selector_2 s616_5(wires_154_4[0], addr_154_4, wires_616_5,addr_616_5);

wire[3:0] wires_617_5;

wire[27:0] addr_617_5;

Selector_2 s617_5(wires_154_4[1], addr_154_4, wires_617_5,addr_617_5);

wire[3:0] wires_618_5;

wire[27:0] addr_618_5;

Selector_2 s618_5(wires_154_4[2], addr_154_4, wires_618_5,addr_618_5);

wire[3:0] wires_619_5;

wire[27:0] addr_619_5;

Selector_2 s619_5(wires_154_4[3], addr_154_4, wires_619_5,addr_619_5);

wire[3:0] wires_620_5;

wire[27:0] addr_620_5;

Selector_2 s620_5(wires_155_4[0], addr_155_4, wires_620_5,addr_620_5);

wire[3:0] wires_621_5;

wire[27:0] addr_621_5;

Selector_2 s621_5(wires_155_4[1], addr_155_4, wires_621_5,addr_621_5);

wire[3:0] wires_622_5;

wire[27:0] addr_622_5;

Selector_2 s622_5(wires_155_4[2], addr_155_4, wires_622_5,addr_622_5);

wire[3:0] wires_623_5;

wire[27:0] addr_623_5;

Selector_2 s623_5(wires_155_4[3], addr_155_4, wires_623_5,addr_623_5);

wire[3:0] wires_624_5;

wire[27:0] addr_624_5;

Selector_2 s624_5(wires_156_4[0], addr_156_4, wires_624_5,addr_624_5);

wire[3:0] wires_625_5;

wire[27:0] addr_625_5;

Selector_2 s625_5(wires_156_4[1], addr_156_4, wires_625_5,addr_625_5);

wire[3:0] wires_626_5;

wire[27:0] addr_626_5;

Selector_2 s626_5(wires_156_4[2], addr_156_4, wires_626_5,addr_626_5);

wire[3:0] wires_627_5;

wire[27:0] addr_627_5;

Selector_2 s627_5(wires_156_4[3], addr_156_4, wires_627_5,addr_627_5);

wire[3:0] wires_628_5;

wire[27:0] addr_628_5;

Selector_2 s628_5(wires_157_4[0], addr_157_4, wires_628_5,addr_628_5);

wire[3:0] wires_629_5;

wire[27:0] addr_629_5;

Selector_2 s629_5(wires_157_4[1], addr_157_4, wires_629_5,addr_629_5);

wire[3:0] wires_630_5;

wire[27:0] addr_630_5;

Selector_2 s630_5(wires_157_4[2], addr_157_4, wires_630_5,addr_630_5);

wire[3:0] wires_631_5;

wire[27:0] addr_631_5;

Selector_2 s631_5(wires_157_4[3], addr_157_4, wires_631_5,addr_631_5);

wire[3:0] wires_632_5;

wire[27:0] addr_632_5;

Selector_2 s632_5(wires_158_4[0], addr_158_4, wires_632_5,addr_632_5);

wire[3:0] wires_633_5;

wire[27:0] addr_633_5;

Selector_2 s633_5(wires_158_4[1], addr_158_4, wires_633_5,addr_633_5);

wire[3:0] wires_634_5;

wire[27:0] addr_634_5;

Selector_2 s634_5(wires_158_4[2], addr_158_4, wires_634_5,addr_634_5);

wire[3:0] wires_635_5;

wire[27:0] addr_635_5;

Selector_2 s635_5(wires_158_4[3], addr_158_4, wires_635_5,addr_635_5);

wire[3:0] wires_636_5;

wire[27:0] addr_636_5;

Selector_2 s636_5(wires_159_4[0], addr_159_4, wires_636_5,addr_636_5);

wire[3:0] wires_637_5;

wire[27:0] addr_637_5;

Selector_2 s637_5(wires_159_4[1], addr_159_4, wires_637_5,addr_637_5);

wire[3:0] wires_638_5;

wire[27:0] addr_638_5;

Selector_2 s638_5(wires_159_4[2], addr_159_4, wires_638_5,addr_638_5);

wire[3:0] wires_639_5;

wire[27:0] addr_639_5;

Selector_2 s639_5(wires_159_4[3], addr_159_4, wires_639_5,addr_639_5);

wire[3:0] wires_640_5;

wire[27:0] addr_640_5;

Selector_2 s640_5(wires_160_4[0], addr_160_4, wires_640_5,addr_640_5);

wire[3:0] wires_641_5;

wire[27:0] addr_641_5;

Selector_2 s641_5(wires_160_4[1], addr_160_4, wires_641_5,addr_641_5);

wire[3:0] wires_642_5;

wire[27:0] addr_642_5;

Selector_2 s642_5(wires_160_4[2], addr_160_4, wires_642_5,addr_642_5);

wire[3:0] wires_643_5;

wire[27:0] addr_643_5;

Selector_2 s643_5(wires_160_4[3], addr_160_4, wires_643_5,addr_643_5);

wire[3:0] wires_644_5;

wire[27:0] addr_644_5;

Selector_2 s644_5(wires_161_4[0], addr_161_4, wires_644_5,addr_644_5);

wire[3:0] wires_645_5;

wire[27:0] addr_645_5;

Selector_2 s645_5(wires_161_4[1], addr_161_4, wires_645_5,addr_645_5);

wire[3:0] wires_646_5;

wire[27:0] addr_646_5;

Selector_2 s646_5(wires_161_4[2], addr_161_4, wires_646_5,addr_646_5);

wire[3:0] wires_647_5;

wire[27:0] addr_647_5;

Selector_2 s647_5(wires_161_4[3], addr_161_4, wires_647_5,addr_647_5);

wire[3:0] wires_648_5;

wire[27:0] addr_648_5;

Selector_2 s648_5(wires_162_4[0], addr_162_4, wires_648_5,addr_648_5);

wire[3:0] wires_649_5;

wire[27:0] addr_649_5;

Selector_2 s649_5(wires_162_4[1], addr_162_4, wires_649_5,addr_649_5);

wire[3:0] wires_650_5;

wire[27:0] addr_650_5;

Selector_2 s650_5(wires_162_4[2], addr_162_4, wires_650_5,addr_650_5);

wire[3:0] wires_651_5;

wire[27:0] addr_651_5;

Selector_2 s651_5(wires_162_4[3], addr_162_4, wires_651_5,addr_651_5);

wire[3:0] wires_652_5;

wire[27:0] addr_652_5;

Selector_2 s652_5(wires_163_4[0], addr_163_4, wires_652_5,addr_652_5);

wire[3:0] wires_653_5;

wire[27:0] addr_653_5;

Selector_2 s653_5(wires_163_4[1], addr_163_4, wires_653_5,addr_653_5);

wire[3:0] wires_654_5;

wire[27:0] addr_654_5;

Selector_2 s654_5(wires_163_4[2], addr_163_4, wires_654_5,addr_654_5);

wire[3:0] wires_655_5;

wire[27:0] addr_655_5;

Selector_2 s655_5(wires_163_4[3], addr_163_4, wires_655_5,addr_655_5);

wire[3:0] wires_656_5;

wire[27:0] addr_656_5;

Selector_2 s656_5(wires_164_4[0], addr_164_4, wires_656_5,addr_656_5);

wire[3:0] wires_657_5;

wire[27:0] addr_657_5;

Selector_2 s657_5(wires_164_4[1], addr_164_4, wires_657_5,addr_657_5);

wire[3:0] wires_658_5;

wire[27:0] addr_658_5;

Selector_2 s658_5(wires_164_4[2], addr_164_4, wires_658_5,addr_658_5);

wire[3:0] wires_659_5;

wire[27:0] addr_659_5;

Selector_2 s659_5(wires_164_4[3], addr_164_4, wires_659_5,addr_659_5);

wire[3:0] wires_660_5;

wire[27:0] addr_660_5;

Selector_2 s660_5(wires_165_4[0], addr_165_4, wires_660_5,addr_660_5);

wire[3:0] wires_661_5;

wire[27:0] addr_661_5;

Selector_2 s661_5(wires_165_4[1], addr_165_4, wires_661_5,addr_661_5);

wire[3:0] wires_662_5;

wire[27:0] addr_662_5;

Selector_2 s662_5(wires_165_4[2], addr_165_4, wires_662_5,addr_662_5);

wire[3:0] wires_663_5;

wire[27:0] addr_663_5;

Selector_2 s663_5(wires_165_4[3], addr_165_4, wires_663_5,addr_663_5);

wire[3:0] wires_664_5;

wire[27:0] addr_664_5;

Selector_2 s664_5(wires_166_4[0], addr_166_4, wires_664_5,addr_664_5);

wire[3:0] wires_665_5;

wire[27:0] addr_665_5;

Selector_2 s665_5(wires_166_4[1], addr_166_4, wires_665_5,addr_665_5);

wire[3:0] wires_666_5;

wire[27:0] addr_666_5;

Selector_2 s666_5(wires_166_4[2], addr_166_4, wires_666_5,addr_666_5);

wire[3:0] wires_667_5;

wire[27:0] addr_667_5;

Selector_2 s667_5(wires_166_4[3], addr_166_4, wires_667_5,addr_667_5);

wire[3:0] wires_668_5;

wire[27:0] addr_668_5;

Selector_2 s668_5(wires_167_4[0], addr_167_4, wires_668_5,addr_668_5);

wire[3:0] wires_669_5;

wire[27:0] addr_669_5;

Selector_2 s669_5(wires_167_4[1], addr_167_4, wires_669_5,addr_669_5);

wire[3:0] wires_670_5;

wire[27:0] addr_670_5;

Selector_2 s670_5(wires_167_4[2], addr_167_4, wires_670_5,addr_670_5);

wire[3:0] wires_671_5;

wire[27:0] addr_671_5;

Selector_2 s671_5(wires_167_4[3], addr_167_4, wires_671_5,addr_671_5);

wire[3:0] wires_672_5;

wire[27:0] addr_672_5;

Selector_2 s672_5(wires_168_4[0], addr_168_4, wires_672_5,addr_672_5);

wire[3:0] wires_673_5;

wire[27:0] addr_673_5;

Selector_2 s673_5(wires_168_4[1], addr_168_4, wires_673_5,addr_673_5);

wire[3:0] wires_674_5;

wire[27:0] addr_674_5;

Selector_2 s674_5(wires_168_4[2], addr_168_4, wires_674_5,addr_674_5);

wire[3:0] wires_675_5;

wire[27:0] addr_675_5;

Selector_2 s675_5(wires_168_4[3], addr_168_4, wires_675_5,addr_675_5);

wire[3:0] wires_676_5;

wire[27:0] addr_676_5;

Selector_2 s676_5(wires_169_4[0], addr_169_4, wires_676_5,addr_676_5);

wire[3:0] wires_677_5;

wire[27:0] addr_677_5;

Selector_2 s677_5(wires_169_4[1], addr_169_4, wires_677_5,addr_677_5);

wire[3:0] wires_678_5;

wire[27:0] addr_678_5;

Selector_2 s678_5(wires_169_4[2], addr_169_4, wires_678_5,addr_678_5);

wire[3:0] wires_679_5;

wire[27:0] addr_679_5;

Selector_2 s679_5(wires_169_4[3], addr_169_4, wires_679_5,addr_679_5);

wire[3:0] wires_680_5;

wire[27:0] addr_680_5;

Selector_2 s680_5(wires_170_4[0], addr_170_4, wires_680_5,addr_680_5);

wire[3:0] wires_681_5;

wire[27:0] addr_681_5;

Selector_2 s681_5(wires_170_4[1], addr_170_4, wires_681_5,addr_681_5);

wire[3:0] wires_682_5;

wire[27:0] addr_682_5;

Selector_2 s682_5(wires_170_4[2], addr_170_4, wires_682_5,addr_682_5);

wire[3:0] wires_683_5;

wire[27:0] addr_683_5;

Selector_2 s683_5(wires_170_4[3], addr_170_4, wires_683_5,addr_683_5);

wire[3:0] wires_684_5;

wire[27:0] addr_684_5;

Selector_2 s684_5(wires_171_4[0], addr_171_4, wires_684_5,addr_684_5);

wire[3:0] wires_685_5;

wire[27:0] addr_685_5;

Selector_2 s685_5(wires_171_4[1], addr_171_4, wires_685_5,addr_685_5);

wire[3:0] wires_686_5;

wire[27:0] addr_686_5;

Selector_2 s686_5(wires_171_4[2], addr_171_4, wires_686_5,addr_686_5);

wire[3:0] wires_687_5;

wire[27:0] addr_687_5;

Selector_2 s687_5(wires_171_4[3], addr_171_4, wires_687_5,addr_687_5);

wire[3:0] wires_688_5;

wire[27:0] addr_688_5;

Selector_2 s688_5(wires_172_4[0], addr_172_4, wires_688_5,addr_688_5);

wire[3:0] wires_689_5;

wire[27:0] addr_689_5;

Selector_2 s689_5(wires_172_4[1], addr_172_4, wires_689_5,addr_689_5);

wire[3:0] wires_690_5;

wire[27:0] addr_690_5;

Selector_2 s690_5(wires_172_4[2], addr_172_4, wires_690_5,addr_690_5);

wire[3:0] wires_691_5;

wire[27:0] addr_691_5;

Selector_2 s691_5(wires_172_4[3], addr_172_4, wires_691_5,addr_691_5);

wire[3:0] wires_692_5;

wire[27:0] addr_692_5;

Selector_2 s692_5(wires_173_4[0], addr_173_4, wires_692_5,addr_692_5);

wire[3:0] wires_693_5;

wire[27:0] addr_693_5;

Selector_2 s693_5(wires_173_4[1], addr_173_4, wires_693_5,addr_693_5);

wire[3:0] wires_694_5;

wire[27:0] addr_694_5;

Selector_2 s694_5(wires_173_4[2], addr_173_4, wires_694_5,addr_694_5);

wire[3:0] wires_695_5;

wire[27:0] addr_695_5;

Selector_2 s695_5(wires_173_4[3], addr_173_4, wires_695_5,addr_695_5);

wire[3:0] wires_696_5;

wire[27:0] addr_696_5;

Selector_2 s696_5(wires_174_4[0], addr_174_4, wires_696_5,addr_696_5);

wire[3:0] wires_697_5;

wire[27:0] addr_697_5;

Selector_2 s697_5(wires_174_4[1], addr_174_4, wires_697_5,addr_697_5);

wire[3:0] wires_698_5;

wire[27:0] addr_698_5;

Selector_2 s698_5(wires_174_4[2], addr_174_4, wires_698_5,addr_698_5);

wire[3:0] wires_699_5;

wire[27:0] addr_699_5;

Selector_2 s699_5(wires_174_4[3], addr_174_4, wires_699_5,addr_699_5);

wire[3:0] wires_700_5;

wire[27:0] addr_700_5;

Selector_2 s700_5(wires_175_4[0], addr_175_4, wires_700_5,addr_700_5);

wire[3:0] wires_701_5;

wire[27:0] addr_701_5;

Selector_2 s701_5(wires_175_4[1], addr_175_4, wires_701_5,addr_701_5);

wire[3:0] wires_702_5;

wire[27:0] addr_702_5;

Selector_2 s702_5(wires_175_4[2], addr_175_4, wires_702_5,addr_702_5);

wire[3:0] wires_703_5;

wire[27:0] addr_703_5;

Selector_2 s703_5(wires_175_4[3], addr_175_4, wires_703_5,addr_703_5);

wire[3:0] wires_704_5;

wire[27:0] addr_704_5;

Selector_2 s704_5(wires_176_4[0], addr_176_4, wires_704_5,addr_704_5);

wire[3:0] wires_705_5;

wire[27:0] addr_705_5;

Selector_2 s705_5(wires_176_4[1], addr_176_4, wires_705_5,addr_705_5);

wire[3:0] wires_706_5;

wire[27:0] addr_706_5;

Selector_2 s706_5(wires_176_4[2], addr_176_4, wires_706_5,addr_706_5);

wire[3:0] wires_707_5;

wire[27:0] addr_707_5;

Selector_2 s707_5(wires_176_4[3], addr_176_4, wires_707_5,addr_707_5);

wire[3:0] wires_708_5;

wire[27:0] addr_708_5;

Selector_2 s708_5(wires_177_4[0], addr_177_4, wires_708_5,addr_708_5);

wire[3:0] wires_709_5;

wire[27:0] addr_709_5;

Selector_2 s709_5(wires_177_4[1], addr_177_4, wires_709_5,addr_709_5);

wire[3:0] wires_710_5;

wire[27:0] addr_710_5;

Selector_2 s710_5(wires_177_4[2], addr_177_4, wires_710_5,addr_710_5);

wire[3:0] wires_711_5;

wire[27:0] addr_711_5;

Selector_2 s711_5(wires_177_4[3], addr_177_4, wires_711_5,addr_711_5);

wire[3:0] wires_712_5;

wire[27:0] addr_712_5;

Selector_2 s712_5(wires_178_4[0], addr_178_4, wires_712_5,addr_712_5);

wire[3:0] wires_713_5;

wire[27:0] addr_713_5;

Selector_2 s713_5(wires_178_4[1], addr_178_4, wires_713_5,addr_713_5);

wire[3:0] wires_714_5;

wire[27:0] addr_714_5;

Selector_2 s714_5(wires_178_4[2], addr_178_4, wires_714_5,addr_714_5);

wire[3:0] wires_715_5;

wire[27:0] addr_715_5;

Selector_2 s715_5(wires_178_4[3], addr_178_4, wires_715_5,addr_715_5);

wire[3:0] wires_716_5;

wire[27:0] addr_716_5;

Selector_2 s716_5(wires_179_4[0], addr_179_4, wires_716_5,addr_716_5);

wire[3:0] wires_717_5;

wire[27:0] addr_717_5;

Selector_2 s717_5(wires_179_4[1], addr_179_4, wires_717_5,addr_717_5);

wire[3:0] wires_718_5;

wire[27:0] addr_718_5;

Selector_2 s718_5(wires_179_4[2], addr_179_4, wires_718_5,addr_718_5);

wire[3:0] wires_719_5;

wire[27:0] addr_719_5;

Selector_2 s719_5(wires_179_4[3], addr_179_4, wires_719_5,addr_719_5);

wire[3:0] wires_720_5;

wire[27:0] addr_720_5;

Selector_2 s720_5(wires_180_4[0], addr_180_4, wires_720_5,addr_720_5);

wire[3:0] wires_721_5;

wire[27:0] addr_721_5;

Selector_2 s721_5(wires_180_4[1], addr_180_4, wires_721_5,addr_721_5);

wire[3:0] wires_722_5;

wire[27:0] addr_722_5;

Selector_2 s722_5(wires_180_4[2], addr_180_4, wires_722_5,addr_722_5);

wire[3:0] wires_723_5;

wire[27:0] addr_723_5;

Selector_2 s723_5(wires_180_4[3], addr_180_4, wires_723_5,addr_723_5);

wire[3:0] wires_724_5;

wire[27:0] addr_724_5;

Selector_2 s724_5(wires_181_4[0], addr_181_4, wires_724_5,addr_724_5);

wire[3:0] wires_725_5;

wire[27:0] addr_725_5;

Selector_2 s725_5(wires_181_4[1], addr_181_4, wires_725_5,addr_725_5);

wire[3:0] wires_726_5;

wire[27:0] addr_726_5;

Selector_2 s726_5(wires_181_4[2], addr_181_4, wires_726_5,addr_726_5);

wire[3:0] wires_727_5;

wire[27:0] addr_727_5;

Selector_2 s727_5(wires_181_4[3], addr_181_4, wires_727_5,addr_727_5);

wire[3:0] wires_728_5;

wire[27:0] addr_728_5;

Selector_2 s728_5(wires_182_4[0], addr_182_4, wires_728_5,addr_728_5);

wire[3:0] wires_729_5;

wire[27:0] addr_729_5;

Selector_2 s729_5(wires_182_4[1], addr_182_4, wires_729_5,addr_729_5);

wire[3:0] wires_730_5;

wire[27:0] addr_730_5;

Selector_2 s730_5(wires_182_4[2], addr_182_4, wires_730_5,addr_730_5);

wire[3:0] wires_731_5;

wire[27:0] addr_731_5;

Selector_2 s731_5(wires_182_4[3], addr_182_4, wires_731_5,addr_731_5);

wire[3:0] wires_732_5;

wire[27:0] addr_732_5;

Selector_2 s732_5(wires_183_4[0], addr_183_4, wires_732_5,addr_732_5);

wire[3:0] wires_733_5;

wire[27:0] addr_733_5;

Selector_2 s733_5(wires_183_4[1], addr_183_4, wires_733_5,addr_733_5);

wire[3:0] wires_734_5;

wire[27:0] addr_734_5;

Selector_2 s734_5(wires_183_4[2], addr_183_4, wires_734_5,addr_734_5);

wire[3:0] wires_735_5;

wire[27:0] addr_735_5;

Selector_2 s735_5(wires_183_4[3], addr_183_4, wires_735_5,addr_735_5);

wire[3:0] wires_736_5;

wire[27:0] addr_736_5;

Selector_2 s736_5(wires_184_4[0], addr_184_4, wires_736_5,addr_736_5);

wire[3:0] wires_737_5;

wire[27:0] addr_737_5;

Selector_2 s737_5(wires_184_4[1], addr_184_4, wires_737_5,addr_737_5);

wire[3:0] wires_738_5;

wire[27:0] addr_738_5;

Selector_2 s738_5(wires_184_4[2], addr_184_4, wires_738_5,addr_738_5);

wire[3:0] wires_739_5;

wire[27:0] addr_739_5;

Selector_2 s739_5(wires_184_4[3], addr_184_4, wires_739_5,addr_739_5);

wire[3:0] wires_740_5;

wire[27:0] addr_740_5;

Selector_2 s740_5(wires_185_4[0], addr_185_4, wires_740_5,addr_740_5);

wire[3:0] wires_741_5;

wire[27:0] addr_741_5;

Selector_2 s741_5(wires_185_4[1], addr_185_4, wires_741_5,addr_741_5);

wire[3:0] wires_742_5;

wire[27:0] addr_742_5;

Selector_2 s742_5(wires_185_4[2], addr_185_4, wires_742_5,addr_742_5);

wire[3:0] wires_743_5;

wire[27:0] addr_743_5;

Selector_2 s743_5(wires_185_4[3], addr_185_4, wires_743_5,addr_743_5);

wire[3:0] wires_744_5;

wire[27:0] addr_744_5;

Selector_2 s744_5(wires_186_4[0], addr_186_4, wires_744_5,addr_744_5);

wire[3:0] wires_745_5;

wire[27:0] addr_745_5;

Selector_2 s745_5(wires_186_4[1], addr_186_4, wires_745_5,addr_745_5);

wire[3:0] wires_746_5;

wire[27:0] addr_746_5;

Selector_2 s746_5(wires_186_4[2], addr_186_4, wires_746_5,addr_746_5);

wire[3:0] wires_747_5;

wire[27:0] addr_747_5;

Selector_2 s747_5(wires_186_4[3], addr_186_4, wires_747_5,addr_747_5);

wire[3:0] wires_748_5;

wire[27:0] addr_748_5;

Selector_2 s748_5(wires_187_4[0], addr_187_4, wires_748_5,addr_748_5);

wire[3:0] wires_749_5;

wire[27:0] addr_749_5;

Selector_2 s749_5(wires_187_4[1], addr_187_4, wires_749_5,addr_749_5);

wire[3:0] wires_750_5;

wire[27:0] addr_750_5;

Selector_2 s750_5(wires_187_4[2], addr_187_4, wires_750_5,addr_750_5);

wire[3:0] wires_751_5;

wire[27:0] addr_751_5;

Selector_2 s751_5(wires_187_4[3], addr_187_4, wires_751_5,addr_751_5);

wire[3:0] wires_752_5;

wire[27:0] addr_752_5;

Selector_2 s752_5(wires_188_4[0], addr_188_4, wires_752_5,addr_752_5);

wire[3:0] wires_753_5;

wire[27:0] addr_753_5;

Selector_2 s753_5(wires_188_4[1], addr_188_4, wires_753_5,addr_753_5);

wire[3:0] wires_754_5;

wire[27:0] addr_754_5;

Selector_2 s754_5(wires_188_4[2], addr_188_4, wires_754_5,addr_754_5);

wire[3:0] wires_755_5;

wire[27:0] addr_755_5;

Selector_2 s755_5(wires_188_4[3], addr_188_4, wires_755_5,addr_755_5);

wire[3:0] wires_756_5;

wire[27:0] addr_756_5;

Selector_2 s756_5(wires_189_4[0], addr_189_4, wires_756_5,addr_756_5);

wire[3:0] wires_757_5;

wire[27:0] addr_757_5;

Selector_2 s757_5(wires_189_4[1], addr_189_4, wires_757_5,addr_757_5);

wire[3:0] wires_758_5;

wire[27:0] addr_758_5;

Selector_2 s758_5(wires_189_4[2], addr_189_4, wires_758_5,addr_758_5);

wire[3:0] wires_759_5;

wire[27:0] addr_759_5;

Selector_2 s759_5(wires_189_4[3], addr_189_4, wires_759_5,addr_759_5);

wire[3:0] wires_760_5;

wire[27:0] addr_760_5;

Selector_2 s760_5(wires_190_4[0], addr_190_4, wires_760_5,addr_760_5);

wire[3:0] wires_761_5;

wire[27:0] addr_761_5;

Selector_2 s761_5(wires_190_4[1], addr_190_4, wires_761_5,addr_761_5);

wire[3:0] wires_762_5;

wire[27:0] addr_762_5;

Selector_2 s762_5(wires_190_4[2], addr_190_4, wires_762_5,addr_762_5);

wire[3:0] wires_763_5;

wire[27:0] addr_763_5;

Selector_2 s763_5(wires_190_4[3], addr_190_4, wires_763_5,addr_763_5);

wire[3:0] wires_764_5;

wire[27:0] addr_764_5;

Selector_2 s764_5(wires_191_4[0], addr_191_4, wires_764_5,addr_764_5);

wire[3:0] wires_765_5;

wire[27:0] addr_765_5;

Selector_2 s765_5(wires_191_4[1], addr_191_4, wires_765_5,addr_765_5);

wire[3:0] wires_766_5;

wire[27:0] addr_766_5;

Selector_2 s766_5(wires_191_4[2], addr_191_4, wires_766_5,addr_766_5);

wire[3:0] wires_767_5;

wire[27:0] addr_767_5;

Selector_2 s767_5(wires_191_4[3], addr_191_4, wires_767_5,addr_767_5);

wire[3:0] wires_768_5;

wire[27:0] addr_768_5;

Selector_2 s768_5(wires_192_4[0], addr_192_4, wires_768_5,addr_768_5);

wire[3:0] wires_769_5;

wire[27:0] addr_769_5;

Selector_2 s769_5(wires_192_4[1], addr_192_4, wires_769_5,addr_769_5);

wire[3:0] wires_770_5;

wire[27:0] addr_770_5;

Selector_2 s770_5(wires_192_4[2], addr_192_4, wires_770_5,addr_770_5);

wire[3:0] wires_771_5;

wire[27:0] addr_771_5;

Selector_2 s771_5(wires_192_4[3], addr_192_4, wires_771_5,addr_771_5);

wire[3:0] wires_772_5;

wire[27:0] addr_772_5;

Selector_2 s772_5(wires_193_4[0], addr_193_4, wires_772_5,addr_772_5);

wire[3:0] wires_773_5;

wire[27:0] addr_773_5;

Selector_2 s773_5(wires_193_4[1], addr_193_4, wires_773_5,addr_773_5);

wire[3:0] wires_774_5;

wire[27:0] addr_774_5;

Selector_2 s774_5(wires_193_4[2], addr_193_4, wires_774_5,addr_774_5);

wire[3:0] wires_775_5;

wire[27:0] addr_775_5;

Selector_2 s775_5(wires_193_4[3], addr_193_4, wires_775_5,addr_775_5);

wire[3:0] wires_776_5;

wire[27:0] addr_776_5;

Selector_2 s776_5(wires_194_4[0], addr_194_4, wires_776_5,addr_776_5);

wire[3:0] wires_777_5;

wire[27:0] addr_777_5;

Selector_2 s777_5(wires_194_4[1], addr_194_4, wires_777_5,addr_777_5);

wire[3:0] wires_778_5;

wire[27:0] addr_778_5;

Selector_2 s778_5(wires_194_4[2], addr_194_4, wires_778_5,addr_778_5);

wire[3:0] wires_779_5;

wire[27:0] addr_779_5;

Selector_2 s779_5(wires_194_4[3], addr_194_4, wires_779_5,addr_779_5);

wire[3:0] wires_780_5;

wire[27:0] addr_780_5;

Selector_2 s780_5(wires_195_4[0], addr_195_4, wires_780_5,addr_780_5);

wire[3:0] wires_781_5;

wire[27:0] addr_781_5;

Selector_2 s781_5(wires_195_4[1], addr_195_4, wires_781_5,addr_781_5);

wire[3:0] wires_782_5;

wire[27:0] addr_782_5;

Selector_2 s782_5(wires_195_4[2], addr_195_4, wires_782_5,addr_782_5);

wire[3:0] wires_783_5;

wire[27:0] addr_783_5;

Selector_2 s783_5(wires_195_4[3], addr_195_4, wires_783_5,addr_783_5);

wire[3:0] wires_784_5;

wire[27:0] addr_784_5;

Selector_2 s784_5(wires_196_4[0], addr_196_4, wires_784_5,addr_784_5);

wire[3:0] wires_785_5;

wire[27:0] addr_785_5;

Selector_2 s785_5(wires_196_4[1], addr_196_4, wires_785_5,addr_785_5);

wire[3:0] wires_786_5;

wire[27:0] addr_786_5;

Selector_2 s786_5(wires_196_4[2], addr_196_4, wires_786_5,addr_786_5);

wire[3:0] wires_787_5;

wire[27:0] addr_787_5;

Selector_2 s787_5(wires_196_4[3], addr_196_4, wires_787_5,addr_787_5);

wire[3:0] wires_788_5;

wire[27:0] addr_788_5;

Selector_2 s788_5(wires_197_4[0], addr_197_4, wires_788_5,addr_788_5);

wire[3:0] wires_789_5;

wire[27:0] addr_789_5;

Selector_2 s789_5(wires_197_4[1], addr_197_4, wires_789_5,addr_789_5);

wire[3:0] wires_790_5;

wire[27:0] addr_790_5;

Selector_2 s790_5(wires_197_4[2], addr_197_4, wires_790_5,addr_790_5);

wire[3:0] wires_791_5;

wire[27:0] addr_791_5;

Selector_2 s791_5(wires_197_4[3], addr_197_4, wires_791_5,addr_791_5);

wire[3:0] wires_792_5;

wire[27:0] addr_792_5;

Selector_2 s792_5(wires_198_4[0], addr_198_4, wires_792_5,addr_792_5);

wire[3:0] wires_793_5;

wire[27:0] addr_793_5;

Selector_2 s793_5(wires_198_4[1], addr_198_4, wires_793_5,addr_793_5);

wire[3:0] wires_794_5;

wire[27:0] addr_794_5;

Selector_2 s794_5(wires_198_4[2], addr_198_4, wires_794_5,addr_794_5);

wire[3:0] wires_795_5;

wire[27:0] addr_795_5;

Selector_2 s795_5(wires_198_4[3], addr_198_4, wires_795_5,addr_795_5);

wire[3:0] wires_796_5;

wire[27:0] addr_796_5;

Selector_2 s796_5(wires_199_4[0], addr_199_4, wires_796_5,addr_796_5);

wire[3:0] wires_797_5;

wire[27:0] addr_797_5;

Selector_2 s797_5(wires_199_4[1], addr_199_4, wires_797_5,addr_797_5);

wire[3:0] wires_798_5;

wire[27:0] addr_798_5;

Selector_2 s798_5(wires_199_4[2], addr_199_4, wires_798_5,addr_798_5);

wire[3:0] wires_799_5;

wire[27:0] addr_799_5;

Selector_2 s799_5(wires_199_4[3], addr_199_4, wires_799_5,addr_799_5);

wire[3:0] wires_800_5;

wire[27:0] addr_800_5;

Selector_2 s800_5(wires_200_4[0], addr_200_4, wires_800_5,addr_800_5);

wire[3:0] wires_801_5;

wire[27:0] addr_801_5;

Selector_2 s801_5(wires_200_4[1], addr_200_4, wires_801_5,addr_801_5);

wire[3:0] wires_802_5;

wire[27:0] addr_802_5;

Selector_2 s802_5(wires_200_4[2], addr_200_4, wires_802_5,addr_802_5);

wire[3:0] wires_803_5;

wire[27:0] addr_803_5;

Selector_2 s803_5(wires_200_4[3], addr_200_4, wires_803_5,addr_803_5);

wire[3:0] wires_804_5;

wire[27:0] addr_804_5;

Selector_2 s804_5(wires_201_4[0], addr_201_4, wires_804_5,addr_804_5);

wire[3:0] wires_805_5;

wire[27:0] addr_805_5;

Selector_2 s805_5(wires_201_4[1], addr_201_4, wires_805_5,addr_805_5);

wire[3:0] wires_806_5;

wire[27:0] addr_806_5;

Selector_2 s806_5(wires_201_4[2], addr_201_4, wires_806_5,addr_806_5);

wire[3:0] wires_807_5;

wire[27:0] addr_807_5;

Selector_2 s807_5(wires_201_4[3], addr_201_4, wires_807_5,addr_807_5);

wire[3:0] wires_808_5;

wire[27:0] addr_808_5;

Selector_2 s808_5(wires_202_4[0], addr_202_4, wires_808_5,addr_808_5);

wire[3:0] wires_809_5;

wire[27:0] addr_809_5;

Selector_2 s809_5(wires_202_4[1], addr_202_4, wires_809_5,addr_809_5);

wire[3:0] wires_810_5;

wire[27:0] addr_810_5;

Selector_2 s810_5(wires_202_4[2], addr_202_4, wires_810_5,addr_810_5);

wire[3:0] wires_811_5;

wire[27:0] addr_811_5;

Selector_2 s811_5(wires_202_4[3], addr_202_4, wires_811_5,addr_811_5);

wire[3:0] wires_812_5;

wire[27:0] addr_812_5;

Selector_2 s812_5(wires_203_4[0], addr_203_4, wires_812_5,addr_812_5);

wire[3:0] wires_813_5;

wire[27:0] addr_813_5;

Selector_2 s813_5(wires_203_4[1], addr_203_4, wires_813_5,addr_813_5);

wire[3:0] wires_814_5;

wire[27:0] addr_814_5;

Selector_2 s814_5(wires_203_4[2], addr_203_4, wires_814_5,addr_814_5);

wire[3:0] wires_815_5;

wire[27:0] addr_815_5;

Selector_2 s815_5(wires_203_4[3], addr_203_4, wires_815_5,addr_815_5);

wire[3:0] wires_816_5;

wire[27:0] addr_816_5;

Selector_2 s816_5(wires_204_4[0], addr_204_4, wires_816_5,addr_816_5);

wire[3:0] wires_817_5;

wire[27:0] addr_817_5;

Selector_2 s817_5(wires_204_4[1], addr_204_4, wires_817_5,addr_817_5);

wire[3:0] wires_818_5;

wire[27:0] addr_818_5;

Selector_2 s818_5(wires_204_4[2], addr_204_4, wires_818_5,addr_818_5);

wire[3:0] wires_819_5;

wire[27:0] addr_819_5;

Selector_2 s819_5(wires_204_4[3], addr_204_4, wires_819_5,addr_819_5);

wire[3:0] wires_820_5;

wire[27:0] addr_820_5;

Selector_2 s820_5(wires_205_4[0], addr_205_4, wires_820_5,addr_820_5);

wire[3:0] wires_821_5;

wire[27:0] addr_821_5;

Selector_2 s821_5(wires_205_4[1], addr_205_4, wires_821_5,addr_821_5);

wire[3:0] wires_822_5;

wire[27:0] addr_822_5;

Selector_2 s822_5(wires_205_4[2], addr_205_4, wires_822_5,addr_822_5);

wire[3:0] wires_823_5;

wire[27:0] addr_823_5;

Selector_2 s823_5(wires_205_4[3], addr_205_4, wires_823_5,addr_823_5);

wire[3:0] wires_824_5;

wire[27:0] addr_824_5;

Selector_2 s824_5(wires_206_4[0], addr_206_4, wires_824_5,addr_824_5);

wire[3:0] wires_825_5;

wire[27:0] addr_825_5;

Selector_2 s825_5(wires_206_4[1], addr_206_4, wires_825_5,addr_825_5);

wire[3:0] wires_826_5;

wire[27:0] addr_826_5;

Selector_2 s826_5(wires_206_4[2], addr_206_4, wires_826_5,addr_826_5);

wire[3:0] wires_827_5;

wire[27:0] addr_827_5;

Selector_2 s827_5(wires_206_4[3], addr_206_4, wires_827_5,addr_827_5);

wire[3:0] wires_828_5;

wire[27:0] addr_828_5;

Selector_2 s828_5(wires_207_4[0], addr_207_4, wires_828_5,addr_828_5);

wire[3:0] wires_829_5;

wire[27:0] addr_829_5;

Selector_2 s829_5(wires_207_4[1], addr_207_4, wires_829_5,addr_829_5);

wire[3:0] wires_830_5;

wire[27:0] addr_830_5;

Selector_2 s830_5(wires_207_4[2], addr_207_4, wires_830_5,addr_830_5);

wire[3:0] wires_831_5;

wire[27:0] addr_831_5;

Selector_2 s831_5(wires_207_4[3], addr_207_4, wires_831_5,addr_831_5);

wire[3:0] wires_832_5;

wire[27:0] addr_832_5;

Selector_2 s832_5(wires_208_4[0], addr_208_4, wires_832_5,addr_832_5);

wire[3:0] wires_833_5;

wire[27:0] addr_833_5;

Selector_2 s833_5(wires_208_4[1], addr_208_4, wires_833_5,addr_833_5);

wire[3:0] wires_834_5;

wire[27:0] addr_834_5;

Selector_2 s834_5(wires_208_4[2], addr_208_4, wires_834_5,addr_834_5);

wire[3:0] wires_835_5;

wire[27:0] addr_835_5;

Selector_2 s835_5(wires_208_4[3], addr_208_4, wires_835_5,addr_835_5);

wire[3:0] wires_836_5;

wire[27:0] addr_836_5;

Selector_2 s836_5(wires_209_4[0], addr_209_4, wires_836_5,addr_836_5);

wire[3:0] wires_837_5;

wire[27:0] addr_837_5;

Selector_2 s837_5(wires_209_4[1], addr_209_4, wires_837_5,addr_837_5);

wire[3:0] wires_838_5;

wire[27:0] addr_838_5;

Selector_2 s838_5(wires_209_4[2], addr_209_4, wires_838_5,addr_838_5);

wire[3:0] wires_839_5;

wire[27:0] addr_839_5;

Selector_2 s839_5(wires_209_4[3], addr_209_4, wires_839_5,addr_839_5);

wire[3:0] wires_840_5;

wire[27:0] addr_840_5;

Selector_2 s840_5(wires_210_4[0], addr_210_4, wires_840_5,addr_840_5);

wire[3:0] wires_841_5;

wire[27:0] addr_841_5;

Selector_2 s841_5(wires_210_4[1], addr_210_4, wires_841_5,addr_841_5);

wire[3:0] wires_842_5;

wire[27:0] addr_842_5;

Selector_2 s842_5(wires_210_4[2], addr_210_4, wires_842_5,addr_842_5);

wire[3:0] wires_843_5;

wire[27:0] addr_843_5;

Selector_2 s843_5(wires_210_4[3], addr_210_4, wires_843_5,addr_843_5);

wire[3:0] wires_844_5;

wire[27:0] addr_844_5;

Selector_2 s844_5(wires_211_4[0], addr_211_4, wires_844_5,addr_844_5);

wire[3:0] wires_845_5;

wire[27:0] addr_845_5;

Selector_2 s845_5(wires_211_4[1], addr_211_4, wires_845_5,addr_845_5);

wire[3:0] wires_846_5;

wire[27:0] addr_846_5;

Selector_2 s846_5(wires_211_4[2], addr_211_4, wires_846_5,addr_846_5);

wire[3:0] wires_847_5;

wire[27:0] addr_847_5;

Selector_2 s847_5(wires_211_4[3], addr_211_4, wires_847_5,addr_847_5);

wire[3:0] wires_848_5;

wire[27:0] addr_848_5;

Selector_2 s848_5(wires_212_4[0], addr_212_4, wires_848_5,addr_848_5);

wire[3:0] wires_849_5;

wire[27:0] addr_849_5;

Selector_2 s849_5(wires_212_4[1], addr_212_4, wires_849_5,addr_849_5);

wire[3:0] wires_850_5;

wire[27:0] addr_850_5;

Selector_2 s850_5(wires_212_4[2], addr_212_4, wires_850_5,addr_850_5);

wire[3:0] wires_851_5;

wire[27:0] addr_851_5;

Selector_2 s851_5(wires_212_4[3], addr_212_4, wires_851_5,addr_851_5);

wire[3:0] wires_852_5;

wire[27:0] addr_852_5;

Selector_2 s852_5(wires_213_4[0], addr_213_4, wires_852_5,addr_852_5);

wire[3:0] wires_853_5;

wire[27:0] addr_853_5;

Selector_2 s853_5(wires_213_4[1], addr_213_4, wires_853_5,addr_853_5);

wire[3:0] wires_854_5;

wire[27:0] addr_854_5;

Selector_2 s854_5(wires_213_4[2], addr_213_4, wires_854_5,addr_854_5);

wire[3:0] wires_855_5;

wire[27:0] addr_855_5;

Selector_2 s855_5(wires_213_4[3], addr_213_4, wires_855_5,addr_855_5);

wire[3:0] wires_856_5;

wire[27:0] addr_856_5;

Selector_2 s856_5(wires_214_4[0], addr_214_4, wires_856_5,addr_856_5);

wire[3:0] wires_857_5;

wire[27:0] addr_857_5;

Selector_2 s857_5(wires_214_4[1], addr_214_4, wires_857_5,addr_857_5);

wire[3:0] wires_858_5;

wire[27:0] addr_858_5;

Selector_2 s858_5(wires_214_4[2], addr_214_4, wires_858_5,addr_858_5);

wire[3:0] wires_859_5;

wire[27:0] addr_859_5;

Selector_2 s859_5(wires_214_4[3], addr_214_4, wires_859_5,addr_859_5);

wire[3:0] wires_860_5;

wire[27:0] addr_860_5;

Selector_2 s860_5(wires_215_4[0], addr_215_4, wires_860_5,addr_860_5);

wire[3:0] wires_861_5;

wire[27:0] addr_861_5;

Selector_2 s861_5(wires_215_4[1], addr_215_4, wires_861_5,addr_861_5);

wire[3:0] wires_862_5;

wire[27:0] addr_862_5;

Selector_2 s862_5(wires_215_4[2], addr_215_4, wires_862_5,addr_862_5);

wire[3:0] wires_863_5;

wire[27:0] addr_863_5;

Selector_2 s863_5(wires_215_4[3], addr_215_4, wires_863_5,addr_863_5);

wire[3:0] wires_864_5;

wire[27:0] addr_864_5;

Selector_2 s864_5(wires_216_4[0], addr_216_4, wires_864_5,addr_864_5);

wire[3:0] wires_865_5;

wire[27:0] addr_865_5;

Selector_2 s865_5(wires_216_4[1], addr_216_4, wires_865_5,addr_865_5);

wire[3:0] wires_866_5;

wire[27:0] addr_866_5;

Selector_2 s866_5(wires_216_4[2], addr_216_4, wires_866_5,addr_866_5);

wire[3:0] wires_867_5;

wire[27:0] addr_867_5;

Selector_2 s867_5(wires_216_4[3], addr_216_4, wires_867_5,addr_867_5);

wire[3:0] wires_868_5;

wire[27:0] addr_868_5;

Selector_2 s868_5(wires_217_4[0], addr_217_4, wires_868_5,addr_868_5);

wire[3:0] wires_869_5;

wire[27:0] addr_869_5;

Selector_2 s869_5(wires_217_4[1], addr_217_4, wires_869_5,addr_869_5);

wire[3:0] wires_870_5;

wire[27:0] addr_870_5;

Selector_2 s870_5(wires_217_4[2], addr_217_4, wires_870_5,addr_870_5);

wire[3:0] wires_871_5;

wire[27:0] addr_871_5;

Selector_2 s871_5(wires_217_4[3], addr_217_4, wires_871_5,addr_871_5);

wire[3:0] wires_872_5;

wire[27:0] addr_872_5;

Selector_2 s872_5(wires_218_4[0], addr_218_4, wires_872_5,addr_872_5);

wire[3:0] wires_873_5;

wire[27:0] addr_873_5;

Selector_2 s873_5(wires_218_4[1], addr_218_4, wires_873_5,addr_873_5);

wire[3:0] wires_874_5;

wire[27:0] addr_874_5;

Selector_2 s874_5(wires_218_4[2], addr_218_4, wires_874_5,addr_874_5);

wire[3:0] wires_875_5;

wire[27:0] addr_875_5;

Selector_2 s875_5(wires_218_4[3], addr_218_4, wires_875_5,addr_875_5);

wire[3:0] wires_876_5;

wire[27:0] addr_876_5;

Selector_2 s876_5(wires_219_4[0], addr_219_4, wires_876_5,addr_876_5);

wire[3:0] wires_877_5;

wire[27:0] addr_877_5;

Selector_2 s877_5(wires_219_4[1], addr_219_4, wires_877_5,addr_877_5);

wire[3:0] wires_878_5;

wire[27:0] addr_878_5;

Selector_2 s878_5(wires_219_4[2], addr_219_4, wires_878_5,addr_878_5);

wire[3:0] wires_879_5;

wire[27:0] addr_879_5;

Selector_2 s879_5(wires_219_4[3], addr_219_4, wires_879_5,addr_879_5);

wire[3:0] wires_880_5;

wire[27:0] addr_880_5;

Selector_2 s880_5(wires_220_4[0], addr_220_4, wires_880_5,addr_880_5);

wire[3:0] wires_881_5;

wire[27:0] addr_881_5;

Selector_2 s881_5(wires_220_4[1], addr_220_4, wires_881_5,addr_881_5);

wire[3:0] wires_882_5;

wire[27:0] addr_882_5;

Selector_2 s882_5(wires_220_4[2], addr_220_4, wires_882_5,addr_882_5);

wire[3:0] wires_883_5;

wire[27:0] addr_883_5;

Selector_2 s883_5(wires_220_4[3], addr_220_4, wires_883_5,addr_883_5);

wire[3:0] wires_884_5;

wire[27:0] addr_884_5;

Selector_2 s884_5(wires_221_4[0], addr_221_4, wires_884_5,addr_884_5);

wire[3:0] wires_885_5;

wire[27:0] addr_885_5;

Selector_2 s885_5(wires_221_4[1], addr_221_4, wires_885_5,addr_885_5);

wire[3:0] wires_886_5;

wire[27:0] addr_886_5;

Selector_2 s886_5(wires_221_4[2], addr_221_4, wires_886_5,addr_886_5);

wire[3:0] wires_887_5;

wire[27:0] addr_887_5;

Selector_2 s887_5(wires_221_4[3], addr_221_4, wires_887_5,addr_887_5);

wire[3:0] wires_888_5;

wire[27:0] addr_888_5;

Selector_2 s888_5(wires_222_4[0], addr_222_4, wires_888_5,addr_888_5);

wire[3:0] wires_889_5;

wire[27:0] addr_889_5;

Selector_2 s889_5(wires_222_4[1], addr_222_4, wires_889_5,addr_889_5);

wire[3:0] wires_890_5;

wire[27:0] addr_890_5;

Selector_2 s890_5(wires_222_4[2], addr_222_4, wires_890_5,addr_890_5);

wire[3:0] wires_891_5;

wire[27:0] addr_891_5;

Selector_2 s891_5(wires_222_4[3], addr_222_4, wires_891_5,addr_891_5);

wire[3:0] wires_892_5;

wire[27:0] addr_892_5;

Selector_2 s892_5(wires_223_4[0], addr_223_4, wires_892_5,addr_892_5);

wire[3:0] wires_893_5;

wire[27:0] addr_893_5;

Selector_2 s893_5(wires_223_4[1], addr_223_4, wires_893_5,addr_893_5);

wire[3:0] wires_894_5;

wire[27:0] addr_894_5;

Selector_2 s894_5(wires_223_4[2], addr_223_4, wires_894_5,addr_894_5);

wire[3:0] wires_895_5;

wire[27:0] addr_895_5;

Selector_2 s895_5(wires_223_4[3], addr_223_4, wires_895_5,addr_895_5);

wire[3:0] wires_896_5;

wire[27:0] addr_896_5;

Selector_2 s896_5(wires_224_4[0], addr_224_4, wires_896_5,addr_896_5);

wire[3:0] wires_897_5;

wire[27:0] addr_897_5;

Selector_2 s897_5(wires_224_4[1], addr_224_4, wires_897_5,addr_897_5);

wire[3:0] wires_898_5;

wire[27:0] addr_898_5;

Selector_2 s898_5(wires_224_4[2], addr_224_4, wires_898_5,addr_898_5);

wire[3:0] wires_899_5;

wire[27:0] addr_899_5;

Selector_2 s899_5(wires_224_4[3], addr_224_4, wires_899_5,addr_899_5);

wire[3:0] wires_900_5;

wire[27:0] addr_900_5;

Selector_2 s900_5(wires_225_4[0], addr_225_4, wires_900_5,addr_900_5);

wire[3:0] wires_901_5;

wire[27:0] addr_901_5;

Selector_2 s901_5(wires_225_4[1], addr_225_4, wires_901_5,addr_901_5);

wire[3:0] wires_902_5;

wire[27:0] addr_902_5;

Selector_2 s902_5(wires_225_4[2], addr_225_4, wires_902_5,addr_902_5);

wire[3:0] wires_903_5;

wire[27:0] addr_903_5;

Selector_2 s903_5(wires_225_4[3], addr_225_4, wires_903_5,addr_903_5);

wire[3:0] wires_904_5;

wire[27:0] addr_904_5;

Selector_2 s904_5(wires_226_4[0], addr_226_4, wires_904_5,addr_904_5);

wire[3:0] wires_905_5;

wire[27:0] addr_905_5;

Selector_2 s905_5(wires_226_4[1], addr_226_4, wires_905_5,addr_905_5);

wire[3:0] wires_906_5;

wire[27:0] addr_906_5;

Selector_2 s906_5(wires_226_4[2], addr_226_4, wires_906_5,addr_906_5);

wire[3:0] wires_907_5;

wire[27:0] addr_907_5;

Selector_2 s907_5(wires_226_4[3], addr_226_4, wires_907_5,addr_907_5);

wire[3:0] wires_908_5;

wire[27:0] addr_908_5;

Selector_2 s908_5(wires_227_4[0], addr_227_4, wires_908_5,addr_908_5);

wire[3:0] wires_909_5;

wire[27:0] addr_909_5;

Selector_2 s909_5(wires_227_4[1], addr_227_4, wires_909_5,addr_909_5);

wire[3:0] wires_910_5;

wire[27:0] addr_910_5;

Selector_2 s910_5(wires_227_4[2], addr_227_4, wires_910_5,addr_910_5);

wire[3:0] wires_911_5;

wire[27:0] addr_911_5;

Selector_2 s911_5(wires_227_4[3], addr_227_4, wires_911_5,addr_911_5);

wire[3:0] wires_912_5;

wire[27:0] addr_912_5;

Selector_2 s912_5(wires_228_4[0], addr_228_4, wires_912_5,addr_912_5);

wire[3:0] wires_913_5;

wire[27:0] addr_913_5;

Selector_2 s913_5(wires_228_4[1], addr_228_4, wires_913_5,addr_913_5);

wire[3:0] wires_914_5;

wire[27:0] addr_914_5;

Selector_2 s914_5(wires_228_4[2], addr_228_4, wires_914_5,addr_914_5);

wire[3:0] wires_915_5;

wire[27:0] addr_915_5;

Selector_2 s915_5(wires_228_4[3], addr_228_4, wires_915_5,addr_915_5);

wire[3:0] wires_916_5;

wire[27:0] addr_916_5;

Selector_2 s916_5(wires_229_4[0], addr_229_4, wires_916_5,addr_916_5);

wire[3:0] wires_917_5;

wire[27:0] addr_917_5;

Selector_2 s917_5(wires_229_4[1], addr_229_4, wires_917_5,addr_917_5);

wire[3:0] wires_918_5;

wire[27:0] addr_918_5;

Selector_2 s918_5(wires_229_4[2], addr_229_4, wires_918_5,addr_918_5);

wire[3:0] wires_919_5;

wire[27:0] addr_919_5;

Selector_2 s919_5(wires_229_4[3], addr_229_4, wires_919_5,addr_919_5);

wire[3:0] wires_920_5;

wire[27:0] addr_920_5;

Selector_2 s920_5(wires_230_4[0], addr_230_4, wires_920_5,addr_920_5);

wire[3:0] wires_921_5;

wire[27:0] addr_921_5;

Selector_2 s921_5(wires_230_4[1], addr_230_4, wires_921_5,addr_921_5);

wire[3:0] wires_922_5;

wire[27:0] addr_922_5;

Selector_2 s922_5(wires_230_4[2], addr_230_4, wires_922_5,addr_922_5);

wire[3:0] wires_923_5;

wire[27:0] addr_923_5;

Selector_2 s923_5(wires_230_4[3], addr_230_4, wires_923_5,addr_923_5);

wire[3:0] wires_924_5;

wire[27:0] addr_924_5;

Selector_2 s924_5(wires_231_4[0], addr_231_4, wires_924_5,addr_924_5);

wire[3:0] wires_925_5;

wire[27:0] addr_925_5;

Selector_2 s925_5(wires_231_4[1], addr_231_4, wires_925_5,addr_925_5);

wire[3:0] wires_926_5;

wire[27:0] addr_926_5;

Selector_2 s926_5(wires_231_4[2], addr_231_4, wires_926_5,addr_926_5);

wire[3:0] wires_927_5;

wire[27:0] addr_927_5;

Selector_2 s927_5(wires_231_4[3], addr_231_4, wires_927_5,addr_927_5);

wire[3:0] wires_928_5;

wire[27:0] addr_928_5;

Selector_2 s928_5(wires_232_4[0], addr_232_4, wires_928_5,addr_928_5);

wire[3:0] wires_929_5;

wire[27:0] addr_929_5;

Selector_2 s929_5(wires_232_4[1], addr_232_4, wires_929_5,addr_929_5);

wire[3:0] wires_930_5;

wire[27:0] addr_930_5;

Selector_2 s930_5(wires_232_4[2], addr_232_4, wires_930_5,addr_930_5);

wire[3:0] wires_931_5;

wire[27:0] addr_931_5;

Selector_2 s931_5(wires_232_4[3], addr_232_4, wires_931_5,addr_931_5);

wire[3:0] wires_932_5;

wire[27:0] addr_932_5;

Selector_2 s932_5(wires_233_4[0], addr_233_4, wires_932_5,addr_932_5);

wire[3:0] wires_933_5;

wire[27:0] addr_933_5;

Selector_2 s933_5(wires_233_4[1], addr_233_4, wires_933_5,addr_933_5);

wire[3:0] wires_934_5;

wire[27:0] addr_934_5;

Selector_2 s934_5(wires_233_4[2], addr_233_4, wires_934_5,addr_934_5);

wire[3:0] wires_935_5;

wire[27:0] addr_935_5;

Selector_2 s935_5(wires_233_4[3], addr_233_4, wires_935_5,addr_935_5);

wire[3:0] wires_936_5;

wire[27:0] addr_936_5;

Selector_2 s936_5(wires_234_4[0], addr_234_4, wires_936_5,addr_936_5);

wire[3:0] wires_937_5;

wire[27:0] addr_937_5;

Selector_2 s937_5(wires_234_4[1], addr_234_4, wires_937_5,addr_937_5);

wire[3:0] wires_938_5;

wire[27:0] addr_938_5;

Selector_2 s938_5(wires_234_4[2], addr_234_4, wires_938_5,addr_938_5);

wire[3:0] wires_939_5;

wire[27:0] addr_939_5;

Selector_2 s939_5(wires_234_4[3], addr_234_4, wires_939_5,addr_939_5);

wire[3:0] wires_940_5;

wire[27:0] addr_940_5;

Selector_2 s940_5(wires_235_4[0], addr_235_4, wires_940_5,addr_940_5);

wire[3:0] wires_941_5;

wire[27:0] addr_941_5;

Selector_2 s941_5(wires_235_4[1], addr_235_4, wires_941_5,addr_941_5);

wire[3:0] wires_942_5;

wire[27:0] addr_942_5;

Selector_2 s942_5(wires_235_4[2], addr_235_4, wires_942_5,addr_942_5);

wire[3:0] wires_943_5;

wire[27:0] addr_943_5;

Selector_2 s943_5(wires_235_4[3], addr_235_4, wires_943_5,addr_943_5);

wire[3:0] wires_944_5;

wire[27:0] addr_944_5;

Selector_2 s944_5(wires_236_4[0], addr_236_4, wires_944_5,addr_944_5);

wire[3:0] wires_945_5;

wire[27:0] addr_945_5;

Selector_2 s945_5(wires_236_4[1], addr_236_4, wires_945_5,addr_945_5);

wire[3:0] wires_946_5;

wire[27:0] addr_946_5;

Selector_2 s946_5(wires_236_4[2], addr_236_4, wires_946_5,addr_946_5);

wire[3:0] wires_947_5;

wire[27:0] addr_947_5;

Selector_2 s947_5(wires_236_4[3], addr_236_4, wires_947_5,addr_947_5);

wire[3:0] wires_948_5;

wire[27:0] addr_948_5;

Selector_2 s948_5(wires_237_4[0], addr_237_4, wires_948_5,addr_948_5);

wire[3:0] wires_949_5;

wire[27:0] addr_949_5;

Selector_2 s949_5(wires_237_4[1], addr_237_4, wires_949_5,addr_949_5);

wire[3:0] wires_950_5;

wire[27:0] addr_950_5;

Selector_2 s950_5(wires_237_4[2], addr_237_4, wires_950_5,addr_950_5);

wire[3:0] wires_951_5;

wire[27:0] addr_951_5;

Selector_2 s951_5(wires_237_4[3], addr_237_4, wires_951_5,addr_951_5);

wire[3:0] wires_952_5;

wire[27:0] addr_952_5;

Selector_2 s952_5(wires_238_4[0], addr_238_4, wires_952_5,addr_952_5);

wire[3:0] wires_953_5;

wire[27:0] addr_953_5;

Selector_2 s953_5(wires_238_4[1], addr_238_4, wires_953_5,addr_953_5);

wire[3:0] wires_954_5;

wire[27:0] addr_954_5;

Selector_2 s954_5(wires_238_4[2], addr_238_4, wires_954_5,addr_954_5);

wire[3:0] wires_955_5;

wire[27:0] addr_955_5;

Selector_2 s955_5(wires_238_4[3], addr_238_4, wires_955_5,addr_955_5);

wire[3:0] wires_956_5;

wire[27:0] addr_956_5;

Selector_2 s956_5(wires_239_4[0], addr_239_4, wires_956_5,addr_956_5);

wire[3:0] wires_957_5;

wire[27:0] addr_957_5;

Selector_2 s957_5(wires_239_4[1], addr_239_4, wires_957_5,addr_957_5);

wire[3:0] wires_958_5;

wire[27:0] addr_958_5;

Selector_2 s958_5(wires_239_4[2], addr_239_4, wires_958_5,addr_958_5);

wire[3:0] wires_959_5;

wire[27:0] addr_959_5;

Selector_2 s959_5(wires_239_4[3], addr_239_4, wires_959_5,addr_959_5);

wire[3:0] wires_960_5;

wire[27:0] addr_960_5;

Selector_2 s960_5(wires_240_4[0], addr_240_4, wires_960_5,addr_960_5);

wire[3:0] wires_961_5;

wire[27:0] addr_961_5;

Selector_2 s961_5(wires_240_4[1], addr_240_4, wires_961_5,addr_961_5);

wire[3:0] wires_962_5;

wire[27:0] addr_962_5;

Selector_2 s962_5(wires_240_4[2], addr_240_4, wires_962_5,addr_962_5);

wire[3:0] wires_963_5;

wire[27:0] addr_963_5;

Selector_2 s963_5(wires_240_4[3], addr_240_4, wires_963_5,addr_963_5);

wire[3:0] wires_964_5;

wire[27:0] addr_964_5;

Selector_2 s964_5(wires_241_4[0], addr_241_4, wires_964_5,addr_964_5);

wire[3:0] wires_965_5;

wire[27:0] addr_965_5;

Selector_2 s965_5(wires_241_4[1], addr_241_4, wires_965_5,addr_965_5);

wire[3:0] wires_966_5;

wire[27:0] addr_966_5;

Selector_2 s966_5(wires_241_4[2], addr_241_4, wires_966_5,addr_966_5);

wire[3:0] wires_967_5;

wire[27:0] addr_967_5;

Selector_2 s967_5(wires_241_4[3], addr_241_4, wires_967_5,addr_967_5);

wire[3:0] wires_968_5;

wire[27:0] addr_968_5;

Selector_2 s968_5(wires_242_4[0], addr_242_4, wires_968_5,addr_968_5);

wire[3:0] wires_969_5;

wire[27:0] addr_969_5;

Selector_2 s969_5(wires_242_4[1], addr_242_4, wires_969_5,addr_969_5);

wire[3:0] wires_970_5;

wire[27:0] addr_970_5;

Selector_2 s970_5(wires_242_4[2], addr_242_4, wires_970_5,addr_970_5);

wire[3:0] wires_971_5;

wire[27:0] addr_971_5;

Selector_2 s971_5(wires_242_4[3], addr_242_4, wires_971_5,addr_971_5);

wire[3:0] wires_972_5;

wire[27:0] addr_972_5;

Selector_2 s972_5(wires_243_4[0], addr_243_4, wires_972_5,addr_972_5);

wire[3:0] wires_973_5;

wire[27:0] addr_973_5;

Selector_2 s973_5(wires_243_4[1], addr_243_4, wires_973_5,addr_973_5);

wire[3:0] wires_974_5;

wire[27:0] addr_974_5;

Selector_2 s974_5(wires_243_4[2], addr_243_4, wires_974_5,addr_974_5);

wire[3:0] wires_975_5;

wire[27:0] addr_975_5;

Selector_2 s975_5(wires_243_4[3], addr_243_4, wires_975_5,addr_975_5);

wire[3:0] wires_976_5;

wire[27:0] addr_976_5;

Selector_2 s976_5(wires_244_4[0], addr_244_4, wires_976_5,addr_976_5);

wire[3:0] wires_977_5;

wire[27:0] addr_977_5;

Selector_2 s977_5(wires_244_4[1], addr_244_4, wires_977_5,addr_977_5);

wire[3:0] wires_978_5;

wire[27:0] addr_978_5;

Selector_2 s978_5(wires_244_4[2], addr_244_4, wires_978_5,addr_978_5);

wire[3:0] wires_979_5;

wire[27:0] addr_979_5;

Selector_2 s979_5(wires_244_4[3], addr_244_4, wires_979_5,addr_979_5);

wire[3:0] wires_980_5;

wire[27:0] addr_980_5;

Selector_2 s980_5(wires_245_4[0], addr_245_4, wires_980_5,addr_980_5);

wire[3:0] wires_981_5;

wire[27:0] addr_981_5;

Selector_2 s981_5(wires_245_4[1], addr_245_4, wires_981_5,addr_981_5);

wire[3:0] wires_982_5;

wire[27:0] addr_982_5;

Selector_2 s982_5(wires_245_4[2], addr_245_4, wires_982_5,addr_982_5);

wire[3:0] wires_983_5;

wire[27:0] addr_983_5;

Selector_2 s983_5(wires_245_4[3], addr_245_4, wires_983_5,addr_983_5);

wire[3:0] wires_984_5;

wire[27:0] addr_984_5;

Selector_2 s984_5(wires_246_4[0], addr_246_4, wires_984_5,addr_984_5);

wire[3:0] wires_985_5;

wire[27:0] addr_985_5;

Selector_2 s985_5(wires_246_4[1], addr_246_4, wires_985_5,addr_985_5);

wire[3:0] wires_986_5;

wire[27:0] addr_986_5;

Selector_2 s986_5(wires_246_4[2], addr_246_4, wires_986_5,addr_986_5);

wire[3:0] wires_987_5;

wire[27:0] addr_987_5;

Selector_2 s987_5(wires_246_4[3], addr_246_4, wires_987_5,addr_987_5);

wire[3:0] wires_988_5;

wire[27:0] addr_988_5;

Selector_2 s988_5(wires_247_4[0], addr_247_4, wires_988_5,addr_988_5);

wire[3:0] wires_989_5;

wire[27:0] addr_989_5;

Selector_2 s989_5(wires_247_4[1], addr_247_4, wires_989_5,addr_989_5);

wire[3:0] wires_990_5;

wire[27:0] addr_990_5;

Selector_2 s990_5(wires_247_4[2], addr_247_4, wires_990_5,addr_990_5);

wire[3:0] wires_991_5;

wire[27:0] addr_991_5;

Selector_2 s991_5(wires_247_4[3], addr_247_4, wires_991_5,addr_991_5);

wire[3:0] wires_992_5;

wire[27:0] addr_992_5;

Selector_2 s992_5(wires_248_4[0], addr_248_4, wires_992_5,addr_992_5);

wire[3:0] wires_993_5;

wire[27:0] addr_993_5;

Selector_2 s993_5(wires_248_4[1], addr_248_4, wires_993_5,addr_993_5);

wire[3:0] wires_994_5;

wire[27:0] addr_994_5;

Selector_2 s994_5(wires_248_4[2], addr_248_4, wires_994_5,addr_994_5);

wire[3:0] wires_995_5;

wire[27:0] addr_995_5;

Selector_2 s995_5(wires_248_4[3], addr_248_4, wires_995_5,addr_995_5);

wire[3:0] wires_996_5;

wire[27:0] addr_996_5;

Selector_2 s996_5(wires_249_4[0], addr_249_4, wires_996_5,addr_996_5);

wire[3:0] wires_997_5;

wire[27:0] addr_997_5;

Selector_2 s997_5(wires_249_4[1], addr_249_4, wires_997_5,addr_997_5);

wire[3:0] wires_998_5;

wire[27:0] addr_998_5;

Selector_2 s998_5(wires_249_4[2], addr_249_4, wires_998_5,addr_998_5);

wire[3:0] wires_999_5;

wire[27:0] addr_999_5;

Selector_2 s999_5(wires_249_4[3], addr_249_4, wires_999_5,addr_999_5);

wire[3:0] wires_1000_5;

wire[27:0] addr_1000_5;

Selector_2 s1000_5(wires_250_4[0], addr_250_4, wires_1000_5,addr_1000_5);

wire[3:0] wires_1001_5;

wire[27:0] addr_1001_5;

Selector_2 s1001_5(wires_250_4[1], addr_250_4, wires_1001_5,addr_1001_5);

wire[3:0] wires_1002_5;

wire[27:0] addr_1002_5;

Selector_2 s1002_5(wires_250_4[2], addr_250_4, wires_1002_5,addr_1002_5);

wire[3:0] wires_1003_5;

wire[27:0] addr_1003_5;

Selector_2 s1003_5(wires_250_4[3], addr_250_4, wires_1003_5,addr_1003_5);

wire[3:0] wires_1004_5;

wire[27:0] addr_1004_5;

Selector_2 s1004_5(wires_251_4[0], addr_251_4, wires_1004_5,addr_1004_5);

wire[3:0] wires_1005_5;

wire[27:0] addr_1005_5;

Selector_2 s1005_5(wires_251_4[1], addr_251_4, wires_1005_5,addr_1005_5);

wire[3:0] wires_1006_5;

wire[27:0] addr_1006_5;

Selector_2 s1006_5(wires_251_4[2], addr_251_4, wires_1006_5,addr_1006_5);

wire[3:0] wires_1007_5;

wire[27:0] addr_1007_5;

Selector_2 s1007_5(wires_251_4[3], addr_251_4, wires_1007_5,addr_1007_5);

wire[3:0] wires_1008_5;

wire[27:0] addr_1008_5;

Selector_2 s1008_5(wires_252_4[0], addr_252_4, wires_1008_5,addr_1008_5);

wire[3:0] wires_1009_5;

wire[27:0] addr_1009_5;

Selector_2 s1009_5(wires_252_4[1], addr_252_4, wires_1009_5,addr_1009_5);

wire[3:0] wires_1010_5;

wire[27:0] addr_1010_5;

Selector_2 s1010_5(wires_252_4[2], addr_252_4, wires_1010_5,addr_1010_5);

wire[3:0] wires_1011_5;

wire[27:0] addr_1011_5;

Selector_2 s1011_5(wires_252_4[3], addr_252_4, wires_1011_5,addr_1011_5);

wire[3:0] wires_1012_5;

wire[27:0] addr_1012_5;

Selector_2 s1012_5(wires_253_4[0], addr_253_4, wires_1012_5,addr_1012_5);

wire[3:0] wires_1013_5;

wire[27:0] addr_1013_5;

Selector_2 s1013_5(wires_253_4[1], addr_253_4, wires_1013_5,addr_1013_5);

wire[3:0] wires_1014_5;

wire[27:0] addr_1014_5;

Selector_2 s1014_5(wires_253_4[2], addr_253_4, wires_1014_5,addr_1014_5);

wire[3:0] wires_1015_5;

wire[27:0] addr_1015_5;

Selector_2 s1015_5(wires_253_4[3], addr_253_4, wires_1015_5,addr_1015_5);

wire[3:0] wires_1016_5;

wire[27:0] addr_1016_5;

Selector_2 s1016_5(wires_254_4[0], addr_254_4, wires_1016_5,addr_1016_5);

wire[3:0] wires_1017_5;

wire[27:0] addr_1017_5;

Selector_2 s1017_5(wires_254_4[1], addr_254_4, wires_1017_5,addr_1017_5);

wire[3:0] wires_1018_5;

wire[27:0] addr_1018_5;

Selector_2 s1018_5(wires_254_4[2], addr_254_4, wires_1018_5,addr_1018_5);

wire[3:0] wires_1019_5;

wire[27:0] addr_1019_5;

Selector_2 s1019_5(wires_254_4[3], addr_254_4, wires_1019_5,addr_1019_5);

wire[3:0] wires_1020_5;

wire[27:0] addr_1020_5;

Selector_2 s1020_5(wires_255_4[0], addr_255_4, wires_1020_5,addr_1020_5);

wire[3:0] wires_1021_5;

wire[27:0] addr_1021_5;

Selector_2 s1021_5(wires_255_4[1], addr_255_4, wires_1021_5,addr_1021_5);

wire[3:0] wires_1022_5;

wire[27:0] addr_1022_5;

Selector_2 s1022_5(wires_255_4[2], addr_255_4, wires_1022_5,addr_1022_5);

wire[3:0] wires_1023_5;

wire[27:0] addr_1023_5;

Selector_2 s1023_5(wires_255_4[3], addr_255_4, wires_1023_5,addr_1023_5);

wire[27:0] addr_0_6;

Selector_2 s0_6(wires_0_5[0], addr_0_5, addr_positional[3:0], addr_0_6);

wire[27:0] addr_1_6;

Selector_2 s1_6(wires_0_5[1], addr_0_5, addr_positional[7:4], addr_1_6);

wire[27:0] addr_2_6;

Selector_2 s2_6(wires_0_5[2], addr_0_5, addr_positional[11:8], addr_2_6);

wire[27:0] addr_3_6;

Selector_2 s3_6(wires_0_5[3], addr_0_5, addr_positional[15:12], addr_3_6);

wire[27:0] addr_4_6;

Selector_2 s4_6(wires_1_5[0], addr_1_5, addr_positional[19:16], addr_4_6);

wire[27:0] addr_5_6;

Selector_2 s5_6(wires_1_5[1], addr_1_5, addr_positional[23:20], addr_5_6);

wire[27:0] addr_6_6;

Selector_2 s6_6(wires_1_5[2], addr_1_5, addr_positional[27:24], addr_6_6);

wire[27:0] addr_7_6;

Selector_2 s7_6(wires_1_5[3], addr_1_5, addr_positional[31:28], addr_7_6);

wire[27:0] addr_8_6;

Selector_2 s8_6(wires_2_5[0], addr_2_5, addr_positional[35:32], addr_8_6);

wire[27:0] addr_9_6;

Selector_2 s9_6(wires_2_5[1], addr_2_5, addr_positional[39:36], addr_9_6);

wire[27:0] addr_10_6;

Selector_2 s10_6(wires_2_5[2], addr_2_5, addr_positional[43:40], addr_10_6);

wire[27:0] addr_11_6;

Selector_2 s11_6(wires_2_5[3], addr_2_5, addr_positional[47:44], addr_11_6);

wire[27:0] addr_12_6;

Selector_2 s12_6(wires_3_5[0], addr_3_5, addr_positional[51:48], addr_12_6);

wire[27:0] addr_13_6;

Selector_2 s13_6(wires_3_5[1], addr_3_5, addr_positional[55:52], addr_13_6);

wire[27:0] addr_14_6;

Selector_2 s14_6(wires_3_5[2], addr_3_5, addr_positional[59:56], addr_14_6);

wire[27:0] addr_15_6;

Selector_2 s15_6(wires_3_5[3], addr_3_5, addr_positional[63:60], addr_15_6);

wire[27:0] addr_16_6;

Selector_2 s16_6(wires_4_5[0], addr_4_5, addr_positional[67:64], addr_16_6);

wire[27:0] addr_17_6;

Selector_2 s17_6(wires_4_5[1], addr_4_5, addr_positional[71:68], addr_17_6);

wire[27:0] addr_18_6;

Selector_2 s18_6(wires_4_5[2], addr_4_5, addr_positional[75:72], addr_18_6);

wire[27:0] addr_19_6;

Selector_2 s19_6(wires_4_5[3], addr_4_5, addr_positional[79:76], addr_19_6);

wire[27:0] addr_20_6;

Selector_2 s20_6(wires_5_5[0], addr_5_5, addr_positional[83:80], addr_20_6);

wire[27:0] addr_21_6;

Selector_2 s21_6(wires_5_5[1], addr_5_5, addr_positional[87:84], addr_21_6);

wire[27:0] addr_22_6;

Selector_2 s22_6(wires_5_5[2], addr_5_5, addr_positional[91:88], addr_22_6);

wire[27:0] addr_23_6;

Selector_2 s23_6(wires_5_5[3], addr_5_5, addr_positional[95:92], addr_23_6);

wire[27:0] addr_24_6;

Selector_2 s24_6(wires_6_5[0], addr_6_5, addr_positional[99:96], addr_24_6);

wire[27:0] addr_25_6;

Selector_2 s25_6(wires_6_5[1], addr_6_5, addr_positional[103:100], addr_25_6);

wire[27:0] addr_26_6;

Selector_2 s26_6(wires_6_5[2], addr_6_5, addr_positional[107:104], addr_26_6);

wire[27:0] addr_27_6;

Selector_2 s27_6(wires_6_5[3], addr_6_5, addr_positional[111:108], addr_27_6);

wire[27:0] addr_28_6;

Selector_2 s28_6(wires_7_5[0], addr_7_5, addr_positional[115:112], addr_28_6);

wire[27:0] addr_29_6;

Selector_2 s29_6(wires_7_5[1], addr_7_5, addr_positional[119:116], addr_29_6);

wire[27:0] addr_30_6;

Selector_2 s30_6(wires_7_5[2], addr_7_5, addr_positional[123:120], addr_30_6);

wire[27:0] addr_31_6;

Selector_2 s31_6(wires_7_5[3], addr_7_5, addr_positional[127:124], addr_31_6);

wire[27:0] addr_32_6;

Selector_2 s32_6(wires_8_5[0], addr_8_5, addr_positional[131:128], addr_32_6);

wire[27:0] addr_33_6;

Selector_2 s33_6(wires_8_5[1], addr_8_5, addr_positional[135:132], addr_33_6);

wire[27:0] addr_34_6;

Selector_2 s34_6(wires_8_5[2], addr_8_5, addr_positional[139:136], addr_34_6);

wire[27:0] addr_35_6;

Selector_2 s35_6(wires_8_5[3], addr_8_5, addr_positional[143:140], addr_35_6);

wire[27:0] addr_36_6;

Selector_2 s36_6(wires_9_5[0], addr_9_5, addr_positional[147:144], addr_36_6);

wire[27:0] addr_37_6;

Selector_2 s37_6(wires_9_5[1], addr_9_5, addr_positional[151:148], addr_37_6);

wire[27:0] addr_38_6;

Selector_2 s38_6(wires_9_5[2], addr_9_5, addr_positional[155:152], addr_38_6);

wire[27:0] addr_39_6;

Selector_2 s39_6(wires_9_5[3], addr_9_5, addr_positional[159:156], addr_39_6);

wire[27:0] addr_40_6;

Selector_2 s40_6(wires_10_5[0], addr_10_5, addr_positional[163:160], addr_40_6);

wire[27:0] addr_41_6;

Selector_2 s41_6(wires_10_5[1], addr_10_5, addr_positional[167:164], addr_41_6);

wire[27:0] addr_42_6;

Selector_2 s42_6(wires_10_5[2], addr_10_5, addr_positional[171:168], addr_42_6);

wire[27:0] addr_43_6;

Selector_2 s43_6(wires_10_5[3], addr_10_5, addr_positional[175:172], addr_43_6);

wire[27:0] addr_44_6;

Selector_2 s44_6(wires_11_5[0], addr_11_5, addr_positional[179:176], addr_44_6);

wire[27:0] addr_45_6;

Selector_2 s45_6(wires_11_5[1], addr_11_5, addr_positional[183:180], addr_45_6);

wire[27:0] addr_46_6;

Selector_2 s46_6(wires_11_5[2], addr_11_5, addr_positional[187:184], addr_46_6);

wire[27:0] addr_47_6;

Selector_2 s47_6(wires_11_5[3], addr_11_5, addr_positional[191:188], addr_47_6);

wire[27:0] addr_48_6;

Selector_2 s48_6(wires_12_5[0], addr_12_5, addr_positional[195:192], addr_48_6);

wire[27:0] addr_49_6;

Selector_2 s49_6(wires_12_5[1], addr_12_5, addr_positional[199:196], addr_49_6);

wire[27:0] addr_50_6;

Selector_2 s50_6(wires_12_5[2], addr_12_5, addr_positional[203:200], addr_50_6);

wire[27:0] addr_51_6;

Selector_2 s51_6(wires_12_5[3], addr_12_5, addr_positional[207:204], addr_51_6);

wire[27:0] addr_52_6;

Selector_2 s52_6(wires_13_5[0], addr_13_5, addr_positional[211:208], addr_52_6);

wire[27:0] addr_53_6;

Selector_2 s53_6(wires_13_5[1], addr_13_5, addr_positional[215:212], addr_53_6);

wire[27:0] addr_54_6;

Selector_2 s54_6(wires_13_5[2], addr_13_5, addr_positional[219:216], addr_54_6);

wire[27:0] addr_55_6;

Selector_2 s55_6(wires_13_5[3], addr_13_5, addr_positional[223:220], addr_55_6);

wire[27:0] addr_56_6;

Selector_2 s56_6(wires_14_5[0], addr_14_5, addr_positional[227:224], addr_56_6);

wire[27:0] addr_57_6;

Selector_2 s57_6(wires_14_5[1], addr_14_5, addr_positional[231:228], addr_57_6);

wire[27:0] addr_58_6;

Selector_2 s58_6(wires_14_5[2], addr_14_5, addr_positional[235:232], addr_58_6);

wire[27:0] addr_59_6;

Selector_2 s59_6(wires_14_5[3], addr_14_5, addr_positional[239:236], addr_59_6);

wire[27:0] addr_60_6;

Selector_2 s60_6(wires_15_5[0], addr_15_5, addr_positional[243:240], addr_60_6);

wire[27:0] addr_61_6;

Selector_2 s61_6(wires_15_5[1], addr_15_5, addr_positional[247:244], addr_61_6);

wire[27:0] addr_62_6;

Selector_2 s62_6(wires_15_5[2], addr_15_5, addr_positional[251:248], addr_62_6);

wire[27:0] addr_63_6;

Selector_2 s63_6(wires_15_5[3], addr_15_5, addr_positional[255:252], addr_63_6);

wire[27:0] addr_64_6;

Selector_2 s64_6(wires_16_5[0], addr_16_5, addr_positional[259:256], addr_64_6);

wire[27:0] addr_65_6;

Selector_2 s65_6(wires_16_5[1], addr_16_5, addr_positional[263:260], addr_65_6);

wire[27:0] addr_66_6;

Selector_2 s66_6(wires_16_5[2], addr_16_5, addr_positional[267:264], addr_66_6);

wire[27:0] addr_67_6;

Selector_2 s67_6(wires_16_5[3], addr_16_5, addr_positional[271:268], addr_67_6);

wire[27:0] addr_68_6;

Selector_2 s68_6(wires_17_5[0], addr_17_5, addr_positional[275:272], addr_68_6);

wire[27:0] addr_69_6;

Selector_2 s69_6(wires_17_5[1], addr_17_5, addr_positional[279:276], addr_69_6);

wire[27:0] addr_70_6;

Selector_2 s70_6(wires_17_5[2], addr_17_5, addr_positional[283:280], addr_70_6);

wire[27:0] addr_71_6;

Selector_2 s71_6(wires_17_5[3], addr_17_5, addr_positional[287:284], addr_71_6);

wire[27:0] addr_72_6;

Selector_2 s72_6(wires_18_5[0], addr_18_5, addr_positional[291:288], addr_72_6);

wire[27:0] addr_73_6;

Selector_2 s73_6(wires_18_5[1], addr_18_5, addr_positional[295:292], addr_73_6);

wire[27:0] addr_74_6;

Selector_2 s74_6(wires_18_5[2], addr_18_5, addr_positional[299:296], addr_74_6);

wire[27:0] addr_75_6;

Selector_2 s75_6(wires_18_5[3], addr_18_5, addr_positional[303:300], addr_75_6);

wire[27:0] addr_76_6;

Selector_2 s76_6(wires_19_5[0], addr_19_5, addr_positional[307:304], addr_76_6);

wire[27:0] addr_77_6;

Selector_2 s77_6(wires_19_5[1], addr_19_5, addr_positional[311:308], addr_77_6);

wire[27:0] addr_78_6;

Selector_2 s78_6(wires_19_5[2], addr_19_5, addr_positional[315:312], addr_78_6);

wire[27:0] addr_79_6;

Selector_2 s79_6(wires_19_5[3], addr_19_5, addr_positional[319:316], addr_79_6);

wire[27:0] addr_80_6;

Selector_2 s80_6(wires_20_5[0], addr_20_5, addr_positional[323:320], addr_80_6);

wire[27:0] addr_81_6;

Selector_2 s81_6(wires_20_5[1], addr_20_5, addr_positional[327:324], addr_81_6);

wire[27:0] addr_82_6;

Selector_2 s82_6(wires_20_5[2], addr_20_5, addr_positional[331:328], addr_82_6);

wire[27:0] addr_83_6;

Selector_2 s83_6(wires_20_5[3], addr_20_5, addr_positional[335:332], addr_83_6);

wire[27:0] addr_84_6;

Selector_2 s84_6(wires_21_5[0], addr_21_5, addr_positional[339:336], addr_84_6);

wire[27:0] addr_85_6;

Selector_2 s85_6(wires_21_5[1], addr_21_5, addr_positional[343:340], addr_85_6);

wire[27:0] addr_86_6;

Selector_2 s86_6(wires_21_5[2], addr_21_5, addr_positional[347:344], addr_86_6);

wire[27:0] addr_87_6;

Selector_2 s87_6(wires_21_5[3], addr_21_5, addr_positional[351:348], addr_87_6);

wire[27:0] addr_88_6;

Selector_2 s88_6(wires_22_5[0], addr_22_5, addr_positional[355:352], addr_88_6);

wire[27:0] addr_89_6;

Selector_2 s89_6(wires_22_5[1], addr_22_5, addr_positional[359:356], addr_89_6);

wire[27:0] addr_90_6;

Selector_2 s90_6(wires_22_5[2], addr_22_5, addr_positional[363:360], addr_90_6);

wire[27:0] addr_91_6;

Selector_2 s91_6(wires_22_5[3], addr_22_5, addr_positional[367:364], addr_91_6);

wire[27:0] addr_92_6;

Selector_2 s92_6(wires_23_5[0], addr_23_5, addr_positional[371:368], addr_92_6);

wire[27:0] addr_93_6;

Selector_2 s93_6(wires_23_5[1], addr_23_5, addr_positional[375:372], addr_93_6);

wire[27:0] addr_94_6;

Selector_2 s94_6(wires_23_5[2], addr_23_5, addr_positional[379:376], addr_94_6);

wire[27:0] addr_95_6;

Selector_2 s95_6(wires_23_5[3], addr_23_5, addr_positional[383:380], addr_95_6);

wire[27:0] addr_96_6;

Selector_2 s96_6(wires_24_5[0], addr_24_5, addr_positional[387:384], addr_96_6);

wire[27:0] addr_97_6;

Selector_2 s97_6(wires_24_5[1], addr_24_5, addr_positional[391:388], addr_97_6);

wire[27:0] addr_98_6;

Selector_2 s98_6(wires_24_5[2], addr_24_5, addr_positional[395:392], addr_98_6);

wire[27:0] addr_99_6;

Selector_2 s99_6(wires_24_5[3], addr_24_5, addr_positional[399:396], addr_99_6);

wire[27:0] addr_100_6;

Selector_2 s100_6(wires_25_5[0], addr_25_5, addr_positional[403:400], addr_100_6);

wire[27:0] addr_101_6;

Selector_2 s101_6(wires_25_5[1], addr_25_5, addr_positional[407:404], addr_101_6);

wire[27:0] addr_102_6;

Selector_2 s102_6(wires_25_5[2], addr_25_5, addr_positional[411:408], addr_102_6);

wire[27:0] addr_103_6;

Selector_2 s103_6(wires_25_5[3], addr_25_5, addr_positional[415:412], addr_103_6);

wire[27:0] addr_104_6;

Selector_2 s104_6(wires_26_5[0], addr_26_5, addr_positional[419:416], addr_104_6);

wire[27:0] addr_105_6;

Selector_2 s105_6(wires_26_5[1], addr_26_5, addr_positional[423:420], addr_105_6);

wire[27:0] addr_106_6;

Selector_2 s106_6(wires_26_5[2], addr_26_5, addr_positional[427:424], addr_106_6);

wire[27:0] addr_107_6;

Selector_2 s107_6(wires_26_5[3], addr_26_5, addr_positional[431:428], addr_107_6);

wire[27:0] addr_108_6;

Selector_2 s108_6(wires_27_5[0], addr_27_5, addr_positional[435:432], addr_108_6);

wire[27:0] addr_109_6;

Selector_2 s109_6(wires_27_5[1], addr_27_5, addr_positional[439:436], addr_109_6);

wire[27:0] addr_110_6;

Selector_2 s110_6(wires_27_5[2], addr_27_5, addr_positional[443:440], addr_110_6);

wire[27:0] addr_111_6;

Selector_2 s111_6(wires_27_5[3], addr_27_5, addr_positional[447:444], addr_111_6);

wire[27:0] addr_112_6;

Selector_2 s112_6(wires_28_5[0], addr_28_5, addr_positional[451:448], addr_112_6);

wire[27:0] addr_113_6;

Selector_2 s113_6(wires_28_5[1], addr_28_5, addr_positional[455:452], addr_113_6);

wire[27:0] addr_114_6;

Selector_2 s114_6(wires_28_5[2], addr_28_5, addr_positional[459:456], addr_114_6);

wire[27:0] addr_115_6;

Selector_2 s115_6(wires_28_5[3], addr_28_5, addr_positional[463:460], addr_115_6);

wire[27:0] addr_116_6;

Selector_2 s116_6(wires_29_5[0], addr_29_5, addr_positional[467:464], addr_116_6);

wire[27:0] addr_117_6;

Selector_2 s117_6(wires_29_5[1], addr_29_5, addr_positional[471:468], addr_117_6);

wire[27:0] addr_118_6;

Selector_2 s118_6(wires_29_5[2], addr_29_5, addr_positional[475:472], addr_118_6);

wire[27:0] addr_119_6;

Selector_2 s119_6(wires_29_5[3], addr_29_5, addr_positional[479:476], addr_119_6);

wire[27:0] addr_120_6;

Selector_2 s120_6(wires_30_5[0], addr_30_5, addr_positional[483:480], addr_120_6);

wire[27:0] addr_121_6;

Selector_2 s121_6(wires_30_5[1], addr_30_5, addr_positional[487:484], addr_121_6);

wire[27:0] addr_122_6;

Selector_2 s122_6(wires_30_5[2], addr_30_5, addr_positional[491:488], addr_122_6);

wire[27:0] addr_123_6;

Selector_2 s123_6(wires_30_5[3], addr_30_5, addr_positional[495:492], addr_123_6);

wire[27:0] addr_124_6;

Selector_2 s124_6(wires_31_5[0], addr_31_5, addr_positional[499:496], addr_124_6);

wire[27:0] addr_125_6;

Selector_2 s125_6(wires_31_5[1], addr_31_5, addr_positional[503:500], addr_125_6);

wire[27:0] addr_126_6;

Selector_2 s126_6(wires_31_5[2], addr_31_5, addr_positional[507:504], addr_126_6);

wire[27:0] addr_127_6;

Selector_2 s127_6(wires_31_5[3], addr_31_5, addr_positional[511:508], addr_127_6);

wire[27:0] addr_128_6;

Selector_2 s128_6(wires_32_5[0], addr_32_5, addr_positional[515:512], addr_128_6);

wire[27:0] addr_129_6;

Selector_2 s129_6(wires_32_5[1], addr_32_5, addr_positional[519:516], addr_129_6);

wire[27:0] addr_130_6;

Selector_2 s130_6(wires_32_5[2], addr_32_5, addr_positional[523:520], addr_130_6);

wire[27:0] addr_131_6;

Selector_2 s131_6(wires_32_5[3], addr_32_5, addr_positional[527:524], addr_131_6);

wire[27:0] addr_132_6;

Selector_2 s132_6(wires_33_5[0], addr_33_5, addr_positional[531:528], addr_132_6);

wire[27:0] addr_133_6;

Selector_2 s133_6(wires_33_5[1], addr_33_5, addr_positional[535:532], addr_133_6);

wire[27:0] addr_134_6;

Selector_2 s134_6(wires_33_5[2], addr_33_5, addr_positional[539:536], addr_134_6);

wire[27:0] addr_135_6;

Selector_2 s135_6(wires_33_5[3], addr_33_5, addr_positional[543:540], addr_135_6);

wire[27:0] addr_136_6;

Selector_2 s136_6(wires_34_5[0], addr_34_5, addr_positional[547:544], addr_136_6);

wire[27:0] addr_137_6;

Selector_2 s137_6(wires_34_5[1], addr_34_5, addr_positional[551:548], addr_137_6);

wire[27:0] addr_138_6;

Selector_2 s138_6(wires_34_5[2], addr_34_5, addr_positional[555:552], addr_138_6);

wire[27:0] addr_139_6;

Selector_2 s139_6(wires_34_5[3], addr_34_5, addr_positional[559:556], addr_139_6);

wire[27:0] addr_140_6;

Selector_2 s140_6(wires_35_5[0], addr_35_5, addr_positional[563:560], addr_140_6);

wire[27:0] addr_141_6;

Selector_2 s141_6(wires_35_5[1], addr_35_5, addr_positional[567:564], addr_141_6);

wire[27:0] addr_142_6;

Selector_2 s142_6(wires_35_5[2], addr_35_5, addr_positional[571:568], addr_142_6);

wire[27:0] addr_143_6;

Selector_2 s143_6(wires_35_5[3], addr_35_5, addr_positional[575:572], addr_143_6);

wire[27:0] addr_144_6;

Selector_2 s144_6(wires_36_5[0], addr_36_5, addr_positional[579:576], addr_144_6);

wire[27:0] addr_145_6;

Selector_2 s145_6(wires_36_5[1], addr_36_5, addr_positional[583:580], addr_145_6);

wire[27:0] addr_146_6;

Selector_2 s146_6(wires_36_5[2], addr_36_5, addr_positional[587:584], addr_146_6);

wire[27:0] addr_147_6;

Selector_2 s147_6(wires_36_5[3], addr_36_5, addr_positional[591:588], addr_147_6);

wire[27:0] addr_148_6;

Selector_2 s148_6(wires_37_5[0], addr_37_5, addr_positional[595:592], addr_148_6);

wire[27:0] addr_149_6;

Selector_2 s149_6(wires_37_5[1], addr_37_5, addr_positional[599:596], addr_149_6);

wire[27:0] addr_150_6;

Selector_2 s150_6(wires_37_5[2], addr_37_5, addr_positional[603:600], addr_150_6);

wire[27:0] addr_151_6;

Selector_2 s151_6(wires_37_5[3], addr_37_5, addr_positional[607:604], addr_151_6);

wire[27:0] addr_152_6;

Selector_2 s152_6(wires_38_5[0], addr_38_5, addr_positional[611:608], addr_152_6);

wire[27:0] addr_153_6;

Selector_2 s153_6(wires_38_5[1], addr_38_5, addr_positional[615:612], addr_153_6);

wire[27:0] addr_154_6;

Selector_2 s154_6(wires_38_5[2], addr_38_5, addr_positional[619:616], addr_154_6);

wire[27:0] addr_155_6;

Selector_2 s155_6(wires_38_5[3], addr_38_5, addr_positional[623:620], addr_155_6);

wire[27:0] addr_156_6;

Selector_2 s156_6(wires_39_5[0], addr_39_5, addr_positional[627:624], addr_156_6);

wire[27:0] addr_157_6;

Selector_2 s157_6(wires_39_5[1], addr_39_5, addr_positional[631:628], addr_157_6);

wire[27:0] addr_158_6;

Selector_2 s158_6(wires_39_5[2], addr_39_5, addr_positional[635:632], addr_158_6);

wire[27:0] addr_159_6;

Selector_2 s159_6(wires_39_5[3], addr_39_5, addr_positional[639:636], addr_159_6);

wire[27:0] addr_160_6;

Selector_2 s160_6(wires_40_5[0], addr_40_5, addr_positional[643:640], addr_160_6);

wire[27:0] addr_161_6;

Selector_2 s161_6(wires_40_5[1], addr_40_5, addr_positional[647:644], addr_161_6);

wire[27:0] addr_162_6;

Selector_2 s162_6(wires_40_5[2], addr_40_5, addr_positional[651:648], addr_162_6);

wire[27:0] addr_163_6;

Selector_2 s163_6(wires_40_5[3], addr_40_5, addr_positional[655:652], addr_163_6);

wire[27:0] addr_164_6;

Selector_2 s164_6(wires_41_5[0], addr_41_5, addr_positional[659:656], addr_164_6);

wire[27:0] addr_165_6;

Selector_2 s165_6(wires_41_5[1], addr_41_5, addr_positional[663:660], addr_165_6);

wire[27:0] addr_166_6;

Selector_2 s166_6(wires_41_5[2], addr_41_5, addr_positional[667:664], addr_166_6);

wire[27:0] addr_167_6;

Selector_2 s167_6(wires_41_5[3], addr_41_5, addr_positional[671:668], addr_167_6);

wire[27:0] addr_168_6;

Selector_2 s168_6(wires_42_5[0], addr_42_5, addr_positional[675:672], addr_168_6);

wire[27:0] addr_169_6;

Selector_2 s169_6(wires_42_5[1], addr_42_5, addr_positional[679:676], addr_169_6);

wire[27:0] addr_170_6;

Selector_2 s170_6(wires_42_5[2], addr_42_5, addr_positional[683:680], addr_170_6);

wire[27:0] addr_171_6;

Selector_2 s171_6(wires_42_5[3], addr_42_5, addr_positional[687:684], addr_171_6);

wire[27:0] addr_172_6;

Selector_2 s172_6(wires_43_5[0], addr_43_5, addr_positional[691:688], addr_172_6);

wire[27:0] addr_173_6;

Selector_2 s173_6(wires_43_5[1], addr_43_5, addr_positional[695:692], addr_173_6);

wire[27:0] addr_174_6;

Selector_2 s174_6(wires_43_5[2], addr_43_5, addr_positional[699:696], addr_174_6);

wire[27:0] addr_175_6;

Selector_2 s175_6(wires_43_5[3], addr_43_5, addr_positional[703:700], addr_175_6);

wire[27:0] addr_176_6;

Selector_2 s176_6(wires_44_5[0], addr_44_5, addr_positional[707:704], addr_176_6);

wire[27:0] addr_177_6;

Selector_2 s177_6(wires_44_5[1], addr_44_5, addr_positional[711:708], addr_177_6);

wire[27:0] addr_178_6;

Selector_2 s178_6(wires_44_5[2], addr_44_5, addr_positional[715:712], addr_178_6);

wire[27:0] addr_179_6;

Selector_2 s179_6(wires_44_5[3], addr_44_5, addr_positional[719:716], addr_179_6);

wire[27:0] addr_180_6;

Selector_2 s180_6(wires_45_5[0], addr_45_5, addr_positional[723:720], addr_180_6);

wire[27:0] addr_181_6;

Selector_2 s181_6(wires_45_5[1], addr_45_5, addr_positional[727:724], addr_181_6);

wire[27:0] addr_182_6;

Selector_2 s182_6(wires_45_5[2], addr_45_5, addr_positional[731:728], addr_182_6);

wire[27:0] addr_183_6;

Selector_2 s183_6(wires_45_5[3], addr_45_5, addr_positional[735:732], addr_183_6);

wire[27:0] addr_184_6;

Selector_2 s184_6(wires_46_5[0], addr_46_5, addr_positional[739:736], addr_184_6);

wire[27:0] addr_185_6;

Selector_2 s185_6(wires_46_5[1], addr_46_5, addr_positional[743:740], addr_185_6);

wire[27:0] addr_186_6;

Selector_2 s186_6(wires_46_5[2], addr_46_5, addr_positional[747:744], addr_186_6);

wire[27:0] addr_187_6;

Selector_2 s187_6(wires_46_5[3], addr_46_5, addr_positional[751:748], addr_187_6);

wire[27:0] addr_188_6;

Selector_2 s188_6(wires_47_5[0], addr_47_5, addr_positional[755:752], addr_188_6);

wire[27:0] addr_189_6;

Selector_2 s189_6(wires_47_5[1], addr_47_5, addr_positional[759:756], addr_189_6);

wire[27:0] addr_190_6;

Selector_2 s190_6(wires_47_5[2], addr_47_5, addr_positional[763:760], addr_190_6);

wire[27:0] addr_191_6;

Selector_2 s191_6(wires_47_5[3], addr_47_5, addr_positional[767:764], addr_191_6);

wire[27:0] addr_192_6;

Selector_2 s192_6(wires_48_5[0], addr_48_5, addr_positional[771:768], addr_192_6);

wire[27:0] addr_193_6;

Selector_2 s193_6(wires_48_5[1], addr_48_5, addr_positional[775:772], addr_193_6);

wire[27:0] addr_194_6;

Selector_2 s194_6(wires_48_5[2], addr_48_5, addr_positional[779:776], addr_194_6);

wire[27:0] addr_195_6;

Selector_2 s195_6(wires_48_5[3], addr_48_5, addr_positional[783:780], addr_195_6);

wire[27:0] addr_196_6;

Selector_2 s196_6(wires_49_5[0], addr_49_5, addr_positional[787:784], addr_196_6);

wire[27:0] addr_197_6;

Selector_2 s197_6(wires_49_5[1], addr_49_5, addr_positional[791:788], addr_197_6);

wire[27:0] addr_198_6;

Selector_2 s198_6(wires_49_5[2], addr_49_5, addr_positional[795:792], addr_198_6);

wire[27:0] addr_199_6;

Selector_2 s199_6(wires_49_5[3], addr_49_5, addr_positional[799:796], addr_199_6);

wire[27:0] addr_200_6;

Selector_2 s200_6(wires_50_5[0], addr_50_5, addr_positional[803:800], addr_200_6);

wire[27:0] addr_201_6;

Selector_2 s201_6(wires_50_5[1], addr_50_5, addr_positional[807:804], addr_201_6);

wire[27:0] addr_202_6;

Selector_2 s202_6(wires_50_5[2], addr_50_5, addr_positional[811:808], addr_202_6);

wire[27:0] addr_203_6;

Selector_2 s203_6(wires_50_5[3], addr_50_5, addr_positional[815:812], addr_203_6);

wire[27:0] addr_204_6;

Selector_2 s204_6(wires_51_5[0], addr_51_5, addr_positional[819:816], addr_204_6);

wire[27:0] addr_205_6;

Selector_2 s205_6(wires_51_5[1], addr_51_5, addr_positional[823:820], addr_205_6);

wire[27:0] addr_206_6;

Selector_2 s206_6(wires_51_5[2], addr_51_5, addr_positional[827:824], addr_206_6);

wire[27:0] addr_207_6;

Selector_2 s207_6(wires_51_5[3], addr_51_5, addr_positional[831:828], addr_207_6);

wire[27:0] addr_208_6;

Selector_2 s208_6(wires_52_5[0], addr_52_5, addr_positional[835:832], addr_208_6);

wire[27:0] addr_209_6;

Selector_2 s209_6(wires_52_5[1], addr_52_5, addr_positional[839:836], addr_209_6);

wire[27:0] addr_210_6;

Selector_2 s210_6(wires_52_5[2], addr_52_5, addr_positional[843:840], addr_210_6);

wire[27:0] addr_211_6;

Selector_2 s211_6(wires_52_5[3], addr_52_5, addr_positional[847:844], addr_211_6);

wire[27:0] addr_212_6;

Selector_2 s212_6(wires_53_5[0], addr_53_5, addr_positional[851:848], addr_212_6);

wire[27:0] addr_213_6;

Selector_2 s213_6(wires_53_5[1], addr_53_5, addr_positional[855:852], addr_213_6);

wire[27:0] addr_214_6;

Selector_2 s214_6(wires_53_5[2], addr_53_5, addr_positional[859:856], addr_214_6);

wire[27:0] addr_215_6;

Selector_2 s215_6(wires_53_5[3], addr_53_5, addr_positional[863:860], addr_215_6);

wire[27:0] addr_216_6;

Selector_2 s216_6(wires_54_5[0], addr_54_5, addr_positional[867:864], addr_216_6);

wire[27:0] addr_217_6;

Selector_2 s217_6(wires_54_5[1], addr_54_5, addr_positional[871:868], addr_217_6);

wire[27:0] addr_218_6;

Selector_2 s218_6(wires_54_5[2], addr_54_5, addr_positional[875:872], addr_218_6);

wire[27:0] addr_219_6;

Selector_2 s219_6(wires_54_5[3], addr_54_5, addr_positional[879:876], addr_219_6);

wire[27:0] addr_220_6;

Selector_2 s220_6(wires_55_5[0], addr_55_5, addr_positional[883:880], addr_220_6);

wire[27:0] addr_221_6;

Selector_2 s221_6(wires_55_5[1], addr_55_5, addr_positional[887:884], addr_221_6);

wire[27:0] addr_222_6;

Selector_2 s222_6(wires_55_5[2], addr_55_5, addr_positional[891:888], addr_222_6);

wire[27:0] addr_223_6;

Selector_2 s223_6(wires_55_5[3], addr_55_5, addr_positional[895:892], addr_223_6);

wire[27:0] addr_224_6;

Selector_2 s224_6(wires_56_5[0], addr_56_5, addr_positional[899:896], addr_224_6);

wire[27:0] addr_225_6;

Selector_2 s225_6(wires_56_5[1], addr_56_5, addr_positional[903:900], addr_225_6);

wire[27:0] addr_226_6;

Selector_2 s226_6(wires_56_5[2], addr_56_5, addr_positional[907:904], addr_226_6);

wire[27:0] addr_227_6;

Selector_2 s227_6(wires_56_5[3], addr_56_5, addr_positional[911:908], addr_227_6);

wire[27:0] addr_228_6;

Selector_2 s228_6(wires_57_5[0], addr_57_5, addr_positional[915:912], addr_228_6);

wire[27:0] addr_229_6;

Selector_2 s229_6(wires_57_5[1], addr_57_5, addr_positional[919:916], addr_229_6);

wire[27:0] addr_230_6;

Selector_2 s230_6(wires_57_5[2], addr_57_5, addr_positional[923:920], addr_230_6);

wire[27:0] addr_231_6;

Selector_2 s231_6(wires_57_5[3], addr_57_5, addr_positional[927:924], addr_231_6);

wire[27:0] addr_232_6;

Selector_2 s232_6(wires_58_5[0], addr_58_5, addr_positional[931:928], addr_232_6);

wire[27:0] addr_233_6;

Selector_2 s233_6(wires_58_5[1], addr_58_5, addr_positional[935:932], addr_233_6);

wire[27:0] addr_234_6;

Selector_2 s234_6(wires_58_5[2], addr_58_5, addr_positional[939:936], addr_234_6);

wire[27:0] addr_235_6;

Selector_2 s235_6(wires_58_5[3], addr_58_5, addr_positional[943:940], addr_235_6);

wire[27:0] addr_236_6;

Selector_2 s236_6(wires_59_5[0], addr_59_5, addr_positional[947:944], addr_236_6);

wire[27:0] addr_237_6;

Selector_2 s237_6(wires_59_5[1], addr_59_5, addr_positional[951:948], addr_237_6);

wire[27:0] addr_238_6;

Selector_2 s238_6(wires_59_5[2], addr_59_5, addr_positional[955:952], addr_238_6);

wire[27:0] addr_239_6;

Selector_2 s239_6(wires_59_5[3], addr_59_5, addr_positional[959:956], addr_239_6);

wire[27:0] addr_240_6;

Selector_2 s240_6(wires_60_5[0], addr_60_5, addr_positional[963:960], addr_240_6);

wire[27:0] addr_241_6;

Selector_2 s241_6(wires_60_5[1], addr_60_5, addr_positional[967:964], addr_241_6);

wire[27:0] addr_242_6;

Selector_2 s242_6(wires_60_5[2], addr_60_5, addr_positional[971:968], addr_242_6);

wire[27:0] addr_243_6;

Selector_2 s243_6(wires_60_5[3], addr_60_5, addr_positional[975:972], addr_243_6);

wire[27:0] addr_244_6;

Selector_2 s244_6(wires_61_5[0], addr_61_5, addr_positional[979:976], addr_244_6);

wire[27:0] addr_245_6;

Selector_2 s245_6(wires_61_5[1], addr_61_5, addr_positional[983:980], addr_245_6);

wire[27:0] addr_246_6;

Selector_2 s246_6(wires_61_5[2], addr_61_5, addr_positional[987:984], addr_246_6);

wire[27:0] addr_247_6;

Selector_2 s247_6(wires_61_5[3], addr_61_5, addr_positional[991:988], addr_247_6);

wire[27:0] addr_248_6;

Selector_2 s248_6(wires_62_5[0], addr_62_5, addr_positional[995:992], addr_248_6);

wire[27:0] addr_249_6;

Selector_2 s249_6(wires_62_5[1], addr_62_5, addr_positional[999:996], addr_249_6);

wire[27:0] addr_250_6;

Selector_2 s250_6(wires_62_5[2], addr_62_5, addr_positional[1003:1000], addr_250_6);

wire[27:0] addr_251_6;

Selector_2 s251_6(wires_62_5[3], addr_62_5, addr_positional[1007:1004], addr_251_6);

wire[27:0] addr_252_6;

Selector_2 s252_6(wires_63_5[0], addr_63_5, addr_positional[1011:1008], addr_252_6);

wire[27:0] addr_253_6;

Selector_2 s253_6(wires_63_5[1], addr_63_5, addr_positional[1015:1012], addr_253_6);

wire[27:0] addr_254_6;

Selector_2 s254_6(wires_63_5[2], addr_63_5, addr_positional[1019:1016], addr_254_6);

wire[27:0] addr_255_6;

Selector_2 s255_6(wires_63_5[3], addr_63_5, addr_positional[1023:1020], addr_255_6);

wire[27:0] addr_256_6;

Selector_2 s256_6(wires_64_5[0], addr_64_5, addr_positional[1027:1024], addr_256_6);

wire[27:0] addr_257_6;

Selector_2 s257_6(wires_64_5[1], addr_64_5, addr_positional[1031:1028], addr_257_6);

wire[27:0] addr_258_6;

Selector_2 s258_6(wires_64_5[2], addr_64_5, addr_positional[1035:1032], addr_258_6);

wire[27:0] addr_259_6;

Selector_2 s259_6(wires_64_5[3], addr_64_5, addr_positional[1039:1036], addr_259_6);

wire[27:0] addr_260_6;

Selector_2 s260_6(wires_65_5[0], addr_65_5, addr_positional[1043:1040], addr_260_6);

wire[27:0] addr_261_6;

Selector_2 s261_6(wires_65_5[1], addr_65_5, addr_positional[1047:1044], addr_261_6);

wire[27:0] addr_262_6;

Selector_2 s262_6(wires_65_5[2], addr_65_5, addr_positional[1051:1048], addr_262_6);

wire[27:0] addr_263_6;

Selector_2 s263_6(wires_65_5[3], addr_65_5, addr_positional[1055:1052], addr_263_6);

wire[27:0] addr_264_6;

Selector_2 s264_6(wires_66_5[0], addr_66_5, addr_positional[1059:1056], addr_264_6);

wire[27:0] addr_265_6;

Selector_2 s265_6(wires_66_5[1], addr_66_5, addr_positional[1063:1060], addr_265_6);

wire[27:0] addr_266_6;

Selector_2 s266_6(wires_66_5[2], addr_66_5, addr_positional[1067:1064], addr_266_6);

wire[27:0] addr_267_6;

Selector_2 s267_6(wires_66_5[3], addr_66_5, addr_positional[1071:1068], addr_267_6);

wire[27:0] addr_268_6;

Selector_2 s268_6(wires_67_5[0], addr_67_5, addr_positional[1075:1072], addr_268_6);

wire[27:0] addr_269_6;

Selector_2 s269_6(wires_67_5[1], addr_67_5, addr_positional[1079:1076], addr_269_6);

wire[27:0] addr_270_6;

Selector_2 s270_6(wires_67_5[2], addr_67_5, addr_positional[1083:1080], addr_270_6);

wire[27:0] addr_271_6;

Selector_2 s271_6(wires_67_5[3], addr_67_5, addr_positional[1087:1084], addr_271_6);

wire[27:0] addr_272_6;

Selector_2 s272_6(wires_68_5[0], addr_68_5, addr_positional[1091:1088], addr_272_6);

wire[27:0] addr_273_6;

Selector_2 s273_6(wires_68_5[1], addr_68_5, addr_positional[1095:1092], addr_273_6);

wire[27:0] addr_274_6;

Selector_2 s274_6(wires_68_5[2], addr_68_5, addr_positional[1099:1096], addr_274_6);

wire[27:0] addr_275_6;

Selector_2 s275_6(wires_68_5[3], addr_68_5, addr_positional[1103:1100], addr_275_6);

wire[27:0] addr_276_6;

Selector_2 s276_6(wires_69_5[0], addr_69_5, addr_positional[1107:1104], addr_276_6);

wire[27:0] addr_277_6;

Selector_2 s277_6(wires_69_5[1], addr_69_5, addr_positional[1111:1108], addr_277_6);

wire[27:0] addr_278_6;

Selector_2 s278_6(wires_69_5[2], addr_69_5, addr_positional[1115:1112], addr_278_6);

wire[27:0] addr_279_6;

Selector_2 s279_6(wires_69_5[3], addr_69_5, addr_positional[1119:1116], addr_279_6);

wire[27:0] addr_280_6;

Selector_2 s280_6(wires_70_5[0], addr_70_5, addr_positional[1123:1120], addr_280_6);

wire[27:0] addr_281_6;

Selector_2 s281_6(wires_70_5[1], addr_70_5, addr_positional[1127:1124], addr_281_6);

wire[27:0] addr_282_6;

Selector_2 s282_6(wires_70_5[2], addr_70_5, addr_positional[1131:1128], addr_282_6);

wire[27:0] addr_283_6;

Selector_2 s283_6(wires_70_5[3], addr_70_5, addr_positional[1135:1132], addr_283_6);

wire[27:0] addr_284_6;

Selector_2 s284_6(wires_71_5[0], addr_71_5, addr_positional[1139:1136], addr_284_6);

wire[27:0] addr_285_6;

Selector_2 s285_6(wires_71_5[1], addr_71_5, addr_positional[1143:1140], addr_285_6);

wire[27:0] addr_286_6;

Selector_2 s286_6(wires_71_5[2], addr_71_5, addr_positional[1147:1144], addr_286_6);

wire[27:0] addr_287_6;

Selector_2 s287_6(wires_71_5[3], addr_71_5, addr_positional[1151:1148], addr_287_6);

wire[27:0] addr_288_6;

Selector_2 s288_6(wires_72_5[0], addr_72_5, addr_positional[1155:1152], addr_288_6);

wire[27:0] addr_289_6;

Selector_2 s289_6(wires_72_5[1], addr_72_5, addr_positional[1159:1156], addr_289_6);

wire[27:0] addr_290_6;

Selector_2 s290_6(wires_72_5[2], addr_72_5, addr_positional[1163:1160], addr_290_6);

wire[27:0] addr_291_6;

Selector_2 s291_6(wires_72_5[3], addr_72_5, addr_positional[1167:1164], addr_291_6);

wire[27:0] addr_292_6;

Selector_2 s292_6(wires_73_5[0], addr_73_5, addr_positional[1171:1168], addr_292_6);

wire[27:0] addr_293_6;

Selector_2 s293_6(wires_73_5[1], addr_73_5, addr_positional[1175:1172], addr_293_6);

wire[27:0] addr_294_6;

Selector_2 s294_6(wires_73_5[2], addr_73_5, addr_positional[1179:1176], addr_294_6);

wire[27:0] addr_295_6;

Selector_2 s295_6(wires_73_5[3], addr_73_5, addr_positional[1183:1180], addr_295_6);

wire[27:0] addr_296_6;

Selector_2 s296_6(wires_74_5[0], addr_74_5, addr_positional[1187:1184], addr_296_6);

wire[27:0] addr_297_6;

Selector_2 s297_6(wires_74_5[1], addr_74_5, addr_positional[1191:1188], addr_297_6);

wire[27:0] addr_298_6;

Selector_2 s298_6(wires_74_5[2], addr_74_5, addr_positional[1195:1192], addr_298_6);

wire[27:0] addr_299_6;

Selector_2 s299_6(wires_74_5[3], addr_74_5, addr_positional[1199:1196], addr_299_6);

wire[27:0] addr_300_6;

Selector_2 s300_6(wires_75_5[0], addr_75_5, addr_positional[1203:1200], addr_300_6);

wire[27:0] addr_301_6;

Selector_2 s301_6(wires_75_5[1], addr_75_5, addr_positional[1207:1204], addr_301_6);

wire[27:0] addr_302_6;

Selector_2 s302_6(wires_75_5[2], addr_75_5, addr_positional[1211:1208], addr_302_6);

wire[27:0] addr_303_6;

Selector_2 s303_6(wires_75_5[3], addr_75_5, addr_positional[1215:1212], addr_303_6);

wire[27:0] addr_304_6;

Selector_2 s304_6(wires_76_5[0], addr_76_5, addr_positional[1219:1216], addr_304_6);

wire[27:0] addr_305_6;

Selector_2 s305_6(wires_76_5[1], addr_76_5, addr_positional[1223:1220], addr_305_6);

wire[27:0] addr_306_6;

Selector_2 s306_6(wires_76_5[2], addr_76_5, addr_positional[1227:1224], addr_306_6);

wire[27:0] addr_307_6;

Selector_2 s307_6(wires_76_5[3], addr_76_5, addr_positional[1231:1228], addr_307_6);

wire[27:0] addr_308_6;

Selector_2 s308_6(wires_77_5[0], addr_77_5, addr_positional[1235:1232], addr_308_6);

wire[27:0] addr_309_6;

Selector_2 s309_6(wires_77_5[1], addr_77_5, addr_positional[1239:1236], addr_309_6);

wire[27:0] addr_310_6;

Selector_2 s310_6(wires_77_5[2], addr_77_5, addr_positional[1243:1240], addr_310_6);

wire[27:0] addr_311_6;

Selector_2 s311_6(wires_77_5[3], addr_77_5, addr_positional[1247:1244], addr_311_6);

wire[27:0] addr_312_6;

Selector_2 s312_6(wires_78_5[0], addr_78_5, addr_positional[1251:1248], addr_312_6);

wire[27:0] addr_313_6;

Selector_2 s313_6(wires_78_5[1], addr_78_5, addr_positional[1255:1252], addr_313_6);

wire[27:0] addr_314_6;

Selector_2 s314_6(wires_78_5[2], addr_78_5, addr_positional[1259:1256], addr_314_6);

wire[27:0] addr_315_6;

Selector_2 s315_6(wires_78_5[3], addr_78_5, addr_positional[1263:1260], addr_315_6);

wire[27:0] addr_316_6;

Selector_2 s316_6(wires_79_5[0], addr_79_5, addr_positional[1267:1264], addr_316_6);

wire[27:0] addr_317_6;

Selector_2 s317_6(wires_79_5[1], addr_79_5, addr_positional[1271:1268], addr_317_6);

wire[27:0] addr_318_6;

Selector_2 s318_6(wires_79_5[2], addr_79_5, addr_positional[1275:1272], addr_318_6);

wire[27:0] addr_319_6;

Selector_2 s319_6(wires_79_5[3], addr_79_5, addr_positional[1279:1276], addr_319_6);

wire[27:0] addr_320_6;

Selector_2 s320_6(wires_80_5[0], addr_80_5, addr_positional[1283:1280], addr_320_6);

wire[27:0] addr_321_6;

Selector_2 s321_6(wires_80_5[1], addr_80_5, addr_positional[1287:1284], addr_321_6);

wire[27:0] addr_322_6;

Selector_2 s322_6(wires_80_5[2], addr_80_5, addr_positional[1291:1288], addr_322_6);

wire[27:0] addr_323_6;

Selector_2 s323_6(wires_80_5[3], addr_80_5, addr_positional[1295:1292], addr_323_6);

wire[27:0] addr_324_6;

Selector_2 s324_6(wires_81_5[0], addr_81_5, addr_positional[1299:1296], addr_324_6);

wire[27:0] addr_325_6;

Selector_2 s325_6(wires_81_5[1], addr_81_5, addr_positional[1303:1300], addr_325_6);

wire[27:0] addr_326_6;

Selector_2 s326_6(wires_81_5[2], addr_81_5, addr_positional[1307:1304], addr_326_6);

wire[27:0] addr_327_6;

Selector_2 s327_6(wires_81_5[3], addr_81_5, addr_positional[1311:1308], addr_327_6);

wire[27:0] addr_328_6;

Selector_2 s328_6(wires_82_5[0], addr_82_5, addr_positional[1315:1312], addr_328_6);

wire[27:0] addr_329_6;

Selector_2 s329_6(wires_82_5[1], addr_82_5, addr_positional[1319:1316], addr_329_6);

wire[27:0] addr_330_6;

Selector_2 s330_6(wires_82_5[2], addr_82_5, addr_positional[1323:1320], addr_330_6);

wire[27:0] addr_331_6;

Selector_2 s331_6(wires_82_5[3], addr_82_5, addr_positional[1327:1324], addr_331_6);

wire[27:0] addr_332_6;

Selector_2 s332_6(wires_83_5[0], addr_83_5, addr_positional[1331:1328], addr_332_6);

wire[27:0] addr_333_6;

Selector_2 s333_6(wires_83_5[1], addr_83_5, addr_positional[1335:1332], addr_333_6);

wire[27:0] addr_334_6;

Selector_2 s334_6(wires_83_5[2], addr_83_5, addr_positional[1339:1336], addr_334_6);

wire[27:0] addr_335_6;

Selector_2 s335_6(wires_83_5[3], addr_83_5, addr_positional[1343:1340], addr_335_6);

wire[27:0] addr_336_6;

Selector_2 s336_6(wires_84_5[0], addr_84_5, addr_positional[1347:1344], addr_336_6);

wire[27:0] addr_337_6;

Selector_2 s337_6(wires_84_5[1], addr_84_5, addr_positional[1351:1348], addr_337_6);

wire[27:0] addr_338_6;

Selector_2 s338_6(wires_84_5[2], addr_84_5, addr_positional[1355:1352], addr_338_6);

wire[27:0] addr_339_6;

Selector_2 s339_6(wires_84_5[3], addr_84_5, addr_positional[1359:1356], addr_339_6);

wire[27:0] addr_340_6;

Selector_2 s340_6(wires_85_5[0], addr_85_5, addr_positional[1363:1360], addr_340_6);

wire[27:0] addr_341_6;

Selector_2 s341_6(wires_85_5[1], addr_85_5, addr_positional[1367:1364], addr_341_6);

wire[27:0] addr_342_6;

Selector_2 s342_6(wires_85_5[2], addr_85_5, addr_positional[1371:1368], addr_342_6);

wire[27:0] addr_343_6;

Selector_2 s343_6(wires_85_5[3], addr_85_5, addr_positional[1375:1372], addr_343_6);

wire[27:0] addr_344_6;

Selector_2 s344_6(wires_86_5[0], addr_86_5, addr_positional[1379:1376], addr_344_6);

wire[27:0] addr_345_6;

Selector_2 s345_6(wires_86_5[1], addr_86_5, addr_positional[1383:1380], addr_345_6);

wire[27:0] addr_346_6;

Selector_2 s346_6(wires_86_5[2], addr_86_5, addr_positional[1387:1384], addr_346_6);

wire[27:0] addr_347_6;

Selector_2 s347_6(wires_86_5[3], addr_86_5, addr_positional[1391:1388], addr_347_6);

wire[27:0] addr_348_6;

Selector_2 s348_6(wires_87_5[0], addr_87_5, addr_positional[1395:1392], addr_348_6);

wire[27:0] addr_349_6;

Selector_2 s349_6(wires_87_5[1], addr_87_5, addr_positional[1399:1396], addr_349_6);

wire[27:0] addr_350_6;

Selector_2 s350_6(wires_87_5[2], addr_87_5, addr_positional[1403:1400], addr_350_6);

wire[27:0] addr_351_6;

Selector_2 s351_6(wires_87_5[3], addr_87_5, addr_positional[1407:1404], addr_351_6);

wire[27:0] addr_352_6;

Selector_2 s352_6(wires_88_5[0], addr_88_5, addr_positional[1411:1408], addr_352_6);

wire[27:0] addr_353_6;

Selector_2 s353_6(wires_88_5[1], addr_88_5, addr_positional[1415:1412], addr_353_6);

wire[27:0] addr_354_6;

Selector_2 s354_6(wires_88_5[2], addr_88_5, addr_positional[1419:1416], addr_354_6);

wire[27:0] addr_355_6;

Selector_2 s355_6(wires_88_5[3], addr_88_5, addr_positional[1423:1420], addr_355_6);

wire[27:0] addr_356_6;

Selector_2 s356_6(wires_89_5[0], addr_89_5, addr_positional[1427:1424], addr_356_6);

wire[27:0] addr_357_6;

Selector_2 s357_6(wires_89_5[1], addr_89_5, addr_positional[1431:1428], addr_357_6);

wire[27:0] addr_358_6;

Selector_2 s358_6(wires_89_5[2], addr_89_5, addr_positional[1435:1432], addr_358_6);

wire[27:0] addr_359_6;

Selector_2 s359_6(wires_89_5[3], addr_89_5, addr_positional[1439:1436], addr_359_6);

wire[27:0] addr_360_6;

Selector_2 s360_6(wires_90_5[0], addr_90_5, addr_positional[1443:1440], addr_360_6);

wire[27:0] addr_361_6;

Selector_2 s361_6(wires_90_5[1], addr_90_5, addr_positional[1447:1444], addr_361_6);

wire[27:0] addr_362_6;

Selector_2 s362_6(wires_90_5[2], addr_90_5, addr_positional[1451:1448], addr_362_6);

wire[27:0] addr_363_6;

Selector_2 s363_6(wires_90_5[3], addr_90_5, addr_positional[1455:1452], addr_363_6);

wire[27:0] addr_364_6;

Selector_2 s364_6(wires_91_5[0], addr_91_5, addr_positional[1459:1456], addr_364_6);

wire[27:0] addr_365_6;

Selector_2 s365_6(wires_91_5[1], addr_91_5, addr_positional[1463:1460], addr_365_6);

wire[27:0] addr_366_6;

Selector_2 s366_6(wires_91_5[2], addr_91_5, addr_positional[1467:1464], addr_366_6);

wire[27:0] addr_367_6;

Selector_2 s367_6(wires_91_5[3], addr_91_5, addr_positional[1471:1468], addr_367_6);

wire[27:0] addr_368_6;

Selector_2 s368_6(wires_92_5[0], addr_92_5, addr_positional[1475:1472], addr_368_6);

wire[27:0] addr_369_6;

Selector_2 s369_6(wires_92_5[1], addr_92_5, addr_positional[1479:1476], addr_369_6);

wire[27:0] addr_370_6;

Selector_2 s370_6(wires_92_5[2], addr_92_5, addr_positional[1483:1480], addr_370_6);

wire[27:0] addr_371_6;

Selector_2 s371_6(wires_92_5[3], addr_92_5, addr_positional[1487:1484], addr_371_6);

wire[27:0] addr_372_6;

Selector_2 s372_6(wires_93_5[0], addr_93_5, addr_positional[1491:1488], addr_372_6);

wire[27:0] addr_373_6;

Selector_2 s373_6(wires_93_5[1], addr_93_5, addr_positional[1495:1492], addr_373_6);

wire[27:0] addr_374_6;

Selector_2 s374_6(wires_93_5[2], addr_93_5, addr_positional[1499:1496], addr_374_6);

wire[27:0] addr_375_6;

Selector_2 s375_6(wires_93_5[3], addr_93_5, addr_positional[1503:1500], addr_375_6);

wire[27:0] addr_376_6;

Selector_2 s376_6(wires_94_5[0], addr_94_5, addr_positional[1507:1504], addr_376_6);

wire[27:0] addr_377_6;

Selector_2 s377_6(wires_94_5[1], addr_94_5, addr_positional[1511:1508], addr_377_6);

wire[27:0] addr_378_6;

Selector_2 s378_6(wires_94_5[2], addr_94_5, addr_positional[1515:1512], addr_378_6);

wire[27:0] addr_379_6;

Selector_2 s379_6(wires_94_5[3], addr_94_5, addr_positional[1519:1516], addr_379_6);

wire[27:0] addr_380_6;

Selector_2 s380_6(wires_95_5[0], addr_95_5, addr_positional[1523:1520], addr_380_6);

wire[27:0] addr_381_6;

Selector_2 s381_6(wires_95_5[1], addr_95_5, addr_positional[1527:1524], addr_381_6);

wire[27:0] addr_382_6;

Selector_2 s382_6(wires_95_5[2], addr_95_5, addr_positional[1531:1528], addr_382_6);

wire[27:0] addr_383_6;

Selector_2 s383_6(wires_95_5[3], addr_95_5, addr_positional[1535:1532], addr_383_6);

wire[27:0] addr_384_6;

Selector_2 s384_6(wires_96_5[0], addr_96_5, addr_positional[1539:1536], addr_384_6);

wire[27:0] addr_385_6;

Selector_2 s385_6(wires_96_5[1], addr_96_5, addr_positional[1543:1540], addr_385_6);

wire[27:0] addr_386_6;

Selector_2 s386_6(wires_96_5[2], addr_96_5, addr_positional[1547:1544], addr_386_6);

wire[27:0] addr_387_6;

Selector_2 s387_6(wires_96_5[3], addr_96_5, addr_positional[1551:1548], addr_387_6);

wire[27:0] addr_388_6;

Selector_2 s388_6(wires_97_5[0], addr_97_5, addr_positional[1555:1552], addr_388_6);

wire[27:0] addr_389_6;

Selector_2 s389_6(wires_97_5[1], addr_97_5, addr_positional[1559:1556], addr_389_6);

wire[27:0] addr_390_6;

Selector_2 s390_6(wires_97_5[2], addr_97_5, addr_positional[1563:1560], addr_390_6);

wire[27:0] addr_391_6;

Selector_2 s391_6(wires_97_5[3], addr_97_5, addr_positional[1567:1564], addr_391_6);

wire[27:0] addr_392_6;

Selector_2 s392_6(wires_98_5[0], addr_98_5, addr_positional[1571:1568], addr_392_6);

wire[27:0] addr_393_6;

Selector_2 s393_6(wires_98_5[1], addr_98_5, addr_positional[1575:1572], addr_393_6);

wire[27:0] addr_394_6;

Selector_2 s394_6(wires_98_5[2], addr_98_5, addr_positional[1579:1576], addr_394_6);

wire[27:0] addr_395_6;

Selector_2 s395_6(wires_98_5[3], addr_98_5, addr_positional[1583:1580], addr_395_6);

wire[27:0] addr_396_6;

Selector_2 s396_6(wires_99_5[0], addr_99_5, addr_positional[1587:1584], addr_396_6);

wire[27:0] addr_397_6;

Selector_2 s397_6(wires_99_5[1], addr_99_5, addr_positional[1591:1588], addr_397_6);

wire[27:0] addr_398_6;

Selector_2 s398_6(wires_99_5[2], addr_99_5, addr_positional[1595:1592], addr_398_6);

wire[27:0] addr_399_6;

Selector_2 s399_6(wires_99_5[3], addr_99_5, addr_positional[1599:1596], addr_399_6);

wire[27:0] addr_400_6;

Selector_2 s400_6(wires_100_5[0], addr_100_5, addr_positional[1603:1600], addr_400_6);

wire[27:0] addr_401_6;

Selector_2 s401_6(wires_100_5[1], addr_100_5, addr_positional[1607:1604], addr_401_6);

wire[27:0] addr_402_6;

Selector_2 s402_6(wires_100_5[2], addr_100_5, addr_positional[1611:1608], addr_402_6);

wire[27:0] addr_403_6;

Selector_2 s403_6(wires_100_5[3], addr_100_5, addr_positional[1615:1612], addr_403_6);

wire[27:0] addr_404_6;

Selector_2 s404_6(wires_101_5[0], addr_101_5, addr_positional[1619:1616], addr_404_6);

wire[27:0] addr_405_6;

Selector_2 s405_6(wires_101_5[1], addr_101_5, addr_positional[1623:1620], addr_405_6);

wire[27:0] addr_406_6;

Selector_2 s406_6(wires_101_5[2], addr_101_5, addr_positional[1627:1624], addr_406_6);

wire[27:0] addr_407_6;

Selector_2 s407_6(wires_101_5[3], addr_101_5, addr_positional[1631:1628], addr_407_6);

wire[27:0] addr_408_6;

Selector_2 s408_6(wires_102_5[0], addr_102_5, addr_positional[1635:1632], addr_408_6);

wire[27:0] addr_409_6;

Selector_2 s409_6(wires_102_5[1], addr_102_5, addr_positional[1639:1636], addr_409_6);

wire[27:0] addr_410_6;

Selector_2 s410_6(wires_102_5[2], addr_102_5, addr_positional[1643:1640], addr_410_6);

wire[27:0] addr_411_6;

Selector_2 s411_6(wires_102_5[3], addr_102_5, addr_positional[1647:1644], addr_411_6);

wire[27:0] addr_412_6;

Selector_2 s412_6(wires_103_5[0], addr_103_5, addr_positional[1651:1648], addr_412_6);

wire[27:0] addr_413_6;

Selector_2 s413_6(wires_103_5[1], addr_103_5, addr_positional[1655:1652], addr_413_6);

wire[27:0] addr_414_6;

Selector_2 s414_6(wires_103_5[2], addr_103_5, addr_positional[1659:1656], addr_414_6);

wire[27:0] addr_415_6;

Selector_2 s415_6(wires_103_5[3], addr_103_5, addr_positional[1663:1660], addr_415_6);

wire[27:0] addr_416_6;

Selector_2 s416_6(wires_104_5[0], addr_104_5, addr_positional[1667:1664], addr_416_6);

wire[27:0] addr_417_6;

Selector_2 s417_6(wires_104_5[1], addr_104_5, addr_positional[1671:1668], addr_417_6);

wire[27:0] addr_418_6;

Selector_2 s418_6(wires_104_5[2], addr_104_5, addr_positional[1675:1672], addr_418_6);

wire[27:0] addr_419_6;

Selector_2 s419_6(wires_104_5[3], addr_104_5, addr_positional[1679:1676], addr_419_6);

wire[27:0] addr_420_6;

Selector_2 s420_6(wires_105_5[0], addr_105_5, addr_positional[1683:1680], addr_420_6);

wire[27:0] addr_421_6;

Selector_2 s421_6(wires_105_5[1], addr_105_5, addr_positional[1687:1684], addr_421_6);

wire[27:0] addr_422_6;

Selector_2 s422_6(wires_105_5[2], addr_105_5, addr_positional[1691:1688], addr_422_6);

wire[27:0] addr_423_6;

Selector_2 s423_6(wires_105_5[3], addr_105_5, addr_positional[1695:1692], addr_423_6);

wire[27:0] addr_424_6;

Selector_2 s424_6(wires_106_5[0], addr_106_5, addr_positional[1699:1696], addr_424_6);

wire[27:0] addr_425_6;

Selector_2 s425_6(wires_106_5[1], addr_106_5, addr_positional[1703:1700], addr_425_6);

wire[27:0] addr_426_6;

Selector_2 s426_6(wires_106_5[2], addr_106_5, addr_positional[1707:1704], addr_426_6);

wire[27:0] addr_427_6;

Selector_2 s427_6(wires_106_5[3], addr_106_5, addr_positional[1711:1708], addr_427_6);

wire[27:0] addr_428_6;

Selector_2 s428_6(wires_107_5[0], addr_107_5, addr_positional[1715:1712], addr_428_6);

wire[27:0] addr_429_6;

Selector_2 s429_6(wires_107_5[1], addr_107_5, addr_positional[1719:1716], addr_429_6);

wire[27:0] addr_430_6;

Selector_2 s430_6(wires_107_5[2], addr_107_5, addr_positional[1723:1720], addr_430_6);

wire[27:0] addr_431_6;

Selector_2 s431_6(wires_107_5[3], addr_107_5, addr_positional[1727:1724], addr_431_6);

wire[27:0] addr_432_6;

Selector_2 s432_6(wires_108_5[0], addr_108_5, addr_positional[1731:1728], addr_432_6);

wire[27:0] addr_433_6;

Selector_2 s433_6(wires_108_5[1], addr_108_5, addr_positional[1735:1732], addr_433_6);

wire[27:0] addr_434_6;

Selector_2 s434_6(wires_108_5[2], addr_108_5, addr_positional[1739:1736], addr_434_6);

wire[27:0] addr_435_6;

Selector_2 s435_6(wires_108_5[3], addr_108_5, addr_positional[1743:1740], addr_435_6);

wire[27:0] addr_436_6;

Selector_2 s436_6(wires_109_5[0], addr_109_5, addr_positional[1747:1744], addr_436_6);

wire[27:0] addr_437_6;

Selector_2 s437_6(wires_109_5[1], addr_109_5, addr_positional[1751:1748], addr_437_6);

wire[27:0] addr_438_6;

Selector_2 s438_6(wires_109_5[2], addr_109_5, addr_positional[1755:1752], addr_438_6);

wire[27:0] addr_439_6;

Selector_2 s439_6(wires_109_5[3], addr_109_5, addr_positional[1759:1756], addr_439_6);

wire[27:0] addr_440_6;

Selector_2 s440_6(wires_110_5[0], addr_110_5, addr_positional[1763:1760], addr_440_6);

wire[27:0] addr_441_6;

Selector_2 s441_6(wires_110_5[1], addr_110_5, addr_positional[1767:1764], addr_441_6);

wire[27:0] addr_442_6;

Selector_2 s442_6(wires_110_5[2], addr_110_5, addr_positional[1771:1768], addr_442_6);

wire[27:0] addr_443_6;

Selector_2 s443_6(wires_110_5[3], addr_110_5, addr_positional[1775:1772], addr_443_6);

wire[27:0] addr_444_6;

Selector_2 s444_6(wires_111_5[0], addr_111_5, addr_positional[1779:1776], addr_444_6);

wire[27:0] addr_445_6;

Selector_2 s445_6(wires_111_5[1], addr_111_5, addr_positional[1783:1780], addr_445_6);

wire[27:0] addr_446_6;

Selector_2 s446_6(wires_111_5[2], addr_111_5, addr_positional[1787:1784], addr_446_6);

wire[27:0] addr_447_6;

Selector_2 s447_6(wires_111_5[3], addr_111_5, addr_positional[1791:1788], addr_447_6);

wire[27:0] addr_448_6;

Selector_2 s448_6(wires_112_5[0], addr_112_5, addr_positional[1795:1792], addr_448_6);

wire[27:0] addr_449_6;

Selector_2 s449_6(wires_112_5[1], addr_112_5, addr_positional[1799:1796], addr_449_6);

wire[27:0] addr_450_6;

Selector_2 s450_6(wires_112_5[2], addr_112_5, addr_positional[1803:1800], addr_450_6);

wire[27:0] addr_451_6;

Selector_2 s451_6(wires_112_5[3], addr_112_5, addr_positional[1807:1804], addr_451_6);

wire[27:0] addr_452_6;

Selector_2 s452_6(wires_113_5[0], addr_113_5, addr_positional[1811:1808], addr_452_6);

wire[27:0] addr_453_6;

Selector_2 s453_6(wires_113_5[1], addr_113_5, addr_positional[1815:1812], addr_453_6);

wire[27:0] addr_454_6;

Selector_2 s454_6(wires_113_5[2], addr_113_5, addr_positional[1819:1816], addr_454_6);

wire[27:0] addr_455_6;

Selector_2 s455_6(wires_113_5[3], addr_113_5, addr_positional[1823:1820], addr_455_6);

wire[27:0] addr_456_6;

Selector_2 s456_6(wires_114_5[0], addr_114_5, addr_positional[1827:1824], addr_456_6);

wire[27:0] addr_457_6;

Selector_2 s457_6(wires_114_5[1], addr_114_5, addr_positional[1831:1828], addr_457_6);

wire[27:0] addr_458_6;

Selector_2 s458_6(wires_114_5[2], addr_114_5, addr_positional[1835:1832], addr_458_6);

wire[27:0] addr_459_6;

Selector_2 s459_6(wires_114_5[3], addr_114_5, addr_positional[1839:1836], addr_459_6);

wire[27:0] addr_460_6;

Selector_2 s460_6(wires_115_5[0], addr_115_5, addr_positional[1843:1840], addr_460_6);

wire[27:0] addr_461_6;

Selector_2 s461_6(wires_115_5[1], addr_115_5, addr_positional[1847:1844], addr_461_6);

wire[27:0] addr_462_6;

Selector_2 s462_6(wires_115_5[2], addr_115_5, addr_positional[1851:1848], addr_462_6);

wire[27:0] addr_463_6;

Selector_2 s463_6(wires_115_5[3], addr_115_5, addr_positional[1855:1852], addr_463_6);

wire[27:0] addr_464_6;

Selector_2 s464_6(wires_116_5[0], addr_116_5, addr_positional[1859:1856], addr_464_6);

wire[27:0] addr_465_6;

Selector_2 s465_6(wires_116_5[1], addr_116_5, addr_positional[1863:1860], addr_465_6);

wire[27:0] addr_466_6;

Selector_2 s466_6(wires_116_5[2], addr_116_5, addr_positional[1867:1864], addr_466_6);

wire[27:0] addr_467_6;

Selector_2 s467_6(wires_116_5[3], addr_116_5, addr_positional[1871:1868], addr_467_6);

wire[27:0] addr_468_6;

Selector_2 s468_6(wires_117_5[0], addr_117_5, addr_positional[1875:1872], addr_468_6);

wire[27:0] addr_469_6;

Selector_2 s469_6(wires_117_5[1], addr_117_5, addr_positional[1879:1876], addr_469_6);

wire[27:0] addr_470_6;

Selector_2 s470_6(wires_117_5[2], addr_117_5, addr_positional[1883:1880], addr_470_6);

wire[27:0] addr_471_6;

Selector_2 s471_6(wires_117_5[3], addr_117_5, addr_positional[1887:1884], addr_471_6);

wire[27:0] addr_472_6;

Selector_2 s472_6(wires_118_5[0], addr_118_5, addr_positional[1891:1888], addr_472_6);

wire[27:0] addr_473_6;

Selector_2 s473_6(wires_118_5[1], addr_118_5, addr_positional[1895:1892], addr_473_6);

wire[27:0] addr_474_6;

Selector_2 s474_6(wires_118_5[2], addr_118_5, addr_positional[1899:1896], addr_474_6);

wire[27:0] addr_475_6;

Selector_2 s475_6(wires_118_5[3], addr_118_5, addr_positional[1903:1900], addr_475_6);

wire[27:0] addr_476_6;

Selector_2 s476_6(wires_119_5[0], addr_119_5, addr_positional[1907:1904], addr_476_6);

wire[27:0] addr_477_6;

Selector_2 s477_6(wires_119_5[1], addr_119_5, addr_positional[1911:1908], addr_477_6);

wire[27:0] addr_478_6;

Selector_2 s478_6(wires_119_5[2], addr_119_5, addr_positional[1915:1912], addr_478_6);

wire[27:0] addr_479_6;

Selector_2 s479_6(wires_119_5[3], addr_119_5, addr_positional[1919:1916], addr_479_6);

wire[27:0] addr_480_6;

Selector_2 s480_6(wires_120_5[0], addr_120_5, addr_positional[1923:1920], addr_480_6);

wire[27:0] addr_481_6;

Selector_2 s481_6(wires_120_5[1], addr_120_5, addr_positional[1927:1924], addr_481_6);

wire[27:0] addr_482_6;

Selector_2 s482_6(wires_120_5[2], addr_120_5, addr_positional[1931:1928], addr_482_6);

wire[27:0] addr_483_6;

Selector_2 s483_6(wires_120_5[3], addr_120_5, addr_positional[1935:1932], addr_483_6);

wire[27:0] addr_484_6;

Selector_2 s484_6(wires_121_5[0], addr_121_5, addr_positional[1939:1936], addr_484_6);

wire[27:0] addr_485_6;

Selector_2 s485_6(wires_121_5[1], addr_121_5, addr_positional[1943:1940], addr_485_6);

wire[27:0] addr_486_6;

Selector_2 s486_6(wires_121_5[2], addr_121_5, addr_positional[1947:1944], addr_486_6);

wire[27:0] addr_487_6;

Selector_2 s487_6(wires_121_5[3], addr_121_5, addr_positional[1951:1948], addr_487_6);

wire[27:0] addr_488_6;

Selector_2 s488_6(wires_122_5[0], addr_122_5, addr_positional[1955:1952], addr_488_6);

wire[27:0] addr_489_6;

Selector_2 s489_6(wires_122_5[1], addr_122_5, addr_positional[1959:1956], addr_489_6);

wire[27:0] addr_490_6;

Selector_2 s490_6(wires_122_5[2], addr_122_5, addr_positional[1963:1960], addr_490_6);

wire[27:0] addr_491_6;

Selector_2 s491_6(wires_122_5[3], addr_122_5, addr_positional[1967:1964], addr_491_6);

wire[27:0] addr_492_6;

Selector_2 s492_6(wires_123_5[0], addr_123_5, addr_positional[1971:1968], addr_492_6);

wire[27:0] addr_493_6;

Selector_2 s493_6(wires_123_5[1], addr_123_5, addr_positional[1975:1972], addr_493_6);

wire[27:0] addr_494_6;

Selector_2 s494_6(wires_123_5[2], addr_123_5, addr_positional[1979:1976], addr_494_6);

wire[27:0] addr_495_6;

Selector_2 s495_6(wires_123_5[3], addr_123_5, addr_positional[1983:1980], addr_495_6);

wire[27:0] addr_496_6;

Selector_2 s496_6(wires_124_5[0], addr_124_5, addr_positional[1987:1984], addr_496_6);

wire[27:0] addr_497_6;

Selector_2 s497_6(wires_124_5[1], addr_124_5, addr_positional[1991:1988], addr_497_6);

wire[27:0] addr_498_6;

Selector_2 s498_6(wires_124_5[2], addr_124_5, addr_positional[1995:1992], addr_498_6);

wire[27:0] addr_499_6;

Selector_2 s499_6(wires_124_5[3], addr_124_5, addr_positional[1999:1996], addr_499_6);

wire[27:0] addr_500_6;

Selector_2 s500_6(wires_125_5[0], addr_125_5, addr_positional[2003:2000], addr_500_6);

wire[27:0] addr_501_6;

Selector_2 s501_6(wires_125_5[1], addr_125_5, addr_positional[2007:2004], addr_501_6);

wire[27:0] addr_502_6;

Selector_2 s502_6(wires_125_5[2], addr_125_5, addr_positional[2011:2008], addr_502_6);

wire[27:0] addr_503_6;

Selector_2 s503_6(wires_125_5[3], addr_125_5, addr_positional[2015:2012], addr_503_6);

wire[27:0] addr_504_6;

Selector_2 s504_6(wires_126_5[0], addr_126_5, addr_positional[2019:2016], addr_504_6);

wire[27:0] addr_505_6;

Selector_2 s505_6(wires_126_5[1], addr_126_5, addr_positional[2023:2020], addr_505_6);

wire[27:0] addr_506_6;

Selector_2 s506_6(wires_126_5[2], addr_126_5, addr_positional[2027:2024], addr_506_6);

wire[27:0] addr_507_6;

Selector_2 s507_6(wires_126_5[3], addr_126_5, addr_positional[2031:2028], addr_507_6);

wire[27:0] addr_508_6;

Selector_2 s508_6(wires_127_5[0], addr_127_5, addr_positional[2035:2032], addr_508_6);

wire[27:0] addr_509_6;

Selector_2 s509_6(wires_127_5[1], addr_127_5, addr_positional[2039:2036], addr_509_6);

wire[27:0] addr_510_6;

Selector_2 s510_6(wires_127_5[2], addr_127_5, addr_positional[2043:2040], addr_510_6);

wire[27:0] addr_511_6;

Selector_2 s511_6(wires_127_5[3], addr_127_5, addr_positional[2047:2044], addr_511_6);

wire[27:0] addr_512_6;

Selector_2 s512_6(wires_128_5[0], addr_128_5, addr_positional[2051:2048], addr_512_6);

wire[27:0] addr_513_6;

Selector_2 s513_6(wires_128_5[1], addr_128_5, addr_positional[2055:2052], addr_513_6);

wire[27:0] addr_514_6;

Selector_2 s514_6(wires_128_5[2], addr_128_5, addr_positional[2059:2056], addr_514_6);

wire[27:0] addr_515_6;

Selector_2 s515_6(wires_128_5[3], addr_128_5, addr_positional[2063:2060], addr_515_6);

wire[27:0] addr_516_6;

Selector_2 s516_6(wires_129_5[0], addr_129_5, addr_positional[2067:2064], addr_516_6);

wire[27:0] addr_517_6;

Selector_2 s517_6(wires_129_5[1], addr_129_5, addr_positional[2071:2068], addr_517_6);

wire[27:0] addr_518_6;

Selector_2 s518_6(wires_129_5[2], addr_129_5, addr_positional[2075:2072], addr_518_6);

wire[27:0] addr_519_6;

Selector_2 s519_6(wires_129_5[3], addr_129_5, addr_positional[2079:2076], addr_519_6);

wire[27:0] addr_520_6;

Selector_2 s520_6(wires_130_5[0], addr_130_5, addr_positional[2083:2080], addr_520_6);

wire[27:0] addr_521_6;

Selector_2 s521_6(wires_130_5[1], addr_130_5, addr_positional[2087:2084], addr_521_6);

wire[27:0] addr_522_6;

Selector_2 s522_6(wires_130_5[2], addr_130_5, addr_positional[2091:2088], addr_522_6);

wire[27:0] addr_523_6;

Selector_2 s523_6(wires_130_5[3], addr_130_5, addr_positional[2095:2092], addr_523_6);

wire[27:0] addr_524_6;

Selector_2 s524_6(wires_131_5[0], addr_131_5, addr_positional[2099:2096], addr_524_6);

wire[27:0] addr_525_6;

Selector_2 s525_6(wires_131_5[1], addr_131_5, addr_positional[2103:2100], addr_525_6);

wire[27:0] addr_526_6;

Selector_2 s526_6(wires_131_5[2], addr_131_5, addr_positional[2107:2104], addr_526_6);

wire[27:0] addr_527_6;

Selector_2 s527_6(wires_131_5[3], addr_131_5, addr_positional[2111:2108], addr_527_6);

wire[27:0] addr_528_6;

Selector_2 s528_6(wires_132_5[0], addr_132_5, addr_positional[2115:2112], addr_528_6);

wire[27:0] addr_529_6;

Selector_2 s529_6(wires_132_5[1], addr_132_5, addr_positional[2119:2116], addr_529_6);

wire[27:0] addr_530_6;

Selector_2 s530_6(wires_132_5[2], addr_132_5, addr_positional[2123:2120], addr_530_6);

wire[27:0] addr_531_6;

Selector_2 s531_6(wires_132_5[3], addr_132_5, addr_positional[2127:2124], addr_531_6);

wire[27:0] addr_532_6;

Selector_2 s532_6(wires_133_5[0], addr_133_5, addr_positional[2131:2128], addr_532_6);

wire[27:0] addr_533_6;

Selector_2 s533_6(wires_133_5[1], addr_133_5, addr_positional[2135:2132], addr_533_6);

wire[27:0] addr_534_6;

Selector_2 s534_6(wires_133_5[2], addr_133_5, addr_positional[2139:2136], addr_534_6);

wire[27:0] addr_535_6;

Selector_2 s535_6(wires_133_5[3], addr_133_5, addr_positional[2143:2140], addr_535_6);

wire[27:0] addr_536_6;

Selector_2 s536_6(wires_134_5[0], addr_134_5, addr_positional[2147:2144], addr_536_6);

wire[27:0] addr_537_6;

Selector_2 s537_6(wires_134_5[1], addr_134_5, addr_positional[2151:2148], addr_537_6);

wire[27:0] addr_538_6;

Selector_2 s538_6(wires_134_5[2], addr_134_5, addr_positional[2155:2152], addr_538_6);

wire[27:0] addr_539_6;

Selector_2 s539_6(wires_134_5[3], addr_134_5, addr_positional[2159:2156], addr_539_6);

wire[27:0] addr_540_6;

Selector_2 s540_6(wires_135_5[0], addr_135_5, addr_positional[2163:2160], addr_540_6);

wire[27:0] addr_541_6;

Selector_2 s541_6(wires_135_5[1], addr_135_5, addr_positional[2167:2164], addr_541_6);

wire[27:0] addr_542_6;

Selector_2 s542_6(wires_135_5[2], addr_135_5, addr_positional[2171:2168], addr_542_6);

wire[27:0] addr_543_6;

Selector_2 s543_6(wires_135_5[3], addr_135_5, addr_positional[2175:2172], addr_543_6);

wire[27:0] addr_544_6;

Selector_2 s544_6(wires_136_5[0], addr_136_5, addr_positional[2179:2176], addr_544_6);

wire[27:0] addr_545_6;

Selector_2 s545_6(wires_136_5[1], addr_136_5, addr_positional[2183:2180], addr_545_6);

wire[27:0] addr_546_6;

Selector_2 s546_6(wires_136_5[2], addr_136_5, addr_positional[2187:2184], addr_546_6);

wire[27:0] addr_547_6;

Selector_2 s547_6(wires_136_5[3], addr_136_5, addr_positional[2191:2188], addr_547_6);

wire[27:0] addr_548_6;

Selector_2 s548_6(wires_137_5[0], addr_137_5, addr_positional[2195:2192], addr_548_6);

wire[27:0] addr_549_6;

Selector_2 s549_6(wires_137_5[1], addr_137_5, addr_positional[2199:2196], addr_549_6);

wire[27:0] addr_550_6;

Selector_2 s550_6(wires_137_5[2], addr_137_5, addr_positional[2203:2200], addr_550_6);

wire[27:0] addr_551_6;

Selector_2 s551_6(wires_137_5[3], addr_137_5, addr_positional[2207:2204], addr_551_6);

wire[27:0] addr_552_6;

Selector_2 s552_6(wires_138_5[0], addr_138_5, addr_positional[2211:2208], addr_552_6);

wire[27:0] addr_553_6;

Selector_2 s553_6(wires_138_5[1], addr_138_5, addr_positional[2215:2212], addr_553_6);

wire[27:0] addr_554_6;

Selector_2 s554_6(wires_138_5[2], addr_138_5, addr_positional[2219:2216], addr_554_6);

wire[27:0] addr_555_6;

Selector_2 s555_6(wires_138_5[3], addr_138_5, addr_positional[2223:2220], addr_555_6);

wire[27:0] addr_556_6;

Selector_2 s556_6(wires_139_5[0], addr_139_5, addr_positional[2227:2224], addr_556_6);

wire[27:0] addr_557_6;

Selector_2 s557_6(wires_139_5[1], addr_139_5, addr_positional[2231:2228], addr_557_6);

wire[27:0] addr_558_6;

Selector_2 s558_6(wires_139_5[2], addr_139_5, addr_positional[2235:2232], addr_558_6);

wire[27:0] addr_559_6;

Selector_2 s559_6(wires_139_5[3], addr_139_5, addr_positional[2239:2236], addr_559_6);

wire[27:0] addr_560_6;

Selector_2 s560_6(wires_140_5[0], addr_140_5, addr_positional[2243:2240], addr_560_6);

wire[27:0] addr_561_6;

Selector_2 s561_6(wires_140_5[1], addr_140_5, addr_positional[2247:2244], addr_561_6);

wire[27:0] addr_562_6;

Selector_2 s562_6(wires_140_5[2], addr_140_5, addr_positional[2251:2248], addr_562_6);

wire[27:0] addr_563_6;

Selector_2 s563_6(wires_140_5[3], addr_140_5, addr_positional[2255:2252], addr_563_6);

wire[27:0] addr_564_6;

Selector_2 s564_6(wires_141_5[0], addr_141_5, addr_positional[2259:2256], addr_564_6);

wire[27:0] addr_565_6;

Selector_2 s565_6(wires_141_5[1], addr_141_5, addr_positional[2263:2260], addr_565_6);

wire[27:0] addr_566_6;

Selector_2 s566_6(wires_141_5[2], addr_141_5, addr_positional[2267:2264], addr_566_6);

wire[27:0] addr_567_6;

Selector_2 s567_6(wires_141_5[3], addr_141_5, addr_positional[2271:2268], addr_567_6);

wire[27:0] addr_568_6;

Selector_2 s568_6(wires_142_5[0], addr_142_5, addr_positional[2275:2272], addr_568_6);

wire[27:0] addr_569_6;

Selector_2 s569_6(wires_142_5[1], addr_142_5, addr_positional[2279:2276], addr_569_6);

wire[27:0] addr_570_6;

Selector_2 s570_6(wires_142_5[2], addr_142_5, addr_positional[2283:2280], addr_570_6);

wire[27:0] addr_571_6;

Selector_2 s571_6(wires_142_5[3], addr_142_5, addr_positional[2287:2284], addr_571_6);

wire[27:0] addr_572_6;

Selector_2 s572_6(wires_143_5[0], addr_143_5, addr_positional[2291:2288], addr_572_6);

wire[27:0] addr_573_6;

Selector_2 s573_6(wires_143_5[1], addr_143_5, addr_positional[2295:2292], addr_573_6);

wire[27:0] addr_574_6;

Selector_2 s574_6(wires_143_5[2], addr_143_5, addr_positional[2299:2296], addr_574_6);

wire[27:0] addr_575_6;

Selector_2 s575_6(wires_143_5[3], addr_143_5, addr_positional[2303:2300], addr_575_6);

wire[27:0] addr_576_6;

Selector_2 s576_6(wires_144_5[0], addr_144_5, addr_positional[2307:2304], addr_576_6);

wire[27:0] addr_577_6;

Selector_2 s577_6(wires_144_5[1], addr_144_5, addr_positional[2311:2308], addr_577_6);

wire[27:0] addr_578_6;

Selector_2 s578_6(wires_144_5[2], addr_144_5, addr_positional[2315:2312], addr_578_6);

wire[27:0] addr_579_6;

Selector_2 s579_6(wires_144_5[3], addr_144_5, addr_positional[2319:2316], addr_579_6);

wire[27:0] addr_580_6;

Selector_2 s580_6(wires_145_5[0], addr_145_5, addr_positional[2323:2320], addr_580_6);

wire[27:0] addr_581_6;

Selector_2 s581_6(wires_145_5[1], addr_145_5, addr_positional[2327:2324], addr_581_6);

wire[27:0] addr_582_6;

Selector_2 s582_6(wires_145_5[2], addr_145_5, addr_positional[2331:2328], addr_582_6);

wire[27:0] addr_583_6;

Selector_2 s583_6(wires_145_5[3], addr_145_5, addr_positional[2335:2332], addr_583_6);

wire[27:0] addr_584_6;

Selector_2 s584_6(wires_146_5[0], addr_146_5, addr_positional[2339:2336], addr_584_6);

wire[27:0] addr_585_6;

Selector_2 s585_6(wires_146_5[1], addr_146_5, addr_positional[2343:2340], addr_585_6);

wire[27:0] addr_586_6;

Selector_2 s586_6(wires_146_5[2], addr_146_5, addr_positional[2347:2344], addr_586_6);

wire[27:0] addr_587_6;

Selector_2 s587_6(wires_146_5[3], addr_146_5, addr_positional[2351:2348], addr_587_6);

wire[27:0] addr_588_6;

Selector_2 s588_6(wires_147_5[0], addr_147_5, addr_positional[2355:2352], addr_588_6);

wire[27:0] addr_589_6;

Selector_2 s589_6(wires_147_5[1], addr_147_5, addr_positional[2359:2356], addr_589_6);

wire[27:0] addr_590_6;

Selector_2 s590_6(wires_147_5[2], addr_147_5, addr_positional[2363:2360], addr_590_6);

wire[27:0] addr_591_6;

Selector_2 s591_6(wires_147_5[3], addr_147_5, addr_positional[2367:2364], addr_591_6);

wire[27:0] addr_592_6;

Selector_2 s592_6(wires_148_5[0], addr_148_5, addr_positional[2371:2368], addr_592_6);

wire[27:0] addr_593_6;

Selector_2 s593_6(wires_148_5[1], addr_148_5, addr_positional[2375:2372], addr_593_6);

wire[27:0] addr_594_6;

Selector_2 s594_6(wires_148_5[2], addr_148_5, addr_positional[2379:2376], addr_594_6);

wire[27:0] addr_595_6;

Selector_2 s595_6(wires_148_5[3], addr_148_5, addr_positional[2383:2380], addr_595_6);

wire[27:0] addr_596_6;

Selector_2 s596_6(wires_149_5[0], addr_149_5, addr_positional[2387:2384], addr_596_6);

wire[27:0] addr_597_6;

Selector_2 s597_6(wires_149_5[1], addr_149_5, addr_positional[2391:2388], addr_597_6);

wire[27:0] addr_598_6;

Selector_2 s598_6(wires_149_5[2], addr_149_5, addr_positional[2395:2392], addr_598_6);

wire[27:0] addr_599_6;

Selector_2 s599_6(wires_149_5[3], addr_149_5, addr_positional[2399:2396], addr_599_6);

wire[27:0] addr_600_6;

Selector_2 s600_6(wires_150_5[0], addr_150_5, addr_positional[2403:2400], addr_600_6);

wire[27:0] addr_601_6;

Selector_2 s601_6(wires_150_5[1], addr_150_5, addr_positional[2407:2404], addr_601_6);

wire[27:0] addr_602_6;

Selector_2 s602_6(wires_150_5[2], addr_150_5, addr_positional[2411:2408], addr_602_6);

wire[27:0] addr_603_6;

Selector_2 s603_6(wires_150_5[3], addr_150_5, addr_positional[2415:2412], addr_603_6);

wire[27:0] addr_604_6;

Selector_2 s604_6(wires_151_5[0], addr_151_5, addr_positional[2419:2416], addr_604_6);

wire[27:0] addr_605_6;

Selector_2 s605_6(wires_151_5[1], addr_151_5, addr_positional[2423:2420], addr_605_6);

wire[27:0] addr_606_6;

Selector_2 s606_6(wires_151_5[2], addr_151_5, addr_positional[2427:2424], addr_606_6);

wire[27:0] addr_607_6;

Selector_2 s607_6(wires_151_5[3], addr_151_5, addr_positional[2431:2428], addr_607_6);

wire[27:0] addr_608_6;

Selector_2 s608_6(wires_152_5[0], addr_152_5, addr_positional[2435:2432], addr_608_6);

wire[27:0] addr_609_6;

Selector_2 s609_6(wires_152_5[1], addr_152_5, addr_positional[2439:2436], addr_609_6);

wire[27:0] addr_610_6;

Selector_2 s610_6(wires_152_5[2], addr_152_5, addr_positional[2443:2440], addr_610_6);

wire[27:0] addr_611_6;

Selector_2 s611_6(wires_152_5[3], addr_152_5, addr_positional[2447:2444], addr_611_6);

wire[27:0] addr_612_6;

Selector_2 s612_6(wires_153_5[0], addr_153_5, addr_positional[2451:2448], addr_612_6);

wire[27:0] addr_613_6;

Selector_2 s613_6(wires_153_5[1], addr_153_5, addr_positional[2455:2452], addr_613_6);

wire[27:0] addr_614_6;

Selector_2 s614_6(wires_153_5[2], addr_153_5, addr_positional[2459:2456], addr_614_6);

wire[27:0] addr_615_6;

Selector_2 s615_6(wires_153_5[3], addr_153_5, addr_positional[2463:2460], addr_615_6);

wire[27:0] addr_616_6;

Selector_2 s616_6(wires_154_5[0], addr_154_5, addr_positional[2467:2464], addr_616_6);

wire[27:0] addr_617_6;

Selector_2 s617_6(wires_154_5[1], addr_154_5, addr_positional[2471:2468], addr_617_6);

wire[27:0] addr_618_6;

Selector_2 s618_6(wires_154_5[2], addr_154_5, addr_positional[2475:2472], addr_618_6);

wire[27:0] addr_619_6;

Selector_2 s619_6(wires_154_5[3], addr_154_5, addr_positional[2479:2476], addr_619_6);

wire[27:0] addr_620_6;

Selector_2 s620_6(wires_155_5[0], addr_155_5, addr_positional[2483:2480], addr_620_6);

wire[27:0] addr_621_6;

Selector_2 s621_6(wires_155_5[1], addr_155_5, addr_positional[2487:2484], addr_621_6);

wire[27:0] addr_622_6;

Selector_2 s622_6(wires_155_5[2], addr_155_5, addr_positional[2491:2488], addr_622_6);

wire[27:0] addr_623_6;

Selector_2 s623_6(wires_155_5[3], addr_155_5, addr_positional[2495:2492], addr_623_6);

wire[27:0] addr_624_6;

Selector_2 s624_6(wires_156_5[0], addr_156_5, addr_positional[2499:2496], addr_624_6);

wire[27:0] addr_625_6;

Selector_2 s625_6(wires_156_5[1], addr_156_5, addr_positional[2503:2500], addr_625_6);

wire[27:0] addr_626_6;

Selector_2 s626_6(wires_156_5[2], addr_156_5, addr_positional[2507:2504], addr_626_6);

wire[27:0] addr_627_6;

Selector_2 s627_6(wires_156_5[3], addr_156_5, addr_positional[2511:2508], addr_627_6);

wire[27:0] addr_628_6;

Selector_2 s628_6(wires_157_5[0], addr_157_5, addr_positional[2515:2512], addr_628_6);

wire[27:0] addr_629_6;

Selector_2 s629_6(wires_157_5[1], addr_157_5, addr_positional[2519:2516], addr_629_6);

wire[27:0] addr_630_6;

Selector_2 s630_6(wires_157_5[2], addr_157_5, addr_positional[2523:2520], addr_630_6);

wire[27:0] addr_631_6;

Selector_2 s631_6(wires_157_5[3], addr_157_5, addr_positional[2527:2524], addr_631_6);

wire[27:0] addr_632_6;

Selector_2 s632_6(wires_158_5[0], addr_158_5, addr_positional[2531:2528], addr_632_6);

wire[27:0] addr_633_6;

Selector_2 s633_6(wires_158_5[1], addr_158_5, addr_positional[2535:2532], addr_633_6);

wire[27:0] addr_634_6;

Selector_2 s634_6(wires_158_5[2], addr_158_5, addr_positional[2539:2536], addr_634_6);

wire[27:0] addr_635_6;

Selector_2 s635_6(wires_158_5[3], addr_158_5, addr_positional[2543:2540], addr_635_6);

wire[27:0] addr_636_6;

Selector_2 s636_6(wires_159_5[0], addr_159_5, addr_positional[2547:2544], addr_636_6);

wire[27:0] addr_637_6;

Selector_2 s637_6(wires_159_5[1], addr_159_5, addr_positional[2551:2548], addr_637_6);

wire[27:0] addr_638_6;

Selector_2 s638_6(wires_159_5[2], addr_159_5, addr_positional[2555:2552], addr_638_6);

wire[27:0] addr_639_6;

Selector_2 s639_6(wires_159_5[3], addr_159_5, addr_positional[2559:2556], addr_639_6);

wire[27:0] addr_640_6;

Selector_2 s640_6(wires_160_5[0], addr_160_5, addr_positional[2563:2560], addr_640_6);

wire[27:0] addr_641_6;

Selector_2 s641_6(wires_160_5[1], addr_160_5, addr_positional[2567:2564], addr_641_6);

wire[27:0] addr_642_6;

Selector_2 s642_6(wires_160_5[2], addr_160_5, addr_positional[2571:2568], addr_642_6);

wire[27:0] addr_643_6;

Selector_2 s643_6(wires_160_5[3], addr_160_5, addr_positional[2575:2572], addr_643_6);

wire[27:0] addr_644_6;

Selector_2 s644_6(wires_161_5[0], addr_161_5, addr_positional[2579:2576], addr_644_6);

wire[27:0] addr_645_6;

Selector_2 s645_6(wires_161_5[1], addr_161_5, addr_positional[2583:2580], addr_645_6);

wire[27:0] addr_646_6;

Selector_2 s646_6(wires_161_5[2], addr_161_5, addr_positional[2587:2584], addr_646_6);

wire[27:0] addr_647_6;

Selector_2 s647_6(wires_161_5[3], addr_161_5, addr_positional[2591:2588], addr_647_6);

wire[27:0] addr_648_6;

Selector_2 s648_6(wires_162_5[0], addr_162_5, addr_positional[2595:2592], addr_648_6);

wire[27:0] addr_649_6;

Selector_2 s649_6(wires_162_5[1], addr_162_5, addr_positional[2599:2596], addr_649_6);

wire[27:0] addr_650_6;

Selector_2 s650_6(wires_162_5[2], addr_162_5, addr_positional[2603:2600], addr_650_6);

wire[27:0] addr_651_6;

Selector_2 s651_6(wires_162_5[3], addr_162_5, addr_positional[2607:2604], addr_651_6);

wire[27:0] addr_652_6;

Selector_2 s652_6(wires_163_5[0], addr_163_5, addr_positional[2611:2608], addr_652_6);

wire[27:0] addr_653_6;

Selector_2 s653_6(wires_163_5[1], addr_163_5, addr_positional[2615:2612], addr_653_6);

wire[27:0] addr_654_6;

Selector_2 s654_6(wires_163_5[2], addr_163_5, addr_positional[2619:2616], addr_654_6);

wire[27:0] addr_655_6;

Selector_2 s655_6(wires_163_5[3], addr_163_5, addr_positional[2623:2620], addr_655_6);

wire[27:0] addr_656_6;

Selector_2 s656_6(wires_164_5[0], addr_164_5, addr_positional[2627:2624], addr_656_6);

wire[27:0] addr_657_6;

Selector_2 s657_6(wires_164_5[1], addr_164_5, addr_positional[2631:2628], addr_657_6);

wire[27:0] addr_658_6;

Selector_2 s658_6(wires_164_5[2], addr_164_5, addr_positional[2635:2632], addr_658_6);

wire[27:0] addr_659_6;

Selector_2 s659_6(wires_164_5[3], addr_164_5, addr_positional[2639:2636], addr_659_6);

wire[27:0] addr_660_6;

Selector_2 s660_6(wires_165_5[0], addr_165_5, addr_positional[2643:2640], addr_660_6);

wire[27:0] addr_661_6;

Selector_2 s661_6(wires_165_5[1], addr_165_5, addr_positional[2647:2644], addr_661_6);

wire[27:0] addr_662_6;

Selector_2 s662_6(wires_165_5[2], addr_165_5, addr_positional[2651:2648], addr_662_6);

wire[27:0] addr_663_6;

Selector_2 s663_6(wires_165_5[3], addr_165_5, addr_positional[2655:2652], addr_663_6);

wire[27:0] addr_664_6;

Selector_2 s664_6(wires_166_5[0], addr_166_5, addr_positional[2659:2656], addr_664_6);

wire[27:0] addr_665_6;

Selector_2 s665_6(wires_166_5[1], addr_166_5, addr_positional[2663:2660], addr_665_6);

wire[27:0] addr_666_6;

Selector_2 s666_6(wires_166_5[2], addr_166_5, addr_positional[2667:2664], addr_666_6);

wire[27:0] addr_667_6;

Selector_2 s667_6(wires_166_5[3], addr_166_5, addr_positional[2671:2668], addr_667_6);

wire[27:0] addr_668_6;

Selector_2 s668_6(wires_167_5[0], addr_167_5, addr_positional[2675:2672], addr_668_6);

wire[27:0] addr_669_6;

Selector_2 s669_6(wires_167_5[1], addr_167_5, addr_positional[2679:2676], addr_669_6);

wire[27:0] addr_670_6;

Selector_2 s670_6(wires_167_5[2], addr_167_5, addr_positional[2683:2680], addr_670_6);

wire[27:0] addr_671_6;

Selector_2 s671_6(wires_167_5[3], addr_167_5, addr_positional[2687:2684], addr_671_6);

wire[27:0] addr_672_6;

Selector_2 s672_6(wires_168_5[0], addr_168_5, addr_positional[2691:2688], addr_672_6);

wire[27:0] addr_673_6;

Selector_2 s673_6(wires_168_5[1], addr_168_5, addr_positional[2695:2692], addr_673_6);

wire[27:0] addr_674_6;

Selector_2 s674_6(wires_168_5[2], addr_168_5, addr_positional[2699:2696], addr_674_6);

wire[27:0] addr_675_6;

Selector_2 s675_6(wires_168_5[3], addr_168_5, addr_positional[2703:2700], addr_675_6);

wire[27:0] addr_676_6;

Selector_2 s676_6(wires_169_5[0], addr_169_5, addr_positional[2707:2704], addr_676_6);

wire[27:0] addr_677_6;

Selector_2 s677_6(wires_169_5[1], addr_169_5, addr_positional[2711:2708], addr_677_6);

wire[27:0] addr_678_6;

Selector_2 s678_6(wires_169_5[2], addr_169_5, addr_positional[2715:2712], addr_678_6);

wire[27:0] addr_679_6;

Selector_2 s679_6(wires_169_5[3], addr_169_5, addr_positional[2719:2716], addr_679_6);

wire[27:0] addr_680_6;

Selector_2 s680_6(wires_170_5[0], addr_170_5, addr_positional[2723:2720], addr_680_6);

wire[27:0] addr_681_6;

Selector_2 s681_6(wires_170_5[1], addr_170_5, addr_positional[2727:2724], addr_681_6);

wire[27:0] addr_682_6;

Selector_2 s682_6(wires_170_5[2], addr_170_5, addr_positional[2731:2728], addr_682_6);

wire[27:0] addr_683_6;

Selector_2 s683_6(wires_170_5[3], addr_170_5, addr_positional[2735:2732], addr_683_6);

wire[27:0] addr_684_6;

Selector_2 s684_6(wires_171_5[0], addr_171_5, addr_positional[2739:2736], addr_684_6);

wire[27:0] addr_685_6;

Selector_2 s685_6(wires_171_5[1], addr_171_5, addr_positional[2743:2740], addr_685_6);

wire[27:0] addr_686_6;

Selector_2 s686_6(wires_171_5[2], addr_171_5, addr_positional[2747:2744], addr_686_6);

wire[27:0] addr_687_6;

Selector_2 s687_6(wires_171_5[3], addr_171_5, addr_positional[2751:2748], addr_687_6);

wire[27:0] addr_688_6;

Selector_2 s688_6(wires_172_5[0], addr_172_5, addr_positional[2755:2752], addr_688_6);

wire[27:0] addr_689_6;

Selector_2 s689_6(wires_172_5[1], addr_172_5, addr_positional[2759:2756], addr_689_6);

wire[27:0] addr_690_6;

Selector_2 s690_6(wires_172_5[2], addr_172_5, addr_positional[2763:2760], addr_690_6);

wire[27:0] addr_691_6;

Selector_2 s691_6(wires_172_5[3], addr_172_5, addr_positional[2767:2764], addr_691_6);

wire[27:0] addr_692_6;

Selector_2 s692_6(wires_173_5[0], addr_173_5, addr_positional[2771:2768], addr_692_6);

wire[27:0] addr_693_6;

Selector_2 s693_6(wires_173_5[1], addr_173_5, addr_positional[2775:2772], addr_693_6);

wire[27:0] addr_694_6;

Selector_2 s694_6(wires_173_5[2], addr_173_5, addr_positional[2779:2776], addr_694_6);

wire[27:0] addr_695_6;

Selector_2 s695_6(wires_173_5[3], addr_173_5, addr_positional[2783:2780], addr_695_6);

wire[27:0] addr_696_6;

Selector_2 s696_6(wires_174_5[0], addr_174_5, addr_positional[2787:2784], addr_696_6);

wire[27:0] addr_697_6;

Selector_2 s697_6(wires_174_5[1], addr_174_5, addr_positional[2791:2788], addr_697_6);

wire[27:0] addr_698_6;

Selector_2 s698_6(wires_174_5[2], addr_174_5, addr_positional[2795:2792], addr_698_6);

wire[27:0] addr_699_6;

Selector_2 s699_6(wires_174_5[3], addr_174_5, addr_positional[2799:2796], addr_699_6);

wire[27:0] addr_700_6;

Selector_2 s700_6(wires_175_5[0], addr_175_5, addr_positional[2803:2800], addr_700_6);

wire[27:0] addr_701_6;

Selector_2 s701_6(wires_175_5[1], addr_175_5, addr_positional[2807:2804], addr_701_6);

wire[27:0] addr_702_6;

Selector_2 s702_6(wires_175_5[2], addr_175_5, addr_positional[2811:2808], addr_702_6);

wire[27:0] addr_703_6;

Selector_2 s703_6(wires_175_5[3], addr_175_5, addr_positional[2815:2812], addr_703_6);

wire[27:0] addr_704_6;

Selector_2 s704_6(wires_176_5[0], addr_176_5, addr_positional[2819:2816], addr_704_6);

wire[27:0] addr_705_6;

Selector_2 s705_6(wires_176_5[1], addr_176_5, addr_positional[2823:2820], addr_705_6);

wire[27:0] addr_706_6;

Selector_2 s706_6(wires_176_5[2], addr_176_5, addr_positional[2827:2824], addr_706_6);

wire[27:0] addr_707_6;

Selector_2 s707_6(wires_176_5[3], addr_176_5, addr_positional[2831:2828], addr_707_6);

wire[27:0] addr_708_6;

Selector_2 s708_6(wires_177_5[0], addr_177_5, addr_positional[2835:2832], addr_708_6);

wire[27:0] addr_709_6;

Selector_2 s709_6(wires_177_5[1], addr_177_5, addr_positional[2839:2836], addr_709_6);

wire[27:0] addr_710_6;

Selector_2 s710_6(wires_177_5[2], addr_177_5, addr_positional[2843:2840], addr_710_6);

wire[27:0] addr_711_6;

Selector_2 s711_6(wires_177_5[3], addr_177_5, addr_positional[2847:2844], addr_711_6);

wire[27:0] addr_712_6;

Selector_2 s712_6(wires_178_5[0], addr_178_5, addr_positional[2851:2848], addr_712_6);

wire[27:0] addr_713_6;

Selector_2 s713_6(wires_178_5[1], addr_178_5, addr_positional[2855:2852], addr_713_6);

wire[27:0] addr_714_6;

Selector_2 s714_6(wires_178_5[2], addr_178_5, addr_positional[2859:2856], addr_714_6);

wire[27:0] addr_715_6;

Selector_2 s715_6(wires_178_5[3], addr_178_5, addr_positional[2863:2860], addr_715_6);

wire[27:0] addr_716_6;

Selector_2 s716_6(wires_179_5[0], addr_179_5, addr_positional[2867:2864], addr_716_6);

wire[27:0] addr_717_6;

Selector_2 s717_6(wires_179_5[1], addr_179_5, addr_positional[2871:2868], addr_717_6);

wire[27:0] addr_718_6;

Selector_2 s718_6(wires_179_5[2], addr_179_5, addr_positional[2875:2872], addr_718_6);

wire[27:0] addr_719_6;

Selector_2 s719_6(wires_179_5[3], addr_179_5, addr_positional[2879:2876], addr_719_6);

wire[27:0] addr_720_6;

Selector_2 s720_6(wires_180_5[0], addr_180_5, addr_positional[2883:2880], addr_720_6);

wire[27:0] addr_721_6;

Selector_2 s721_6(wires_180_5[1], addr_180_5, addr_positional[2887:2884], addr_721_6);

wire[27:0] addr_722_6;

Selector_2 s722_6(wires_180_5[2], addr_180_5, addr_positional[2891:2888], addr_722_6);

wire[27:0] addr_723_6;

Selector_2 s723_6(wires_180_5[3], addr_180_5, addr_positional[2895:2892], addr_723_6);

wire[27:0] addr_724_6;

Selector_2 s724_6(wires_181_5[0], addr_181_5, addr_positional[2899:2896], addr_724_6);

wire[27:0] addr_725_6;

Selector_2 s725_6(wires_181_5[1], addr_181_5, addr_positional[2903:2900], addr_725_6);

wire[27:0] addr_726_6;

Selector_2 s726_6(wires_181_5[2], addr_181_5, addr_positional[2907:2904], addr_726_6);

wire[27:0] addr_727_6;

Selector_2 s727_6(wires_181_5[3], addr_181_5, addr_positional[2911:2908], addr_727_6);

wire[27:0] addr_728_6;

Selector_2 s728_6(wires_182_5[0], addr_182_5, addr_positional[2915:2912], addr_728_6);

wire[27:0] addr_729_6;

Selector_2 s729_6(wires_182_5[1], addr_182_5, addr_positional[2919:2916], addr_729_6);

wire[27:0] addr_730_6;

Selector_2 s730_6(wires_182_5[2], addr_182_5, addr_positional[2923:2920], addr_730_6);

wire[27:0] addr_731_6;

Selector_2 s731_6(wires_182_5[3], addr_182_5, addr_positional[2927:2924], addr_731_6);

wire[27:0] addr_732_6;

Selector_2 s732_6(wires_183_5[0], addr_183_5, addr_positional[2931:2928], addr_732_6);

wire[27:0] addr_733_6;

Selector_2 s733_6(wires_183_5[1], addr_183_5, addr_positional[2935:2932], addr_733_6);

wire[27:0] addr_734_6;

Selector_2 s734_6(wires_183_5[2], addr_183_5, addr_positional[2939:2936], addr_734_6);

wire[27:0] addr_735_6;

Selector_2 s735_6(wires_183_5[3], addr_183_5, addr_positional[2943:2940], addr_735_6);

wire[27:0] addr_736_6;

Selector_2 s736_6(wires_184_5[0], addr_184_5, addr_positional[2947:2944], addr_736_6);

wire[27:0] addr_737_6;

Selector_2 s737_6(wires_184_5[1], addr_184_5, addr_positional[2951:2948], addr_737_6);

wire[27:0] addr_738_6;

Selector_2 s738_6(wires_184_5[2], addr_184_5, addr_positional[2955:2952], addr_738_6);

wire[27:0] addr_739_6;

Selector_2 s739_6(wires_184_5[3], addr_184_5, addr_positional[2959:2956], addr_739_6);

wire[27:0] addr_740_6;

Selector_2 s740_6(wires_185_5[0], addr_185_5, addr_positional[2963:2960], addr_740_6);

wire[27:0] addr_741_6;

Selector_2 s741_6(wires_185_5[1], addr_185_5, addr_positional[2967:2964], addr_741_6);

wire[27:0] addr_742_6;

Selector_2 s742_6(wires_185_5[2], addr_185_5, addr_positional[2971:2968], addr_742_6);

wire[27:0] addr_743_6;

Selector_2 s743_6(wires_185_5[3], addr_185_5, addr_positional[2975:2972], addr_743_6);

wire[27:0] addr_744_6;

Selector_2 s744_6(wires_186_5[0], addr_186_5, addr_positional[2979:2976], addr_744_6);

wire[27:0] addr_745_6;

Selector_2 s745_6(wires_186_5[1], addr_186_5, addr_positional[2983:2980], addr_745_6);

wire[27:0] addr_746_6;

Selector_2 s746_6(wires_186_5[2], addr_186_5, addr_positional[2987:2984], addr_746_6);

wire[27:0] addr_747_6;

Selector_2 s747_6(wires_186_5[3], addr_186_5, addr_positional[2991:2988], addr_747_6);

wire[27:0] addr_748_6;

Selector_2 s748_6(wires_187_5[0], addr_187_5, addr_positional[2995:2992], addr_748_6);

wire[27:0] addr_749_6;

Selector_2 s749_6(wires_187_5[1], addr_187_5, addr_positional[2999:2996], addr_749_6);

wire[27:0] addr_750_6;

Selector_2 s750_6(wires_187_5[2], addr_187_5, addr_positional[3003:3000], addr_750_6);

wire[27:0] addr_751_6;

Selector_2 s751_6(wires_187_5[3], addr_187_5, addr_positional[3007:3004], addr_751_6);

wire[27:0] addr_752_6;

Selector_2 s752_6(wires_188_5[0], addr_188_5, addr_positional[3011:3008], addr_752_6);

wire[27:0] addr_753_6;

Selector_2 s753_6(wires_188_5[1], addr_188_5, addr_positional[3015:3012], addr_753_6);

wire[27:0] addr_754_6;

Selector_2 s754_6(wires_188_5[2], addr_188_5, addr_positional[3019:3016], addr_754_6);

wire[27:0] addr_755_6;

Selector_2 s755_6(wires_188_5[3], addr_188_5, addr_positional[3023:3020], addr_755_6);

wire[27:0] addr_756_6;

Selector_2 s756_6(wires_189_5[0], addr_189_5, addr_positional[3027:3024], addr_756_6);

wire[27:0] addr_757_6;

Selector_2 s757_6(wires_189_5[1], addr_189_5, addr_positional[3031:3028], addr_757_6);

wire[27:0] addr_758_6;

Selector_2 s758_6(wires_189_5[2], addr_189_5, addr_positional[3035:3032], addr_758_6);

wire[27:0] addr_759_6;

Selector_2 s759_6(wires_189_5[3], addr_189_5, addr_positional[3039:3036], addr_759_6);

wire[27:0] addr_760_6;

Selector_2 s760_6(wires_190_5[0], addr_190_5, addr_positional[3043:3040], addr_760_6);

wire[27:0] addr_761_6;

Selector_2 s761_6(wires_190_5[1], addr_190_5, addr_positional[3047:3044], addr_761_6);

wire[27:0] addr_762_6;

Selector_2 s762_6(wires_190_5[2], addr_190_5, addr_positional[3051:3048], addr_762_6);

wire[27:0] addr_763_6;

Selector_2 s763_6(wires_190_5[3], addr_190_5, addr_positional[3055:3052], addr_763_6);

wire[27:0] addr_764_6;

Selector_2 s764_6(wires_191_5[0], addr_191_5, addr_positional[3059:3056], addr_764_6);

wire[27:0] addr_765_6;

Selector_2 s765_6(wires_191_5[1], addr_191_5, addr_positional[3063:3060], addr_765_6);

wire[27:0] addr_766_6;

Selector_2 s766_6(wires_191_5[2], addr_191_5, addr_positional[3067:3064], addr_766_6);

wire[27:0] addr_767_6;

Selector_2 s767_6(wires_191_5[3], addr_191_5, addr_positional[3071:3068], addr_767_6);

wire[27:0] addr_768_6;

Selector_2 s768_6(wires_192_5[0], addr_192_5, addr_positional[3075:3072], addr_768_6);

wire[27:0] addr_769_6;

Selector_2 s769_6(wires_192_5[1], addr_192_5, addr_positional[3079:3076], addr_769_6);

wire[27:0] addr_770_6;

Selector_2 s770_6(wires_192_5[2], addr_192_5, addr_positional[3083:3080], addr_770_6);

wire[27:0] addr_771_6;

Selector_2 s771_6(wires_192_5[3], addr_192_5, addr_positional[3087:3084], addr_771_6);

wire[27:0] addr_772_6;

Selector_2 s772_6(wires_193_5[0], addr_193_5, addr_positional[3091:3088], addr_772_6);

wire[27:0] addr_773_6;

Selector_2 s773_6(wires_193_5[1], addr_193_5, addr_positional[3095:3092], addr_773_6);

wire[27:0] addr_774_6;

Selector_2 s774_6(wires_193_5[2], addr_193_5, addr_positional[3099:3096], addr_774_6);

wire[27:0] addr_775_6;

Selector_2 s775_6(wires_193_5[3], addr_193_5, addr_positional[3103:3100], addr_775_6);

wire[27:0] addr_776_6;

Selector_2 s776_6(wires_194_5[0], addr_194_5, addr_positional[3107:3104], addr_776_6);

wire[27:0] addr_777_6;

Selector_2 s777_6(wires_194_5[1], addr_194_5, addr_positional[3111:3108], addr_777_6);

wire[27:0] addr_778_6;

Selector_2 s778_6(wires_194_5[2], addr_194_5, addr_positional[3115:3112], addr_778_6);

wire[27:0] addr_779_6;

Selector_2 s779_6(wires_194_5[3], addr_194_5, addr_positional[3119:3116], addr_779_6);

wire[27:0] addr_780_6;

Selector_2 s780_6(wires_195_5[0], addr_195_5, addr_positional[3123:3120], addr_780_6);

wire[27:0] addr_781_6;

Selector_2 s781_6(wires_195_5[1], addr_195_5, addr_positional[3127:3124], addr_781_6);

wire[27:0] addr_782_6;

Selector_2 s782_6(wires_195_5[2], addr_195_5, addr_positional[3131:3128], addr_782_6);

wire[27:0] addr_783_6;

Selector_2 s783_6(wires_195_5[3], addr_195_5, addr_positional[3135:3132], addr_783_6);

wire[27:0] addr_784_6;

Selector_2 s784_6(wires_196_5[0], addr_196_5, addr_positional[3139:3136], addr_784_6);

wire[27:0] addr_785_6;

Selector_2 s785_6(wires_196_5[1], addr_196_5, addr_positional[3143:3140], addr_785_6);

wire[27:0] addr_786_6;

Selector_2 s786_6(wires_196_5[2], addr_196_5, addr_positional[3147:3144], addr_786_6);

wire[27:0] addr_787_6;

Selector_2 s787_6(wires_196_5[3], addr_196_5, addr_positional[3151:3148], addr_787_6);

wire[27:0] addr_788_6;

Selector_2 s788_6(wires_197_5[0], addr_197_5, addr_positional[3155:3152], addr_788_6);

wire[27:0] addr_789_6;

Selector_2 s789_6(wires_197_5[1], addr_197_5, addr_positional[3159:3156], addr_789_6);

wire[27:0] addr_790_6;

Selector_2 s790_6(wires_197_5[2], addr_197_5, addr_positional[3163:3160], addr_790_6);

wire[27:0] addr_791_6;

Selector_2 s791_6(wires_197_5[3], addr_197_5, addr_positional[3167:3164], addr_791_6);

wire[27:0] addr_792_6;

Selector_2 s792_6(wires_198_5[0], addr_198_5, addr_positional[3171:3168], addr_792_6);

wire[27:0] addr_793_6;

Selector_2 s793_6(wires_198_5[1], addr_198_5, addr_positional[3175:3172], addr_793_6);

wire[27:0] addr_794_6;

Selector_2 s794_6(wires_198_5[2], addr_198_5, addr_positional[3179:3176], addr_794_6);

wire[27:0] addr_795_6;

Selector_2 s795_6(wires_198_5[3], addr_198_5, addr_positional[3183:3180], addr_795_6);

wire[27:0] addr_796_6;

Selector_2 s796_6(wires_199_5[0], addr_199_5, addr_positional[3187:3184], addr_796_6);

wire[27:0] addr_797_6;

Selector_2 s797_6(wires_199_5[1], addr_199_5, addr_positional[3191:3188], addr_797_6);

wire[27:0] addr_798_6;

Selector_2 s798_6(wires_199_5[2], addr_199_5, addr_positional[3195:3192], addr_798_6);

wire[27:0] addr_799_6;

Selector_2 s799_6(wires_199_5[3], addr_199_5, addr_positional[3199:3196], addr_799_6);

wire[27:0] addr_800_6;

Selector_2 s800_6(wires_200_5[0], addr_200_5, addr_positional[3203:3200], addr_800_6);

wire[27:0] addr_801_6;

Selector_2 s801_6(wires_200_5[1], addr_200_5, addr_positional[3207:3204], addr_801_6);

wire[27:0] addr_802_6;

Selector_2 s802_6(wires_200_5[2], addr_200_5, addr_positional[3211:3208], addr_802_6);

wire[27:0] addr_803_6;

Selector_2 s803_6(wires_200_5[3], addr_200_5, addr_positional[3215:3212], addr_803_6);

wire[27:0] addr_804_6;

Selector_2 s804_6(wires_201_5[0], addr_201_5, addr_positional[3219:3216], addr_804_6);

wire[27:0] addr_805_6;

Selector_2 s805_6(wires_201_5[1], addr_201_5, addr_positional[3223:3220], addr_805_6);

wire[27:0] addr_806_6;

Selector_2 s806_6(wires_201_5[2], addr_201_5, addr_positional[3227:3224], addr_806_6);

wire[27:0] addr_807_6;

Selector_2 s807_6(wires_201_5[3], addr_201_5, addr_positional[3231:3228], addr_807_6);

wire[27:0] addr_808_6;

Selector_2 s808_6(wires_202_5[0], addr_202_5, addr_positional[3235:3232], addr_808_6);

wire[27:0] addr_809_6;

Selector_2 s809_6(wires_202_5[1], addr_202_5, addr_positional[3239:3236], addr_809_6);

wire[27:0] addr_810_6;

Selector_2 s810_6(wires_202_5[2], addr_202_5, addr_positional[3243:3240], addr_810_6);

wire[27:0] addr_811_6;

Selector_2 s811_6(wires_202_5[3], addr_202_5, addr_positional[3247:3244], addr_811_6);

wire[27:0] addr_812_6;

Selector_2 s812_6(wires_203_5[0], addr_203_5, addr_positional[3251:3248], addr_812_6);

wire[27:0] addr_813_6;

Selector_2 s813_6(wires_203_5[1], addr_203_5, addr_positional[3255:3252], addr_813_6);

wire[27:0] addr_814_6;

Selector_2 s814_6(wires_203_5[2], addr_203_5, addr_positional[3259:3256], addr_814_6);

wire[27:0] addr_815_6;

Selector_2 s815_6(wires_203_5[3], addr_203_5, addr_positional[3263:3260], addr_815_6);

wire[27:0] addr_816_6;

Selector_2 s816_6(wires_204_5[0], addr_204_5, addr_positional[3267:3264], addr_816_6);

wire[27:0] addr_817_6;

Selector_2 s817_6(wires_204_5[1], addr_204_5, addr_positional[3271:3268], addr_817_6);

wire[27:0] addr_818_6;

Selector_2 s818_6(wires_204_5[2], addr_204_5, addr_positional[3275:3272], addr_818_6);

wire[27:0] addr_819_6;

Selector_2 s819_6(wires_204_5[3], addr_204_5, addr_positional[3279:3276], addr_819_6);

wire[27:0] addr_820_6;

Selector_2 s820_6(wires_205_5[0], addr_205_5, addr_positional[3283:3280], addr_820_6);

wire[27:0] addr_821_6;

Selector_2 s821_6(wires_205_5[1], addr_205_5, addr_positional[3287:3284], addr_821_6);

wire[27:0] addr_822_6;

Selector_2 s822_6(wires_205_5[2], addr_205_5, addr_positional[3291:3288], addr_822_6);

wire[27:0] addr_823_6;

Selector_2 s823_6(wires_205_5[3], addr_205_5, addr_positional[3295:3292], addr_823_6);

wire[27:0] addr_824_6;

Selector_2 s824_6(wires_206_5[0], addr_206_5, addr_positional[3299:3296], addr_824_6);

wire[27:0] addr_825_6;

Selector_2 s825_6(wires_206_5[1], addr_206_5, addr_positional[3303:3300], addr_825_6);

wire[27:0] addr_826_6;

Selector_2 s826_6(wires_206_5[2], addr_206_5, addr_positional[3307:3304], addr_826_6);

wire[27:0] addr_827_6;

Selector_2 s827_6(wires_206_5[3], addr_206_5, addr_positional[3311:3308], addr_827_6);

wire[27:0] addr_828_6;

Selector_2 s828_6(wires_207_5[0], addr_207_5, addr_positional[3315:3312], addr_828_6);

wire[27:0] addr_829_6;

Selector_2 s829_6(wires_207_5[1], addr_207_5, addr_positional[3319:3316], addr_829_6);

wire[27:0] addr_830_6;

Selector_2 s830_6(wires_207_5[2], addr_207_5, addr_positional[3323:3320], addr_830_6);

wire[27:0] addr_831_6;

Selector_2 s831_6(wires_207_5[3], addr_207_5, addr_positional[3327:3324], addr_831_6);

wire[27:0] addr_832_6;

Selector_2 s832_6(wires_208_5[0], addr_208_5, addr_positional[3331:3328], addr_832_6);

wire[27:0] addr_833_6;

Selector_2 s833_6(wires_208_5[1], addr_208_5, addr_positional[3335:3332], addr_833_6);

wire[27:0] addr_834_6;

Selector_2 s834_6(wires_208_5[2], addr_208_5, addr_positional[3339:3336], addr_834_6);

wire[27:0] addr_835_6;

Selector_2 s835_6(wires_208_5[3], addr_208_5, addr_positional[3343:3340], addr_835_6);

wire[27:0] addr_836_6;

Selector_2 s836_6(wires_209_5[0], addr_209_5, addr_positional[3347:3344], addr_836_6);

wire[27:0] addr_837_6;

Selector_2 s837_6(wires_209_5[1], addr_209_5, addr_positional[3351:3348], addr_837_6);

wire[27:0] addr_838_6;

Selector_2 s838_6(wires_209_5[2], addr_209_5, addr_positional[3355:3352], addr_838_6);

wire[27:0] addr_839_6;

Selector_2 s839_6(wires_209_5[3], addr_209_5, addr_positional[3359:3356], addr_839_6);

wire[27:0] addr_840_6;

Selector_2 s840_6(wires_210_5[0], addr_210_5, addr_positional[3363:3360], addr_840_6);

wire[27:0] addr_841_6;

Selector_2 s841_6(wires_210_5[1], addr_210_5, addr_positional[3367:3364], addr_841_6);

wire[27:0] addr_842_6;

Selector_2 s842_6(wires_210_5[2], addr_210_5, addr_positional[3371:3368], addr_842_6);

wire[27:0] addr_843_6;

Selector_2 s843_6(wires_210_5[3], addr_210_5, addr_positional[3375:3372], addr_843_6);

wire[27:0] addr_844_6;

Selector_2 s844_6(wires_211_5[0], addr_211_5, addr_positional[3379:3376], addr_844_6);

wire[27:0] addr_845_6;

Selector_2 s845_6(wires_211_5[1], addr_211_5, addr_positional[3383:3380], addr_845_6);

wire[27:0] addr_846_6;

Selector_2 s846_6(wires_211_5[2], addr_211_5, addr_positional[3387:3384], addr_846_6);

wire[27:0] addr_847_6;

Selector_2 s847_6(wires_211_5[3], addr_211_5, addr_positional[3391:3388], addr_847_6);

wire[27:0] addr_848_6;

Selector_2 s848_6(wires_212_5[0], addr_212_5, addr_positional[3395:3392], addr_848_6);

wire[27:0] addr_849_6;

Selector_2 s849_6(wires_212_5[1], addr_212_5, addr_positional[3399:3396], addr_849_6);

wire[27:0] addr_850_6;

Selector_2 s850_6(wires_212_5[2], addr_212_5, addr_positional[3403:3400], addr_850_6);

wire[27:0] addr_851_6;

Selector_2 s851_6(wires_212_5[3], addr_212_5, addr_positional[3407:3404], addr_851_6);

wire[27:0] addr_852_6;

Selector_2 s852_6(wires_213_5[0], addr_213_5, addr_positional[3411:3408], addr_852_6);

wire[27:0] addr_853_6;

Selector_2 s853_6(wires_213_5[1], addr_213_5, addr_positional[3415:3412], addr_853_6);

wire[27:0] addr_854_6;

Selector_2 s854_6(wires_213_5[2], addr_213_5, addr_positional[3419:3416], addr_854_6);

wire[27:0] addr_855_6;

Selector_2 s855_6(wires_213_5[3], addr_213_5, addr_positional[3423:3420], addr_855_6);

wire[27:0] addr_856_6;

Selector_2 s856_6(wires_214_5[0], addr_214_5, addr_positional[3427:3424], addr_856_6);

wire[27:0] addr_857_6;

Selector_2 s857_6(wires_214_5[1], addr_214_5, addr_positional[3431:3428], addr_857_6);

wire[27:0] addr_858_6;

Selector_2 s858_6(wires_214_5[2], addr_214_5, addr_positional[3435:3432], addr_858_6);

wire[27:0] addr_859_6;

Selector_2 s859_6(wires_214_5[3], addr_214_5, addr_positional[3439:3436], addr_859_6);

wire[27:0] addr_860_6;

Selector_2 s860_6(wires_215_5[0], addr_215_5, addr_positional[3443:3440], addr_860_6);

wire[27:0] addr_861_6;

Selector_2 s861_6(wires_215_5[1], addr_215_5, addr_positional[3447:3444], addr_861_6);

wire[27:0] addr_862_6;

Selector_2 s862_6(wires_215_5[2], addr_215_5, addr_positional[3451:3448], addr_862_6);

wire[27:0] addr_863_6;

Selector_2 s863_6(wires_215_5[3], addr_215_5, addr_positional[3455:3452], addr_863_6);

wire[27:0] addr_864_6;

Selector_2 s864_6(wires_216_5[0], addr_216_5, addr_positional[3459:3456], addr_864_6);

wire[27:0] addr_865_6;

Selector_2 s865_6(wires_216_5[1], addr_216_5, addr_positional[3463:3460], addr_865_6);

wire[27:0] addr_866_6;

Selector_2 s866_6(wires_216_5[2], addr_216_5, addr_positional[3467:3464], addr_866_6);

wire[27:0] addr_867_6;

Selector_2 s867_6(wires_216_5[3], addr_216_5, addr_positional[3471:3468], addr_867_6);

wire[27:0] addr_868_6;

Selector_2 s868_6(wires_217_5[0], addr_217_5, addr_positional[3475:3472], addr_868_6);

wire[27:0] addr_869_6;

Selector_2 s869_6(wires_217_5[1], addr_217_5, addr_positional[3479:3476], addr_869_6);

wire[27:0] addr_870_6;

Selector_2 s870_6(wires_217_5[2], addr_217_5, addr_positional[3483:3480], addr_870_6);

wire[27:0] addr_871_6;

Selector_2 s871_6(wires_217_5[3], addr_217_5, addr_positional[3487:3484], addr_871_6);

wire[27:0] addr_872_6;

Selector_2 s872_6(wires_218_5[0], addr_218_5, addr_positional[3491:3488], addr_872_6);

wire[27:0] addr_873_6;

Selector_2 s873_6(wires_218_5[1], addr_218_5, addr_positional[3495:3492], addr_873_6);

wire[27:0] addr_874_6;

Selector_2 s874_6(wires_218_5[2], addr_218_5, addr_positional[3499:3496], addr_874_6);

wire[27:0] addr_875_6;

Selector_2 s875_6(wires_218_5[3], addr_218_5, addr_positional[3503:3500], addr_875_6);

wire[27:0] addr_876_6;

Selector_2 s876_6(wires_219_5[0], addr_219_5, addr_positional[3507:3504], addr_876_6);

wire[27:0] addr_877_6;

Selector_2 s877_6(wires_219_5[1], addr_219_5, addr_positional[3511:3508], addr_877_6);

wire[27:0] addr_878_6;

Selector_2 s878_6(wires_219_5[2], addr_219_5, addr_positional[3515:3512], addr_878_6);

wire[27:0] addr_879_6;

Selector_2 s879_6(wires_219_5[3], addr_219_5, addr_positional[3519:3516], addr_879_6);

wire[27:0] addr_880_6;

Selector_2 s880_6(wires_220_5[0], addr_220_5, addr_positional[3523:3520], addr_880_6);

wire[27:0] addr_881_6;

Selector_2 s881_6(wires_220_5[1], addr_220_5, addr_positional[3527:3524], addr_881_6);

wire[27:0] addr_882_6;

Selector_2 s882_6(wires_220_5[2], addr_220_5, addr_positional[3531:3528], addr_882_6);

wire[27:0] addr_883_6;

Selector_2 s883_6(wires_220_5[3], addr_220_5, addr_positional[3535:3532], addr_883_6);

wire[27:0] addr_884_6;

Selector_2 s884_6(wires_221_5[0], addr_221_5, addr_positional[3539:3536], addr_884_6);

wire[27:0] addr_885_6;

Selector_2 s885_6(wires_221_5[1], addr_221_5, addr_positional[3543:3540], addr_885_6);

wire[27:0] addr_886_6;

Selector_2 s886_6(wires_221_5[2], addr_221_5, addr_positional[3547:3544], addr_886_6);

wire[27:0] addr_887_6;

Selector_2 s887_6(wires_221_5[3], addr_221_5, addr_positional[3551:3548], addr_887_6);

wire[27:0] addr_888_6;

Selector_2 s888_6(wires_222_5[0], addr_222_5, addr_positional[3555:3552], addr_888_6);

wire[27:0] addr_889_6;

Selector_2 s889_6(wires_222_5[1], addr_222_5, addr_positional[3559:3556], addr_889_6);

wire[27:0] addr_890_6;

Selector_2 s890_6(wires_222_5[2], addr_222_5, addr_positional[3563:3560], addr_890_6);

wire[27:0] addr_891_6;

Selector_2 s891_6(wires_222_5[3], addr_222_5, addr_positional[3567:3564], addr_891_6);

wire[27:0] addr_892_6;

Selector_2 s892_6(wires_223_5[0], addr_223_5, addr_positional[3571:3568], addr_892_6);

wire[27:0] addr_893_6;

Selector_2 s893_6(wires_223_5[1], addr_223_5, addr_positional[3575:3572], addr_893_6);

wire[27:0] addr_894_6;

Selector_2 s894_6(wires_223_5[2], addr_223_5, addr_positional[3579:3576], addr_894_6);

wire[27:0] addr_895_6;

Selector_2 s895_6(wires_223_5[3], addr_223_5, addr_positional[3583:3580], addr_895_6);

wire[27:0] addr_896_6;

Selector_2 s896_6(wires_224_5[0], addr_224_5, addr_positional[3587:3584], addr_896_6);

wire[27:0] addr_897_6;

Selector_2 s897_6(wires_224_5[1], addr_224_5, addr_positional[3591:3588], addr_897_6);

wire[27:0] addr_898_6;

Selector_2 s898_6(wires_224_5[2], addr_224_5, addr_positional[3595:3592], addr_898_6);

wire[27:0] addr_899_6;

Selector_2 s899_6(wires_224_5[3], addr_224_5, addr_positional[3599:3596], addr_899_6);

wire[27:0] addr_900_6;

Selector_2 s900_6(wires_225_5[0], addr_225_5, addr_positional[3603:3600], addr_900_6);

wire[27:0] addr_901_6;

Selector_2 s901_6(wires_225_5[1], addr_225_5, addr_positional[3607:3604], addr_901_6);

wire[27:0] addr_902_6;

Selector_2 s902_6(wires_225_5[2], addr_225_5, addr_positional[3611:3608], addr_902_6);

wire[27:0] addr_903_6;

Selector_2 s903_6(wires_225_5[3], addr_225_5, addr_positional[3615:3612], addr_903_6);

wire[27:0] addr_904_6;

Selector_2 s904_6(wires_226_5[0], addr_226_5, addr_positional[3619:3616], addr_904_6);

wire[27:0] addr_905_6;

Selector_2 s905_6(wires_226_5[1], addr_226_5, addr_positional[3623:3620], addr_905_6);

wire[27:0] addr_906_6;

Selector_2 s906_6(wires_226_5[2], addr_226_5, addr_positional[3627:3624], addr_906_6);

wire[27:0] addr_907_6;

Selector_2 s907_6(wires_226_5[3], addr_226_5, addr_positional[3631:3628], addr_907_6);

wire[27:0] addr_908_6;

Selector_2 s908_6(wires_227_5[0], addr_227_5, addr_positional[3635:3632], addr_908_6);

wire[27:0] addr_909_6;

Selector_2 s909_6(wires_227_5[1], addr_227_5, addr_positional[3639:3636], addr_909_6);

wire[27:0] addr_910_6;

Selector_2 s910_6(wires_227_5[2], addr_227_5, addr_positional[3643:3640], addr_910_6);

wire[27:0] addr_911_6;

Selector_2 s911_6(wires_227_5[3], addr_227_5, addr_positional[3647:3644], addr_911_6);

wire[27:0] addr_912_6;

Selector_2 s912_6(wires_228_5[0], addr_228_5, addr_positional[3651:3648], addr_912_6);

wire[27:0] addr_913_6;

Selector_2 s913_6(wires_228_5[1], addr_228_5, addr_positional[3655:3652], addr_913_6);

wire[27:0] addr_914_6;

Selector_2 s914_6(wires_228_5[2], addr_228_5, addr_positional[3659:3656], addr_914_6);

wire[27:0] addr_915_6;

Selector_2 s915_6(wires_228_5[3], addr_228_5, addr_positional[3663:3660], addr_915_6);

wire[27:0] addr_916_6;

Selector_2 s916_6(wires_229_5[0], addr_229_5, addr_positional[3667:3664], addr_916_6);

wire[27:0] addr_917_6;

Selector_2 s917_6(wires_229_5[1], addr_229_5, addr_positional[3671:3668], addr_917_6);

wire[27:0] addr_918_6;

Selector_2 s918_6(wires_229_5[2], addr_229_5, addr_positional[3675:3672], addr_918_6);

wire[27:0] addr_919_6;

Selector_2 s919_6(wires_229_5[3], addr_229_5, addr_positional[3679:3676], addr_919_6);

wire[27:0] addr_920_6;

Selector_2 s920_6(wires_230_5[0], addr_230_5, addr_positional[3683:3680], addr_920_6);

wire[27:0] addr_921_6;

Selector_2 s921_6(wires_230_5[1], addr_230_5, addr_positional[3687:3684], addr_921_6);

wire[27:0] addr_922_6;

Selector_2 s922_6(wires_230_5[2], addr_230_5, addr_positional[3691:3688], addr_922_6);

wire[27:0] addr_923_6;

Selector_2 s923_6(wires_230_5[3], addr_230_5, addr_positional[3695:3692], addr_923_6);

wire[27:0] addr_924_6;

Selector_2 s924_6(wires_231_5[0], addr_231_5, addr_positional[3699:3696], addr_924_6);

wire[27:0] addr_925_6;

Selector_2 s925_6(wires_231_5[1], addr_231_5, addr_positional[3703:3700], addr_925_6);

wire[27:0] addr_926_6;

Selector_2 s926_6(wires_231_5[2], addr_231_5, addr_positional[3707:3704], addr_926_6);

wire[27:0] addr_927_6;

Selector_2 s927_6(wires_231_5[3], addr_231_5, addr_positional[3711:3708], addr_927_6);

wire[27:0] addr_928_6;

Selector_2 s928_6(wires_232_5[0], addr_232_5, addr_positional[3715:3712], addr_928_6);

wire[27:0] addr_929_6;

Selector_2 s929_6(wires_232_5[1], addr_232_5, addr_positional[3719:3716], addr_929_6);

wire[27:0] addr_930_6;

Selector_2 s930_6(wires_232_5[2], addr_232_5, addr_positional[3723:3720], addr_930_6);

wire[27:0] addr_931_6;

Selector_2 s931_6(wires_232_5[3], addr_232_5, addr_positional[3727:3724], addr_931_6);

wire[27:0] addr_932_6;

Selector_2 s932_6(wires_233_5[0], addr_233_5, addr_positional[3731:3728], addr_932_6);

wire[27:0] addr_933_6;

Selector_2 s933_6(wires_233_5[1], addr_233_5, addr_positional[3735:3732], addr_933_6);

wire[27:0] addr_934_6;

Selector_2 s934_6(wires_233_5[2], addr_233_5, addr_positional[3739:3736], addr_934_6);

wire[27:0] addr_935_6;

Selector_2 s935_6(wires_233_5[3], addr_233_5, addr_positional[3743:3740], addr_935_6);

wire[27:0] addr_936_6;

Selector_2 s936_6(wires_234_5[0], addr_234_5, addr_positional[3747:3744], addr_936_6);

wire[27:0] addr_937_6;

Selector_2 s937_6(wires_234_5[1], addr_234_5, addr_positional[3751:3748], addr_937_6);

wire[27:0] addr_938_6;

Selector_2 s938_6(wires_234_5[2], addr_234_5, addr_positional[3755:3752], addr_938_6);

wire[27:0] addr_939_6;

Selector_2 s939_6(wires_234_5[3], addr_234_5, addr_positional[3759:3756], addr_939_6);

wire[27:0] addr_940_6;

Selector_2 s940_6(wires_235_5[0], addr_235_5, addr_positional[3763:3760], addr_940_6);

wire[27:0] addr_941_6;

Selector_2 s941_6(wires_235_5[1], addr_235_5, addr_positional[3767:3764], addr_941_6);

wire[27:0] addr_942_6;

Selector_2 s942_6(wires_235_5[2], addr_235_5, addr_positional[3771:3768], addr_942_6);

wire[27:0] addr_943_6;

Selector_2 s943_6(wires_235_5[3], addr_235_5, addr_positional[3775:3772], addr_943_6);

wire[27:0] addr_944_6;

Selector_2 s944_6(wires_236_5[0], addr_236_5, addr_positional[3779:3776], addr_944_6);

wire[27:0] addr_945_6;

Selector_2 s945_6(wires_236_5[1], addr_236_5, addr_positional[3783:3780], addr_945_6);

wire[27:0] addr_946_6;

Selector_2 s946_6(wires_236_5[2], addr_236_5, addr_positional[3787:3784], addr_946_6);

wire[27:0] addr_947_6;

Selector_2 s947_6(wires_236_5[3], addr_236_5, addr_positional[3791:3788], addr_947_6);

wire[27:0] addr_948_6;

Selector_2 s948_6(wires_237_5[0], addr_237_5, addr_positional[3795:3792], addr_948_6);

wire[27:0] addr_949_6;

Selector_2 s949_6(wires_237_5[1], addr_237_5, addr_positional[3799:3796], addr_949_6);

wire[27:0] addr_950_6;

Selector_2 s950_6(wires_237_5[2], addr_237_5, addr_positional[3803:3800], addr_950_6);

wire[27:0] addr_951_6;

Selector_2 s951_6(wires_237_5[3], addr_237_5, addr_positional[3807:3804], addr_951_6);

wire[27:0] addr_952_6;

Selector_2 s952_6(wires_238_5[0], addr_238_5, addr_positional[3811:3808], addr_952_6);

wire[27:0] addr_953_6;

Selector_2 s953_6(wires_238_5[1], addr_238_5, addr_positional[3815:3812], addr_953_6);

wire[27:0] addr_954_6;

Selector_2 s954_6(wires_238_5[2], addr_238_5, addr_positional[3819:3816], addr_954_6);

wire[27:0] addr_955_6;

Selector_2 s955_6(wires_238_5[3], addr_238_5, addr_positional[3823:3820], addr_955_6);

wire[27:0] addr_956_6;

Selector_2 s956_6(wires_239_5[0], addr_239_5, addr_positional[3827:3824], addr_956_6);

wire[27:0] addr_957_6;

Selector_2 s957_6(wires_239_5[1], addr_239_5, addr_positional[3831:3828], addr_957_6);

wire[27:0] addr_958_6;

Selector_2 s958_6(wires_239_5[2], addr_239_5, addr_positional[3835:3832], addr_958_6);

wire[27:0] addr_959_6;

Selector_2 s959_6(wires_239_5[3], addr_239_5, addr_positional[3839:3836], addr_959_6);

wire[27:0] addr_960_6;

Selector_2 s960_6(wires_240_5[0], addr_240_5, addr_positional[3843:3840], addr_960_6);

wire[27:0] addr_961_6;

Selector_2 s961_6(wires_240_5[1], addr_240_5, addr_positional[3847:3844], addr_961_6);

wire[27:0] addr_962_6;

Selector_2 s962_6(wires_240_5[2], addr_240_5, addr_positional[3851:3848], addr_962_6);

wire[27:0] addr_963_6;

Selector_2 s963_6(wires_240_5[3], addr_240_5, addr_positional[3855:3852], addr_963_6);

wire[27:0] addr_964_6;

Selector_2 s964_6(wires_241_5[0], addr_241_5, addr_positional[3859:3856], addr_964_6);

wire[27:0] addr_965_6;

Selector_2 s965_6(wires_241_5[1], addr_241_5, addr_positional[3863:3860], addr_965_6);

wire[27:0] addr_966_6;

Selector_2 s966_6(wires_241_5[2], addr_241_5, addr_positional[3867:3864], addr_966_6);

wire[27:0] addr_967_6;

Selector_2 s967_6(wires_241_5[3], addr_241_5, addr_positional[3871:3868], addr_967_6);

wire[27:0] addr_968_6;

Selector_2 s968_6(wires_242_5[0], addr_242_5, addr_positional[3875:3872], addr_968_6);

wire[27:0] addr_969_6;

Selector_2 s969_6(wires_242_5[1], addr_242_5, addr_positional[3879:3876], addr_969_6);

wire[27:0] addr_970_6;

Selector_2 s970_6(wires_242_5[2], addr_242_5, addr_positional[3883:3880], addr_970_6);

wire[27:0] addr_971_6;

Selector_2 s971_6(wires_242_5[3], addr_242_5, addr_positional[3887:3884], addr_971_6);

wire[27:0] addr_972_6;

Selector_2 s972_6(wires_243_5[0], addr_243_5, addr_positional[3891:3888], addr_972_6);

wire[27:0] addr_973_6;

Selector_2 s973_6(wires_243_5[1], addr_243_5, addr_positional[3895:3892], addr_973_6);

wire[27:0] addr_974_6;

Selector_2 s974_6(wires_243_5[2], addr_243_5, addr_positional[3899:3896], addr_974_6);

wire[27:0] addr_975_6;

Selector_2 s975_6(wires_243_5[3], addr_243_5, addr_positional[3903:3900], addr_975_6);

wire[27:0] addr_976_6;

Selector_2 s976_6(wires_244_5[0], addr_244_5, addr_positional[3907:3904], addr_976_6);

wire[27:0] addr_977_6;

Selector_2 s977_6(wires_244_5[1], addr_244_5, addr_positional[3911:3908], addr_977_6);

wire[27:0] addr_978_6;

Selector_2 s978_6(wires_244_5[2], addr_244_5, addr_positional[3915:3912], addr_978_6);

wire[27:0] addr_979_6;

Selector_2 s979_6(wires_244_5[3], addr_244_5, addr_positional[3919:3916], addr_979_6);

wire[27:0] addr_980_6;

Selector_2 s980_6(wires_245_5[0], addr_245_5, addr_positional[3923:3920], addr_980_6);

wire[27:0] addr_981_6;

Selector_2 s981_6(wires_245_5[1], addr_245_5, addr_positional[3927:3924], addr_981_6);

wire[27:0] addr_982_6;

Selector_2 s982_6(wires_245_5[2], addr_245_5, addr_positional[3931:3928], addr_982_6);

wire[27:0] addr_983_6;

Selector_2 s983_6(wires_245_5[3], addr_245_5, addr_positional[3935:3932], addr_983_6);

wire[27:0] addr_984_6;

Selector_2 s984_6(wires_246_5[0], addr_246_5, addr_positional[3939:3936], addr_984_6);

wire[27:0] addr_985_6;

Selector_2 s985_6(wires_246_5[1], addr_246_5, addr_positional[3943:3940], addr_985_6);

wire[27:0] addr_986_6;

Selector_2 s986_6(wires_246_5[2], addr_246_5, addr_positional[3947:3944], addr_986_6);

wire[27:0] addr_987_6;

Selector_2 s987_6(wires_246_5[3], addr_246_5, addr_positional[3951:3948], addr_987_6);

wire[27:0] addr_988_6;

Selector_2 s988_6(wires_247_5[0], addr_247_5, addr_positional[3955:3952], addr_988_6);

wire[27:0] addr_989_6;

Selector_2 s989_6(wires_247_5[1], addr_247_5, addr_positional[3959:3956], addr_989_6);

wire[27:0] addr_990_6;

Selector_2 s990_6(wires_247_5[2], addr_247_5, addr_positional[3963:3960], addr_990_6);

wire[27:0] addr_991_6;

Selector_2 s991_6(wires_247_5[3], addr_247_5, addr_positional[3967:3964], addr_991_6);

wire[27:0] addr_992_6;

Selector_2 s992_6(wires_248_5[0], addr_248_5, addr_positional[3971:3968], addr_992_6);

wire[27:0] addr_993_6;

Selector_2 s993_6(wires_248_5[1], addr_248_5, addr_positional[3975:3972], addr_993_6);

wire[27:0] addr_994_6;

Selector_2 s994_6(wires_248_5[2], addr_248_5, addr_positional[3979:3976], addr_994_6);

wire[27:0] addr_995_6;

Selector_2 s995_6(wires_248_5[3], addr_248_5, addr_positional[3983:3980], addr_995_6);

wire[27:0] addr_996_6;

Selector_2 s996_6(wires_249_5[0], addr_249_5, addr_positional[3987:3984], addr_996_6);

wire[27:0] addr_997_6;

Selector_2 s997_6(wires_249_5[1], addr_249_5, addr_positional[3991:3988], addr_997_6);

wire[27:0] addr_998_6;

Selector_2 s998_6(wires_249_5[2], addr_249_5, addr_positional[3995:3992], addr_998_6);

wire[27:0] addr_999_6;

Selector_2 s999_6(wires_249_5[3], addr_249_5, addr_positional[3999:3996], addr_999_6);

wire[27:0] addr_1000_6;

Selector_2 s1000_6(wires_250_5[0], addr_250_5, addr_positional[4003:4000], addr_1000_6);

wire[27:0] addr_1001_6;

Selector_2 s1001_6(wires_250_5[1], addr_250_5, addr_positional[4007:4004], addr_1001_6);

wire[27:0] addr_1002_6;

Selector_2 s1002_6(wires_250_5[2], addr_250_5, addr_positional[4011:4008], addr_1002_6);

wire[27:0] addr_1003_6;

Selector_2 s1003_6(wires_250_5[3], addr_250_5, addr_positional[4015:4012], addr_1003_6);

wire[27:0] addr_1004_6;

Selector_2 s1004_6(wires_251_5[0], addr_251_5, addr_positional[4019:4016], addr_1004_6);

wire[27:0] addr_1005_6;

Selector_2 s1005_6(wires_251_5[1], addr_251_5, addr_positional[4023:4020], addr_1005_6);

wire[27:0] addr_1006_6;

Selector_2 s1006_6(wires_251_5[2], addr_251_5, addr_positional[4027:4024], addr_1006_6);

wire[27:0] addr_1007_6;

Selector_2 s1007_6(wires_251_5[3], addr_251_5, addr_positional[4031:4028], addr_1007_6);

wire[27:0] addr_1008_6;

Selector_2 s1008_6(wires_252_5[0], addr_252_5, addr_positional[4035:4032], addr_1008_6);

wire[27:0] addr_1009_6;

Selector_2 s1009_6(wires_252_5[1], addr_252_5, addr_positional[4039:4036], addr_1009_6);

wire[27:0] addr_1010_6;

Selector_2 s1010_6(wires_252_5[2], addr_252_5, addr_positional[4043:4040], addr_1010_6);

wire[27:0] addr_1011_6;

Selector_2 s1011_6(wires_252_5[3], addr_252_5, addr_positional[4047:4044], addr_1011_6);

wire[27:0] addr_1012_6;

Selector_2 s1012_6(wires_253_5[0], addr_253_5, addr_positional[4051:4048], addr_1012_6);

wire[27:0] addr_1013_6;

Selector_2 s1013_6(wires_253_5[1], addr_253_5, addr_positional[4055:4052], addr_1013_6);

wire[27:0] addr_1014_6;

Selector_2 s1014_6(wires_253_5[2], addr_253_5, addr_positional[4059:4056], addr_1014_6);

wire[27:0] addr_1015_6;

Selector_2 s1015_6(wires_253_5[3], addr_253_5, addr_positional[4063:4060], addr_1015_6);

wire[27:0] addr_1016_6;

Selector_2 s1016_6(wires_254_5[0], addr_254_5, addr_positional[4067:4064], addr_1016_6);

wire[27:0] addr_1017_6;

Selector_2 s1017_6(wires_254_5[1], addr_254_5, addr_positional[4071:4068], addr_1017_6);

wire[27:0] addr_1018_6;

Selector_2 s1018_6(wires_254_5[2], addr_254_5, addr_positional[4075:4072], addr_1018_6);

wire[27:0] addr_1019_6;

Selector_2 s1019_6(wires_254_5[3], addr_254_5, addr_positional[4079:4076], addr_1019_6);

wire[27:0] addr_1020_6;

Selector_2 s1020_6(wires_255_5[0], addr_255_5, addr_positional[4083:4080], addr_1020_6);

wire[27:0] addr_1021_6;

Selector_2 s1021_6(wires_255_5[1], addr_255_5, addr_positional[4087:4084], addr_1021_6);

wire[27:0] addr_1022_6;

Selector_2 s1022_6(wires_255_5[2], addr_255_5, addr_positional[4091:4088], addr_1022_6);

wire[27:0] addr_1023_6;

Selector_2 s1023_6(wires_255_5[3], addr_255_5, addr_positional[4095:4092], addr_1023_6);

wire[27:0] addr_1024_6;

Selector_2 s1024_6(wires_256_5[0], addr_256_5, addr_positional[4099:4096], addr_1024_6);

wire[27:0] addr_1025_6;

Selector_2 s1025_6(wires_256_5[1], addr_256_5, addr_positional[4103:4100], addr_1025_6);

wire[27:0] addr_1026_6;

Selector_2 s1026_6(wires_256_5[2], addr_256_5, addr_positional[4107:4104], addr_1026_6);

wire[27:0] addr_1027_6;

Selector_2 s1027_6(wires_256_5[3], addr_256_5, addr_positional[4111:4108], addr_1027_6);

wire[27:0] addr_1028_6;

Selector_2 s1028_6(wires_257_5[0], addr_257_5, addr_positional[4115:4112], addr_1028_6);

wire[27:0] addr_1029_6;

Selector_2 s1029_6(wires_257_5[1], addr_257_5, addr_positional[4119:4116], addr_1029_6);

wire[27:0] addr_1030_6;

Selector_2 s1030_6(wires_257_5[2], addr_257_5, addr_positional[4123:4120], addr_1030_6);

wire[27:0] addr_1031_6;

Selector_2 s1031_6(wires_257_5[3], addr_257_5, addr_positional[4127:4124], addr_1031_6);

wire[27:0] addr_1032_6;

Selector_2 s1032_6(wires_258_5[0], addr_258_5, addr_positional[4131:4128], addr_1032_6);

wire[27:0] addr_1033_6;

Selector_2 s1033_6(wires_258_5[1], addr_258_5, addr_positional[4135:4132], addr_1033_6);

wire[27:0] addr_1034_6;

Selector_2 s1034_6(wires_258_5[2], addr_258_5, addr_positional[4139:4136], addr_1034_6);

wire[27:0] addr_1035_6;

Selector_2 s1035_6(wires_258_5[3], addr_258_5, addr_positional[4143:4140], addr_1035_6);

wire[27:0] addr_1036_6;

Selector_2 s1036_6(wires_259_5[0], addr_259_5, addr_positional[4147:4144], addr_1036_6);

wire[27:0] addr_1037_6;

Selector_2 s1037_6(wires_259_5[1], addr_259_5, addr_positional[4151:4148], addr_1037_6);

wire[27:0] addr_1038_6;

Selector_2 s1038_6(wires_259_5[2], addr_259_5, addr_positional[4155:4152], addr_1038_6);

wire[27:0] addr_1039_6;

Selector_2 s1039_6(wires_259_5[3], addr_259_5, addr_positional[4159:4156], addr_1039_6);

wire[27:0] addr_1040_6;

Selector_2 s1040_6(wires_260_5[0], addr_260_5, addr_positional[4163:4160], addr_1040_6);

wire[27:0] addr_1041_6;

Selector_2 s1041_6(wires_260_5[1], addr_260_5, addr_positional[4167:4164], addr_1041_6);

wire[27:0] addr_1042_6;

Selector_2 s1042_6(wires_260_5[2], addr_260_5, addr_positional[4171:4168], addr_1042_6);

wire[27:0] addr_1043_6;

Selector_2 s1043_6(wires_260_5[3], addr_260_5, addr_positional[4175:4172], addr_1043_6);

wire[27:0] addr_1044_6;

Selector_2 s1044_6(wires_261_5[0], addr_261_5, addr_positional[4179:4176], addr_1044_6);

wire[27:0] addr_1045_6;

Selector_2 s1045_6(wires_261_5[1], addr_261_5, addr_positional[4183:4180], addr_1045_6);

wire[27:0] addr_1046_6;

Selector_2 s1046_6(wires_261_5[2], addr_261_5, addr_positional[4187:4184], addr_1046_6);

wire[27:0] addr_1047_6;

Selector_2 s1047_6(wires_261_5[3], addr_261_5, addr_positional[4191:4188], addr_1047_6);

wire[27:0] addr_1048_6;

Selector_2 s1048_6(wires_262_5[0], addr_262_5, addr_positional[4195:4192], addr_1048_6);

wire[27:0] addr_1049_6;

Selector_2 s1049_6(wires_262_5[1], addr_262_5, addr_positional[4199:4196], addr_1049_6);

wire[27:0] addr_1050_6;

Selector_2 s1050_6(wires_262_5[2], addr_262_5, addr_positional[4203:4200], addr_1050_6);

wire[27:0] addr_1051_6;

Selector_2 s1051_6(wires_262_5[3], addr_262_5, addr_positional[4207:4204], addr_1051_6);

wire[27:0] addr_1052_6;

Selector_2 s1052_6(wires_263_5[0], addr_263_5, addr_positional[4211:4208], addr_1052_6);

wire[27:0] addr_1053_6;

Selector_2 s1053_6(wires_263_5[1], addr_263_5, addr_positional[4215:4212], addr_1053_6);

wire[27:0] addr_1054_6;

Selector_2 s1054_6(wires_263_5[2], addr_263_5, addr_positional[4219:4216], addr_1054_6);

wire[27:0] addr_1055_6;

Selector_2 s1055_6(wires_263_5[3], addr_263_5, addr_positional[4223:4220], addr_1055_6);

wire[27:0] addr_1056_6;

Selector_2 s1056_6(wires_264_5[0], addr_264_5, addr_positional[4227:4224], addr_1056_6);

wire[27:0] addr_1057_6;

Selector_2 s1057_6(wires_264_5[1], addr_264_5, addr_positional[4231:4228], addr_1057_6);

wire[27:0] addr_1058_6;

Selector_2 s1058_6(wires_264_5[2], addr_264_5, addr_positional[4235:4232], addr_1058_6);

wire[27:0] addr_1059_6;

Selector_2 s1059_6(wires_264_5[3], addr_264_5, addr_positional[4239:4236], addr_1059_6);

wire[27:0] addr_1060_6;

Selector_2 s1060_6(wires_265_5[0], addr_265_5, addr_positional[4243:4240], addr_1060_6);

wire[27:0] addr_1061_6;

Selector_2 s1061_6(wires_265_5[1], addr_265_5, addr_positional[4247:4244], addr_1061_6);

wire[27:0] addr_1062_6;

Selector_2 s1062_6(wires_265_5[2], addr_265_5, addr_positional[4251:4248], addr_1062_6);

wire[27:0] addr_1063_6;

Selector_2 s1063_6(wires_265_5[3], addr_265_5, addr_positional[4255:4252], addr_1063_6);

wire[27:0] addr_1064_6;

Selector_2 s1064_6(wires_266_5[0], addr_266_5, addr_positional[4259:4256], addr_1064_6);

wire[27:0] addr_1065_6;

Selector_2 s1065_6(wires_266_5[1], addr_266_5, addr_positional[4263:4260], addr_1065_6);

wire[27:0] addr_1066_6;

Selector_2 s1066_6(wires_266_5[2], addr_266_5, addr_positional[4267:4264], addr_1066_6);

wire[27:0] addr_1067_6;

Selector_2 s1067_6(wires_266_5[3], addr_266_5, addr_positional[4271:4268], addr_1067_6);

wire[27:0] addr_1068_6;

Selector_2 s1068_6(wires_267_5[0], addr_267_5, addr_positional[4275:4272], addr_1068_6);

wire[27:0] addr_1069_6;

Selector_2 s1069_6(wires_267_5[1], addr_267_5, addr_positional[4279:4276], addr_1069_6);

wire[27:0] addr_1070_6;

Selector_2 s1070_6(wires_267_5[2], addr_267_5, addr_positional[4283:4280], addr_1070_6);

wire[27:0] addr_1071_6;

Selector_2 s1071_6(wires_267_5[3], addr_267_5, addr_positional[4287:4284], addr_1071_6);

wire[27:0] addr_1072_6;

Selector_2 s1072_6(wires_268_5[0], addr_268_5, addr_positional[4291:4288], addr_1072_6);

wire[27:0] addr_1073_6;

Selector_2 s1073_6(wires_268_5[1], addr_268_5, addr_positional[4295:4292], addr_1073_6);

wire[27:0] addr_1074_6;

Selector_2 s1074_6(wires_268_5[2], addr_268_5, addr_positional[4299:4296], addr_1074_6);

wire[27:0] addr_1075_6;

Selector_2 s1075_6(wires_268_5[3], addr_268_5, addr_positional[4303:4300], addr_1075_6);

wire[27:0] addr_1076_6;

Selector_2 s1076_6(wires_269_5[0], addr_269_5, addr_positional[4307:4304], addr_1076_6);

wire[27:0] addr_1077_6;

Selector_2 s1077_6(wires_269_5[1], addr_269_5, addr_positional[4311:4308], addr_1077_6);

wire[27:0] addr_1078_6;

Selector_2 s1078_6(wires_269_5[2], addr_269_5, addr_positional[4315:4312], addr_1078_6);

wire[27:0] addr_1079_6;

Selector_2 s1079_6(wires_269_5[3], addr_269_5, addr_positional[4319:4316], addr_1079_6);

wire[27:0] addr_1080_6;

Selector_2 s1080_6(wires_270_5[0], addr_270_5, addr_positional[4323:4320], addr_1080_6);

wire[27:0] addr_1081_6;

Selector_2 s1081_6(wires_270_5[1], addr_270_5, addr_positional[4327:4324], addr_1081_6);

wire[27:0] addr_1082_6;

Selector_2 s1082_6(wires_270_5[2], addr_270_5, addr_positional[4331:4328], addr_1082_6);

wire[27:0] addr_1083_6;

Selector_2 s1083_6(wires_270_5[3], addr_270_5, addr_positional[4335:4332], addr_1083_6);

wire[27:0] addr_1084_6;

Selector_2 s1084_6(wires_271_5[0], addr_271_5, addr_positional[4339:4336], addr_1084_6);

wire[27:0] addr_1085_6;

Selector_2 s1085_6(wires_271_5[1], addr_271_5, addr_positional[4343:4340], addr_1085_6);

wire[27:0] addr_1086_6;

Selector_2 s1086_6(wires_271_5[2], addr_271_5, addr_positional[4347:4344], addr_1086_6);

wire[27:0] addr_1087_6;

Selector_2 s1087_6(wires_271_5[3], addr_271_5, addr_positional[4351:4348], addr_1087_6);

wire[27:0] addr_1088_6;

Selector_2 s1088_6(wires_272_5[0], addr_272_5, addr_positional[4355:4352], addr_1088_6);

wire[27:0] addr_1089_6;

Selector_2 s1089_6(wires_272_5[1], addr_272_5, addr_positional[4359:4356], addr_1089_6);

wire[27:0] addr_1090_6;

Selector_2 s1090_6(wires_272_5[2], addr_272_5, addr_positional[4363:4360], addr_1090_6);

wire[27:0] addr_1091_6;

Selector_2 s1091_6(wires_272_5[3], addr_272_5, addr_positional[4367:4364], addr_1091_6);

wire[27:0] addr_1092_6;

Selector_2 s1092_6(wires_273_5[0], addr_273_5, addr_positional[4371:4368], addr_1092_6);

wire[27:0] addr_1093_6;

Selector_2 s1093_6(wires_273_5[1], addr_273_5, addr_positional[4375:4372], addr_1093_6);

wire[27:0] addr_1094_6;

Selector_2 s1094_6(wires_273_5[2], addr_273_5, addr_positional[4379:4376], addr_1094_6);

wire[27:0] addr_1095_6;

Selector_2 s1095_6(wires_273_5[3], addr_273_5, addr_positional[4383:4380], addr_1095_6);

wire[27:0] addr_1096_6;

Selector_2 s1096_6(wires_274_5[0], addr_274_5, addr_positional[4387:4384], addr_1096_6);

wire[27:0] addr_1097_6;

Selector_2 s1097_6(wires_274_5[1], addr_274_5, addr_positional[4391:4388], addr_1097_6);

wire[27:0] addr_1098_6;

Selector_2 s1098_6(wires_274_5[2], addr_274_5, addr_positional[4395:4392], addr_1098_6);

wire[27:0] addr_1099_6;

Selector_2 s1099_6(wires_274_5[3], addr_274_5, addr_positional[4399:4396], addr_1099_6);

wire[27:0] addr_1100_6;

Selector_2 s1100_6(wires_275_5[0], addr_275_5, addr_positional[4403:4400], addr_1100_6);

wire[27:0] addr_1101_6;

Selector_2 s1101_6(wires_275_5[1], addr_275_5, addr_positional[4407:4404], addr_1101_6);

wire[27:0] addr_1102_6;

Selector_2 s1102_6(wires_275_5[2], addr_275_5, addr_positional[4411:4408], addr_1102_6);

wire[27:0] addr_1103_6;

Selector_2 s1103_6(wires_275_5[3], addr_275_5, addr_positional[4415:4412], addr_1103_6);

wire[27:0] addr_1104_6;

Selector_2 s1104_6(wires_276_5[0], addr_276_5, addr_positional[4419:4416], addr_1104_6);

wire[27:0] addr_1105_6;

Selector_2 s1105_6(wires_276_5[1], addr_276_5, addr_positional[4423:4420], addr_1105_6);

wire[27:0] addr_1106_6;

Selector_2 s1106_6(wires_276_5[2], addr_276_5, addr_positional[4427:4424], addr_1106_6);

wire[27:0] addr_1107_6;

Selector_2 s1107_6(wires_276_5[3], addr_276_5, addr_positional[4431:4428], addr_1107_6);

wire[27:0] addr_1108_6;

Selector_2 s1108_6(wires_277_5[0], addr_277_5, addr_positional[4435:4432], addr_1108_6);

wire[27:0] addr_1109_6;

Selector_2 s1109_6(wires_277_5[1], addr_277_5, addr_positional[4439:4436], addr_1109_6);

wire[27:0] addr_1110_6;

Selector_2 s1110_6(wires_277_5[2], addr_277_5, addr_positional[4443:4440], addr_1110_6);

wire[27:0] addr_1111_6;

Selector_2 s1111_6(wires_277_5[3], addr_277_5, addr_positional[4447:4444], addr_1111_6);

wire[27:0] addr_1112_6;

Selector_2 s1112_6(wires_278_5[0], addr_278_5, addr_positional[4451:4448], addr_1112_6);

wire[27:0] addr_1113_6;

Selector_2 s1113_6(wires_278_5[1], addr_278_5, addr_positional[4455:4452], addr_1113_6);

wire[27:0] addr_1114_6;

Selector_2 s1114_6(wires_278_5[2], addr_278_5, addr_positional[4459:4456], addr_1114_6);

wire[27:0] addr_1115_6;

Selector_2 s1115_6(wires_278_5[3], addr_278_5, addr_positional[4463:4460], addr_1115_6);

wire[27:0] addr_1116_6;

Selector_2 s1116_6(wires_279_5[0], addr_279_5, addr_positional[4467:4464], addr_1116_6);

wire[27:0] addr_1117_6;

Selector_2 s1117_6(wires_279_5[1], addr_279_5, addr_positional[4471:4468], addr_1117_6);

wire[27:0] addr_1118_6;

Selector_2 s1118_6(wires_279_5[2], addr_279_5, addr_positional[4475:4472], addr_1118_6);

wire[27:0] addr_1119_6;

Selector_2 s1119_6(wires_279_5[3], addr_279_5, addr_positional[4479:4476], addr_1119_6);

wire[27:0] addr_1120_6;

Selector_2 s1120_6(wires_280_5[0], addr_280_5, addr_positional[4483:4480], addr_1120_6);

wire[27:0] addr_1121_6;

Selector_2 s1121_6(wires_280_5[1], addr_280_5, addr_positional[4487:4484], addr_1121_6);

wire[27:0] addr_1122_6;

Selector_2 s1122_6(wires_280_5[2], addr_280_5, addr_positional[4491:4488], addr_1122_6);

wire[27:0] addr_1123_6;

Selector_2 s1123_6(wires_280_5[3], addr_280_5, addr_positional[4495:4492], addr_1123_6);

wire[27:0] addr_1124_6;

Selector_2 s1124_6(wires_281_5[0], addr_281_5, addr_positional[4499:4496], addr_1124_6);

wire[27:0] addr_1125_6;

Selector_2 s1125_6(wires_281_5[1], addr_281_5, addr_positional[4503:4500], addr_1125_6);

wire[27:0] addr_1126_6;

Selector_2 s1126_6(wires_281_5[2], addr_281_5, addr_positional[4507:4504], addr_1126_6);

wire[27:0] addr_1127_6;

Selector_2 s1127_6(wires_281_5[3], addr_281_5, addr_positional[4511:4508], addr_1127_6);

wire[27:0] addr_1128_6;

Selector_2 s1128_6(wires_282_5[0], addr_282_5, addr_positional[4515:4512], addr_1128_6);

wire[27:0] addr_1129_6;

Selector_2 s1129_6(wires_282_5[1], addr_282_5, addr_positional[4519:4516], addr_1129_6);

wire[27:0] addr_1130_6;

Selector_2 s1130_6(wires_282_5[2], addr_282_5, addr_positional[4523:4520], addr_1130_6);

wire[27:0] addr_1131_6;

Selector_2 s1131_6(wires_282_5[3], addr_282_5, addr_positional[4527:4524], addr_1131_6);

wire[27:0] addr_1132_6;

Selector_2 s1132_6(wires_283_5[0], addr_283_5, addr_positional[4531:4528], addr_1132_6);

wire[27:0] addr_1133_6;

Selector_2 s1133_6(wires_283_5[1], addr_283_5, addr_positional[4535:4532], addr_1133_6);

wire[27:0] addr_1134_6;

Selector_2 s1134_6(wires_283_5[2], addr_283_5, addr_positional[4539:4536], addr_1134_6);

wire[27:0] addr_1135_6;

Selector_2 s1135_6(wires_283_5[3], addr_283_5, addr_positional[4543:4540], addr_1135_6);

wire[27:0] addr_1136_6;

Selector_2 s1136_6(wires_284_5[0], addr_284_5, addr_positional[4547:4544], addr_1136_6);

wire[27:0] addr_1137_6;

Selector_2 s1137_6(wires_284_5[1], addr_284_5, addr_positional[4551:4548], addr_1137_6);

wire[27:0] addr_1138_6;

Selector_2 s1138_6(wires_284_5[2], addr_284_5, addr_positional[4555:4552], addr_1138_6);

wire[27:0] addr_1139_6;

Selector_2 s1139_6(wires_284_5[3], addr_284_5, addr_positional[4559:4556], addr_1139_6);

wire[27:0] addr_1140_6;

Selector_2 s1140_6(wires_285_5[0], addr_285_5, addr_positional[4563:4560], addr_1140_6);

wire[27:0] addr_1141_6;

Selector_2 s1141_6(wires_285_5[1], addr_285_5, addr_positional[4567:4564], addr_1141_6);

wire[27:0] addr_1142_6;

Selector_2 s1142_6(wires_285_5[2], addr_285_5, addr_positional[4571:4568], addr_1142_6);

wire[27:0] addr_1143_6;

Selector_2 s1143_6(wires_285_5[3], addr_285_5, addr_positional[4575:4572], addr_1143_6);

wire[27:0] addr_1144_6;

Selector_2 s1144_6(wires_286_5[0], addr_286_5, addr_positional[4579:4576], addr_1144_6);

wire[27:0] addr_1145_6;

Selector_2 s1145_6(wires_286_5[1], addr_286_5, addr_positional[4583:4580], addr_1145_6);

wire[27:0] addr_1146_6;

Selector_2 s1146_6(wires_286_5[2], addr_286_5, addr_positional[4587:4584], addr_1146_6);

wire[27:0] addr_1147_6;

Selector_2 s1147_6(wires_286_5[3], addr_286_5, addr_positional[4591:4588], addr_1147_6);

wire[27:0] addr_1148_6;

Selector_2 s1148_6(wires_287_5[0], addr_287_5, addr_positional[4595:4592], addr_1148_6);

wire[27:0] addr_1149_6;

Selector_2 s1149_6(wires_287_5[1], addr_287_5, addr_positional[4599:4596], addr_1149_6);

wire[27:0] addr_1150_6;

Selector_2 s1150_6(wires_287_5[2], addr_287_5, addr_positional[4603:4600], addr_1150_6);

wire[27:0] addr_1151_6;

Selector_2 s1151_6(wires_287_5[3], addr_287_5, addr_positional[4607:4604], addr_1151_6);

wire[27:0] addr_1152_6;

Selector_2 s1152_6(wires_288_5[0], addr_288_5, addr_positional[4611:4608], addr_1152_6);

wire[27:0] addr_1153_6;

Selector_2 s1153_6(wires_288_5[1], addr_288_5, addr_positional[4615:4612], addr_1153_6);

wire[27:0] addr_1154_6;

Selector_2 s1154_6(wires_288_5[2], addr_288_5, addr_positional[4619:4616], addr_1154_6);

wire[27:0] addr_1155_6;

Selector_2 s1155_6(wires_288_5[3], addr_288_5, addr_positional[4623:4620], addr_1155_6);

wire[27:0] addr_1156_6;

Selector_2 s1156_6(wires_289_5[0], addr_289_5, addr_positional[4627:4624], addr_1156_6);

wire[27:0] addr_1157_6;

Selector_2 s1157_6(wires_289_5[1], addr_289_5, addr_positional[4631:4628], addr_1157_6);

wire[27:0] addr_1158_6;

Selector_2 s1158_6(wires_289_5[2], addr_289_5, addr_positional[4635:4632], addr_1158_6);

wire[27:0] addr_1159_6;

Selector_2 s1159_6(wires_289_5[3], addr_289_5, addr_positional[4639:4636], addr_1159_6);

wire[27:0] addr_1160_6;

Selector_2 s1160_6(wires_290_5[0], addr_290_5, addr_positional[4643:4640], addr_1160_6);

wire[27:0] addr_1161_6;

Selector_2 s1161_6(wires_290_5[1], addr_290_5, addr_positional[4647:4644], addr_1161_6);

wire[27:0] addr_1162_6;

Selector_2 s1162_6(wires_290_5[2], addr_290_5, addr_positional[4651:4648], addr_1162_6);

wire[27:0] addr_1163_6;

Selector_2 s1163_6(wires_290_5[3], addr_290_5, addr_positional[4655:4652], addr_1163_6);

wire[27:0] addr_1164_6;

Selector_2 s1164_6(wires_291_5[0], addr_291_5, addr_positional[4659:4656], addr_1164_6);

wire[27:0] addr_1165_6;

Selector_2 s1165_6(wires_291_5[1], addr_291_5, addr_positional[4663:4660], addr_1165_6);

wire[27:0] addr_1166_6;

Selector_2 s1166_6(wires_291_5[2], addr_291_5, addr_positional[4667:4664], addr_1166_6);

wire[27:0] addr_1167_6;

Selector_2 s1167_6(wires_291_5[3], addr_291_5, addr_positional[4671:4668], addr_1167_6);

wire[27:0] addr_1168_6;

Selector_2 s1168_6(wires_292_5[0], addr_292_5, addr_positional[4675:4672], addr_1168_6);

wire[27:0] addr_1169_6;

Selector_2 s1169_6(wires_292_5[1], addr_292_5, addr_positional[4679:4676], addr_1169_6);

wire[27:0] addr_1170_6;

Selector_2 s1170_6(wires_292_5[2], addr_292_5, addr_positional[4683:4680], addr_1170_6);

wire[27:0] addr_1171_6;

Selector_2 s1171_6(wires_292_5[3], addr_292_5, addr_positional[4687:4684], addr_1171_6);

wire[27:0] addr_1172_6;

Selector_2 s1172_6(wires_293_5[0], addr_293_5, addr_positional[4691:4688], addr_1172_6);

wire[27:0] addr_1173_6;

Selector_2 s1173_6(wires_293_5[1], addr_293_5, addr_positional[4695:4692], addr_1173_6);

wire[27:0] addr_1174_6;

Selector_2 s1174_6(wires_293_5[2], addr_293_5, addr_positional[4699:4696], addr_1174_6);

wire[27:0] addr_1175_6;

Selector_2 s1175_6(wires_293_5[3], addr_293_5, addr_positional[4703:4700], addr_1175_6);

wire[27:0] addr_1176_6;

Selector_2 s1176_6(wires_294_5[0], addr_294_5, addr_positional[4707:4704], addr_1176_6);

wire[27:0] addr_1177_6;

Selector_2 s1177_6(wires_294_5[1], addr_294_5, addr_positional[4711:4708], addr_1177_6);

wire[27:0] addr_1178_6;

Selector_2 s1178_6(wires_294_5[2], addr_294_5, addr_positional[4715:4712], addr_1178_6);

wire[27:0] addr_1179_6;

Selector_2 s1179_6(wires_294_5[3], addr_294_5, addr_positional[4719:4716], addr_1179_6);

wire[27:0] addr_1180_6;

Selector_2 s1180_6(wires_295_5[0], addr_295_5, addr_positional[4723:4720], addr_1180_6);

wire[27:0] addr_1181_6;

Selector_2 s1181_6(wires_295_5[1], addr_295_5, addr_positional[4727:4724], addr_1181_6);

wire[27:0] addr_1182_6;

Selector_2 s1182_6(wires_295_5[2], addr_295_5, addr_positional[4731:4728], addr_1182_6);

wire[27:0] addr_1183_6;

Selector_2 s1183_6(wires_295_5[3], addr_295_5, addr_positional[4735:4732], addr_1183_6);

wire[27:0] addr_1184_6;

Selector_2 s1184_6(wires_296_5[0], addr_296_5, addr_positional[4739:4736], addr_1184_6);

wire[27:0] addr_1185_6;

Selector_2 s1185_6(wires_296_5[1], addr_296_5, addr_positional[4743:4740], addr_1185_6);

wire[27:0] addr_1186_6;

Selector_2 s1186_6(wires_296_5[2], addr_296_5, addr_positional[4747:4744], addr_1186_6);

wire[27:0] addr_1187_6;

Selector_2 s1187_6(wires_296_5[3], addr_296_5, addr_positional[4751:4748], addr_1187_6);

wire[27:0] addr_1188_6;

Selector_2 s1188_6(wires_297_5[0], addr_297_5, addr_positional[4755:4752], addr_1188_6);

wire[27:0] addr_1189_6;

Selector_2 s1189_6(wires_297_5[1], addr_297_5, addr_positional[4759:4756], addr_1189_6);

wire[27:0] addr_1190_6;

Selector_2 s1190_6(wires_297_5[2], addr_297_5, addr_positional[4763:4760], addr_1190_6);

wire[27:0] addr_1191_6;

Selector_2 s1191_6(wires_297_5[3], addr_297_5, addr_positional[4767:4764], addr_1191_6);

wire[27:0] addr_1192_6;

Selector_2 s1192_6(wires_298_5[0], addr_298_5, addr_positional[4771:4768], addr_1192_6);

wire[27:0] addr_1193_6;

Selector_2 s1193_6(wires_298_5[1], addr_298_5, addr_positional[4775:4772], addr_1193_6);

wire[27:0] addr_1194_6;

Selector_2 s1194_6(wires_298_5[2], addr_298_5, addr_positional[4779:4776], addr_1194_6);

wire[27:0] addr_1195_6;

Selector_2 s1195_6(wires_298_5[3], addr_298_5, addr_positional[4783:4780], addr_1195_6);

wire[27:0] addr_1196_6;

Selector_2 s1196_6(wires_299_5[0], addr_299_5, addr_positional[4787:4784], addr_1196_6);

wire[27:0] addr_1197_6;

Selector_2 s1197_6(wires_299_5[1], addr_299_5, addr_positional[4791:4788], addr_1197_6);

wire[27:0] addr_1198_6;

Selector_2 s1198_6(wires_299_5[2], addr_299_5, addr_positional[4795:4792], addr_1198_6);

wire[27:0] addr_1199_6;

Selector_2 s1199_6(wires_299_5[3], addr_299_5, addr_positional[4799:4796], addr_1199_6);

wire[27:0] addr_1200_6;

Selector_2 s1200_6(wires_300_5[0], addr_300_5, addr_positional[4803:4800], addr_1200_6);

wire[27:0] addr_1201_6;

Selector_2 s1201_6(wires_300_5[1], addr_300_5, addr_positional[4807:4804], addr_1201_6);

wire[27:0] addr_1202_6;

Selector_2 s1202_6(wires_300_5[2], addr_300_5, addr_positional[4811:4808], addr_1202_6);

wire[27:0] addr_1203_6;

Selector_2 s1203_6(wires_300_5[3], addr_300_5, addr_positional[4815:4812], addr_1203_6);

wire[27:0] addr_1204_6;

Selector_2 s1204_6(wires_301_5[0], addr_301_5, addr_positional[4819:4816], addr_1204_6);

wire[27:0] addr_1205_6;

Selector_2 s1205_6(wires_301_5[1], addr_301_5, addr_positional[4823:4820], addr_1205_6);

wire[27:0] addr_1206_6;

Selector_2 s1206_6(wires_301_5[2], addr_301_5, addr_positional[4827:4824], addr_1206_6);

wire[27:0] addr_1207_6;

Selector_2 s1207_6(wires_301_5[3], addr_301_5, addr_positional[4831:4828], addr_1207_6);

wire[27:0] addr_1208_6;

Selector_2 s1208_6(wires_302_5[0], addr_302_5, addr_positional[4835:4832], addr_1208_6);

wire[27:0] addr_1209_6;

Selector_2 s1209_6(wires_302_5[1], addr_302_5, addr_positional[4839:4836], addr_1209_6);

wire[27:0] addr_1210_6;

Selector_2 s1210_6(wires_302_5[2], addr_302_5, addr_positional[4843:4840], addr_1210_6);

wire[27:0] addr_1211_6;

Selector_2 s1211_6(wires_302_5[3], addr_302_5, addr_positional[4847:4844], addr_1211_6);

wire[27:0] addr_1212_6;

Selector_2 s1212_6(wires_303_5[0], addr_303_5, addr_positional[4851:4848], addr_1212_6);

wire[27:0] addr_1213_6;

Selector_2 s1213_6(wires_303_5[1], addr_303_5, addr_positional[4855:4852], addr_1213_6);

wire[27:0] addr_1214_6;

Selector_2 s1214_6(wires_303_5[2], addr_303_5, addr_positional[4859:4856], addr_1214_6);

wire[27:0] addr_1215_6;

Selector_2 s1215_6(wires_303_5[3], addr_303_5, addr_positional[4863:4860], addr_1215_6);

wire[27:0] addr_1216_6;

Selector_2 s1216_6(wires_304_5[0], addr_304_5, addr_positional[4867:4864], addr_1216_6);

wire[27:0] addr_1217_6;

Selector_2 s1217_6(wires_304_5[1], addr_304_5, addr_positional[4871:4868], addr_1217_6);

wire[27:0] addr_1218_6;

Selector_2 s1218_6(wires_304_5[2], addr_304_5, addr_positional[4875:4872], addr_1218_6);

wire[27:0] addr_1219_6;

Selector_2 s1219_6(wires_304_5[3], addr_304_5, addr_positional[4879:4876], addr_1219_6);

wire[27:0] addr_1220_6;

Selector_2 s1220_6(wires_305_5[0], addr_305_5, addr_positional[4883:4880], addr_1220_6);

wire[27:0] addr_1221_6;

Selector_2 s1221_6(wires_305_5[1], addr_305_5, addr_positional[4887:4884], addr_1221_6);

wire[27:0] addr_1222_6;

Selector_2 s1222_6(wires_305_5[2], addr_305_5, addr_positional[4891:4888], addr_1222_6);

wire[27:0] addr_1223_6;

Selector_2 s1223_6(wires_305_5[3], addr_305_5, addr_positional[4895:4892], addr_1223_6);

wire[27:0] addr_1224_6;

Selector_2 s1224_6(wires_306_5[0], addr_306_5, addr_positional[4899:4896], addr_1224_6);

wire[27:0] addr_1225_6;

Selector_2 s1225_6(wires_306_5[1], addr_306_5, addr_positional[4903:4900], addr_1225_6);

wire[27:0] addr_1226_6;

Selector_2 s1226_6(wires_306_5[2], addr_306_5, addr_positional[4907:4904], addr_1226_6);

wire[27:0] addr_1227_6;

Selector_2 s1227_6(wires_306_5[3], addr_306_5, addr_positional[4911:4908], addr_1227_6);

wire[27:0] addr_1228_6;

Selector_2 s1228_6(wires_307_5[0], addr_307_5, addr_positional[4915:4912], addr_1228_6);

wire[27:0] addr_1229_6;

Selector_2 s1229_6(wires_307_5[1], addr_307_5, addr_positional[4919:4916], addr_1229_6);

wire[27:0] addr_1230_6;

Selector_2 s1230_6(wires_307_5[2], addr_307_5, addr_positional[4923:4920], addr_1230_6);

wire[27:0] addr_1231_6;

Selector_2 s1231_6(wires_307_5[3], addr_307_5, addr_positional[4927:4924], addr_1231_6);

wire[27:0] addr_1232_6;

Selector_2 s1232_6(wires_308_5[0], addr_308_5, addr_positional[4931:4928], addr_1232_6);

wire[27:0] addr_1233_6;

Selector_2 s1233_6(wires_308_5[1], addr_308_5, addr_positional[4935:4932], addr_1233_6);

wire[27:0] addr_1234_6;

Selector_2 s1234_6(wires_308_5[2], addr_308_5, addr_positional[4939:4936], addr_1234_6);

wire[27:0] addr_1235_6;

Selector_2 s1235_6(wires_308_5[3], addr_308_5, addr_positional[4943:4940], addr_1235_6);

wire[27:0] addr_1236_6;

Selector_2 s1236_6(wires_309_5[0], addr_309_5, addr_positional[4947:4944], addr_1236_6);

wire[27:0] addr_1237_6;

Selector_2 s1237_6(wires_309_5[1], addr_309_5, addr_positional[4951:4948], addr_1237_6);

wire[27:0] addr_1238_6;

Selector_2 s1238_6(wires_309_5[2], addr_309_5, addr_positional[4955:4952], addr_1238_6);

wire[27:0] addr_1239_6;

Selector_2 s1239_6(wires_309_5[3], addr_309_5, addr_positional[4959:4956], addr_1239_6);

wire[27:0] addr_1240_6;

Selector_2 s1240_6(wires_310_5[0], addr_310_5, addr_positional[4963:4960], addr_1240_6);

wire[27:0] addr_1241_6;

Selector_2 s1241_6(wires_310_5[1], addr_310_5, addr_positional[4967:4964], addr_1241_6);

wire[27:0] addr_1242_6;

Selector_2 s1242_6(wires_310_5[2], addr_310_5, addr_positional[4971:4968], addr_1242_6);

wire[27:0] addr_1243_6;

Selector_2 s1243_6(wires_310_5[3], addr_310_5, addr_positional[4975:4972], addr_1243_6);

wire[27:0] addr_1244_6;

Selector_2 s1244_6(wires_311_5[0], addr_311_5, addr_positional[4979:4976], addr_1244_6);

wire[27:0] addr_1245_6;

Selector_2 s1245_6(wires_311_5[1], addr_311_5, addr_positional[4983:4980], addr_1245_6);

wire[27:0] addr_1246_6;

Selector_2 s1246_6(wires_311_5[2], addr_311_5, addr_positional[4987:4984], addr_1246_6);

wire[27:0] addr_1247_6;

Selector_2 s1247_6(wires_311_5[3], addr_311_5, addr_positional[4991:4988], addr_1247_6);

wire[27:0] addr_1248_6;

Selector_2 s1248_6(wires_312_5[0], addr_312_5, addr_positional[4995:4992], addr_1248_6);

wire[27:0] addr_1249_6;

Selector_2 s1249_6(wires_312_5[1], addr_312_5, addr_positional[4999:4996], addr_1249_6);

wire[27:0] addr_1250_6;

Selector_2 s1250_6(wires_312_5[2], addr_312_5, addr_positional[5003:5000], addr_1250_6);

wire[27:0] addr_1251_6;

Selector_2 s1251_6(wires_312_5[3], addr_312_5, addr_positional[5007:5004], addr_1251_6);

wire[27:0] addr_1252_6;

Selector_2 s1252_6(wires_313_5[0], addr_313_5, addr_positional[5011:5008], addr_1252_6);

wire[27:0] addr_1253_6;

Selector_2 s1253_6(wires_313_5[1], addr_313_5, addr_positional[5015:5012], addr_1253_6);

wire[27:0] addr_1254_6;

Selector_2 s1254_6(wires_313_5[2], addr_313_5, addr_positional[5019:5016], addr_1254_6);

wire[27:0] addr_1255_6;

Selector_2 s1255_6(wires_313_5[3], addr_313_5, addr_positional[5023:5020], addr_1255_6);

wire[27:0] addr_1256_6;

Selector_2 s1256_6(wires_314_5[0], addr_314_5, addr_positional[5027:5024], addr_1256_6);

wire[27:0] addr_1257_6;

Selector_2 s1257_6(wires_314_5[1], addr_314_5, addr_positional[5031:5028], addr_1257_6);

wire[27:0] addr_1258_6;

Selector_2 s1258_6(wires_314_5[2], addr_314_5, addr_positional[5035:5032], addr_1258_6);

wire[27:0] addr_1259_6;

Selector_2 s1259_6(wires_314_5[3], addr_314_5, addr_positional[5039:5036], addr_1259_6);

wire[27:0] addr_1260_6;

Selector_2 s1260_6(wires_315_5[0], addr_315_5, addr_positional[5043:5040], addr_1260_6);

wire[27:0] addr_1261_6;

Selector_2 s1261_6(wires_315_5[1], addr_315_5, addr_positional[5047:5044], addr_1261_6);

wire[27:0] addr_1262_6;

Selector_2 s1262_6(wires_315_5[2], addr_315_5, addr_positional[5051:5048], addr_1262_6);

wire[27:0] addr_1263_6;

Selector_2 s1263_6(wires_315_5[3], addr_315_5, addr_positional[5055:5052], addr_1263_6);

wire[27:0] addr_1264_6;

Selector_2 s1264_6(wires_316_5[0], addr_316_5, addr_positional[5059:5056], addr_1264_6);

wire[27:0] addr_1265_6;

Selector_2 s1265_6(wires_316_5[1], addr_316_5, addr_positional[5063:5060], addr_1265_6);

wire[27:0] addr_1266_6;

Selector_2 s1266_6(wires_316_5[2], addr_316_5, addr_positional[5067:5064], addr_1266_6);

wire[27:0] addr_1267_6;

Selector_2 s1267_6(wires_316_5[3], addr_316_5, addr_positional[5071:5068], addr_1267_6);

wire[27:0] addr_1268_6;

Selector_2 s1268_6(wires_317_5[0], addr_317_5, addr_positional[5075:5072], addr_1268_6);

wire[27:0] addr_1269_6;

Selector_2 s1269_6(wires_317_5[1], addr_317_5, addr_positional[5079:5076], addr_1269_6);

wire[27:0] addr_1270_6;

Selector_2 s1270_6(wires_317_5[2], addr_317_5, addr_positional[5083:5080], addr_1270_6);

wire[27:0] addr_1271_6;

Selector_2 s1271_6(wires_317_5[3], addr_317_5, addr_positional[5087:5084], addr_1271_6);

wire[27:0] addr_1272_6;

Selector_2 s1272_6(wires_318_5[0], addr_318_5, addr_positional[5091:5088], addr_1272_6);

wire[27:0] addr_1273_6;

Selector_2 s1273_6(wires_318_5[1], addr_318_5, addr_positional[5095:5092], addr_1273_6);

wire[27:0] addr_1274_6;

Selector_2 s1274_6(wires_318_5[2], addr_318_5, addr_positional[5099:5096], addr_1274_6);

wire[27:0] addr_1275_6;

Selector_2 s1275_6(wires_318_5[3], addr_318_5, addr_positional[5103:5100], addr_1275_6);

wire[27:0] addr_1276_6;

Selector_2 s1276_6(wires_319_5[0], addr_319_5, addr_positional[5107:5104], addr_1276_6);

wire[27:0] addr_1277_6;

Selector_2 s1277_6(wires_319_5[1], addr_319_5, addr_positional[5111:5108], addr_1277_6);

wire[27:0] addr_1278_6;

Selector_2 s1278_6(wires_319_5[2], addr_319_5, addr_positional[5115:5112], addr_1278_6);

wire[27:0] addr_1279_6;

Selector_2 s1279_6(wires_319_5[3], addr_319_5, addr_positional[5119:5116], addr_1279_6);

wire[27:0] addr_1280_6;

Selector_2 s1280_6(wires_320_5[0], addr_320_5, addr_positional[5123:5120], addr_1280_6);

wire[27:0] addr_1281_6;

Selector_2 s1281_6(wires_320_5[1], addr_320_5, addr_positional[5127:5124], addr_1281_6);

wire[27:0] addr_1282_6;

Selector_2 s1282_6(wires_320_5[2], addr_320_5, addr_positional[5131:5128], addr_1282_6);

wire[27:0] addr_1283_6;

Selector_2 s1283_6(wires_320_5[3], addr_320_5, addr_positional[5135:5132], addr_1283_6);

wire[27:0] addr_1284_6;

Selector_2 s1284_6(wires_321_5[0], addr_321_5, addr_positional[5139:5136], addr_1284_6);

wire[27:0] addr_1285_6;

Selector_2 s1285_6(wires_321_5[1], addr_321_5, addr_positional[5143:5140], addr_1285_6);

wire[27:0] addr_1286_6;

Selector_2 s1286_6(wires_321_5[2], addr_321_5, addr_positional[5147:5144], addr_1286_6);

wire[27:0] addr_1287_6;

Selector_2 s1287_6(wires_321_5[3], addr_321_5, addr_positional[5151:5148], addr_1287_6);

wire[27:0] addr_1288_6;

Selector_2 s1288_6(wires_322_5[0], addr_322_5, addr_positional[5155:5152], addr_1288_6);

wire[27:0] addr_1289_6;

Selector_2 s1289_6(wires_322_5[1], addr_322_5, addr_positional[5159:5156], addr_1289_6);

wire[27:0] addr_1290_6;

Selector_2 s1290_6(wires_322_5[2], addr_322_5, addr_positional[5163:5160], addr_1290_6);

wire[27:0] addr_1291_6;

Selector_2 s1291_6(wires_322_5[3], addr_322_5, addr_positional[5167:5164], addr_1291_6);

wire[27:0] addr_1292_6;

Selector_2 s1292_6(wires_323_5[0], addr_323_5, addr_positional[5171:5168], addr_1292_6);

wire[27:0] addr_1293_6;

Selector_2 s1293_6(wires_323_5[1], addr_323_5, addr_positional[5175:5172], addr_1293_6);

wire[27:0] addr_1294_6;

Selector_2 s1294_6(wires_323_5[2], addr_323_5, addr_positional[5179:5176], addr_1294_6);

wire[27:0] addr_1295_6;

Selector_2 s1295_6(wires_323_5[3], addr_323_5, addr_positional[5183:5180], addr_1295_6);

wire[27:0] addr_1296_6;

Selector_2 s1296_6(wires_324_5[0], addr_324_5, addr_positional[5187:5184], addr_1296_6);

wire[27:0] addr_1297_6;

Selector_2 s1297_6(wires_324_5[1], addr_324_5, addr_positional[5191:5188], addr_1297_6);

wire[27:0] addr_1298_6;

Selector_2 s1298_6(wires_324_5[2], addr_324_5, addr_positional[5195:5192], addr_1298_6);

wire[27:0] addr_1299_6;

Selector_2 s1299_6(wires_324_5[3], addr_324_5, addr_positional[5199:5196], addr_1299_6);

wire[27:0] addr_1300_6;

Selector_2 s1300_6(wires_325_5[0], addr_325_5, addr_positional[5203:5200], addr_1300_6);

wire[27:0] addr_1301_6;

Selector_2 s1301_6(wires_325_5[1], addr_325_5, addr_positional[5207:5204], addr_1301_6);

wire[27:0] addr_1302_6;

Selector_2 s1302_6(wires_325_5[2], addr_325_5, addr_positional[5211:5208], addr_1302_6);

wire[27:0] addr_1303_6;

Selector_2 s1303_6(wires_325_5[3], addr_325_5, addr_positional[5215:5212], addr_1303_6);

wire[27:0] addr_1304_6;

Selector_2 s1304_6(wires_326_5[0], addr_326_5, addr_positional[5219:5216], addr_1304_6);

wire[27:0] addr_1305_6;

Selector_2 s1305_6(wires_326_5[1], addr_326_5, addr_positional[5223:5220], addr_1305_6);

wire[27:0] addr_1306_6;

Selector_2 s1306_6(wires_326_5[2], addr_326_5, addr_positional[5227:5224], addr_1306_6);

wire[27:0] addr_1307_6;

Selector_2 s1307_6(wires_326_5[3], addr_326_5, addr_positional[5231:5228], addr_1307_6);

wire[27:0] addr_1308_6;

Selector_2 s1308_6(wires_327_5[0], addr_327_5, addr_positional[5235:5232], addr_1308_6);

wire[27:0] addr_1309_6;

Selector_2 s1309_6(wires_327_5[1], addr_327_5, addr_positional[5239:5236], addr_1309_6);

wire[27:0] addr_1310_6;

Selector_2 s1310_6(wires_327_5[2], addr_327_5, addr_positional[5243:5240], addr_1310_6);

wire[27:0] addr_1311_6;

Selector_2 s1311_6(wires_327_5[3], addr_327_5, addr_positional[5247:5244], addr_1311_6);

wire[27:0] addr_1312_6;

Selector_2 s1312_6(wires_328_5[0], addr_328_5, addr_positional[5251:5248], addr_1312_6);

wire[27:0] addr_1313_6;

Selector_2 s1313_6(wires_328_5[1], addr_328_5, addr_positional[5255:5252], addr_1313_6);

wire[27:0] addr_1314_6;

Selector_2 s1314_6(wires_328_5[2], addr_328_5, addr_positional[5259:5256], addr_1314_6);

wire[27:0] addr_1315_6;

Selector_2 s1315_6(wires_328_5[3], addr_328_5, addr_positional[5263:5260], addr_1315_6);

wire[27:0] addr_1316_6;

Selector_2 s1316_6(wires_329_5[0], addr_329_5, addr_positional[5267:5264], addr_1316_6);

wire[27:0] addr_1317_6;

Selector_2 s1317_6(wires_329_5[1], addr_329_5, addr_positional[5271:5268], addr_1317_6);

wire[27:0] addr_1318_6;

Selector_2 s1318_6(wires_329_5[2], addr_329_5, addr_positional[5275:5272], addr_1318_6);

wire[27:0] addr_1319_6;

Selector_2 s1319_6(wires_329_5[3], addr_329_5, addr_positional[5279:5276], addr_1319_6);

wire[27:0] addr_1320_6;

Selector_2 s1320_6(wires_330_5[0], addr_330_5, addr_positional[5283:5280], addr_1320_6);

wire[27:0] addr_1321_6;

Selector_2 s1321_6(wires_330_5[1], addr_330_5, addr_positional[5287:5284], addr_1321_6);

wire[27:0] addr_1322_6;

Selector_2 s1322_6(wires_330_5[2], addr_330_5, addr_positional[5291:5288], addr_1322_6);

wire[27:0] addr_1323_6;

Selector_2 s1323_6(wires_330_5[3], addr_330_5, addr_positional[5295:5292], addr_1323_6);

wire[27:0] addr_1324_6;

Selector_2 s1324_6(wires_331_5[0], addr_331_5, addr_positional[5299:5296], addr_1324_6);

wire[27:0] addr_1325_6;

Selector_2 s1325_6(wires_331_5[1], addr_331_5, addr_positional[5303:5300], addr_1325_6);

wire[27:0] addr_1326_6;

Selector_2 s1326_6(wires_331_5[2], addr_331_5, addr_positional[5307:5304], addr_1326_6);

wire[27:0] addr_1327_6;

Selector_2 s1327_6(wires_331_5[3], addr_331_5, addr_positional[5311:5308], addr_1327_6);

wire[27:0] addr_1328_6;

Selector_2 s1328_6(wires_332_5[0], addr_332_5, addr_positional[5315:5312], addr_1328_6);

wire[27:0] addr_1329_6;

Selector_2 s1329_6(wires_332_5[1], addr_332_5, addr_positional[5319:5316], addr_1329_6);

wire[27:0] addr_1330_6;

Selector_2 s1330_6(wires_332_5[2], addr_332_5, addr_positional[5323:5320], addr_1330_6);

wire[27:0] addr_1331_6;

Selector_2 s1331_6(wires_332_5[3], addr_332_5, addr_positional[5327:5324], addr_1331_6);

wire[27:0] addr_1332_6;

Selector_2 s1332_6(wires_333_5[0], addr_333_5, addr_positional[5331:5328], addr_1332_6);

wire[27:0] addr_1333_6;

Selector_2 s1333_6(wires_333_5[1], addr_333_5, addr_positional[5335:5332], addr_1333_6);

wire[27:0] addr_1334_6;

Selector_2 s1334_6(wires_333_5[2], addr_333_5, addr_positional[5339:5336], addr_1334_6);

wire[27:0] addr_1335_6;

Selector_2 s1335_6(wires_333_5[3], addr_333_5, addr_positional[5343:5340], addr_1335_6);

wire[27:0] addr_1336_6;

Selector_2 s1336_6(wires_334_5[0], addr_334_5, addr_positional[5347:5344], addr_1336_6);

wire[27:0] addr_1337_6;

Selector_2 s1337_6(wires_334_5[1], addr_334_5, addr_positional[5351:5348], addr_1337_6);

wire[27:0] addr_1338_6;

Selector_2 s1338_6(wires_334_5[2], addr_334_5, addr_positional[5355:5352], addr_1338_6);

wire[27:0] addr_1339_6;

Selector_2 s1339_6(wires_334_5[3], addr_334_5, addr_positional[5359:5356], addr_1339_6);

wire[27:0] addr_1340_6;

Selector_2 s1340_6(wires_335_5[0], addr_335_5, addr_positional[5363:5360], addr_1340_6);

wire[27:0] addr_1341_6;

Selector_2 s1341_6(wires_335_5[1], addr_335_5, addr_positional[5367:5364], addr_1341_6);

wire[27:0] addr_1342_6;

Selector_2 s1342_6(wires_335_5[2], addr_335_5, addr_positional[5371:5368], addr_1342_6);

wire[27:0] addr_1343_6;

Selector_2 s1343_6(wires_335_5[3], addr_335_5, addr_positional[5375:5372], addr_1343_6);

wire[27:0] addr_1344_6;

Selector_2 s1344_6(wires_336_5[0], addr_336_5, addr_positional[5379:5376], addr_1344_6);

wire[27:0] addr_1345_6;

Selector_2 s1345_6(wires_336_5[1], addr_336_5, addr_positional[5383:5380], addr_1345_6);

wire[27:0] addr_1346_6;

Selector_2 s1346_6(wires_336_5[2], addr_336_5, addr_positional[5387:5384], addr_1346_6);

wire[27:0] addr_1347_6;

Selector_2 s1347_6(wires_336_5[3], addr_336_5, addr_positional[5391:5388], addr_1347_6);

wire[27:0] addr_1348_6;

Selector_2 s1348_6(wires_337_5[0], addr_337_5, addr_positional[5395:5392], addr_1348_6);

wire[27:0] addr_1349_6;

Selector_2 s1349_6(wires_337_5[1], addr_337_5, addr_positional[5399:5396], addr_1349_6);

wire[27:0] addr_1350_6;

Selector_2 s1350_6(wires_337_5[2], addr_337_5, addr_positional[5403:5400], addr_1350_6);

wire[27:0] addr_1351_6;

Selector_2 s1351_6(wires_337_5[3], addr_337_5, addr_positional[5407:5404], addr_1351_6);

wire[27:0] addr_1352_6;

Selector_2 s1352_6(wires_338_5[0], addr_338_5, addr_positional[5411:5408], addr_1352_6);

wire[27:0] addr_1353_6;

Selector_2 s1353_6(wires_338_5[1], addr_338_5, addr_positional[5415:5412], addr_1353_6);

wire[27:0] addr_1354_6;

Selector_2 s1354_6(wires_338_5[2], addr_338_5, addr_positional[5419:5416], addr_1354_6);

wire[27:0] addr_1355_6;

Selector_2 s1355_6(wires_338_5[3], addr_338_5, addr_positional[5423:5420], addr_1355_6);

wire[27:0] addr_1356_6;

Selector_2 s1356_6(wires_339_5[0], addr_339_5, addr_positional[5427:5424], addr_1356_6);

wire[27:0] addr_1357_6;

Selector_2 s1357_6(wires_339_5[1], addr_339_5, addr_positional[5431:5428], addr_1357_6);

wire[27:0] addr_1358_6;

Selector_2 s1358_6(wires_339_5[2], addr_339_5, addr_positional[5435:5432], addr_1358_6);

wire[27:0] addr_1359_6;

Selector_2 s1359_6(wires_339_5[3], addr_339_5, addr_positional[5439:5436], addr_1359_6);

wire[27:0] addr_1360_6;

Selector_2 s1360_6(wires_340_5[0], addr_340_5, addr_positional[5443:5440], addr_1360_6);

wire[27:0] addr_1361_6;

Selector_2 s1361_6(wires_340_5[1], addr_340_5, addr_positional[5447:5444], addr_1361_6);

wire[27:0] addr_1362_6;

Selector_2 s1362_6(wires_340_5[2], addr_340_5, addr_positional[5451:5448], addr_1362_6);

wire[27:0] addr_1363_6;

Selector_2 s1363_6(wires_340_5[3], addr_340_5, addr_positional[5455:5452], addr_1363_6);

wire[27:0] addr_1364_6;

Selector_2 s1364_6(wires_341_5[0], addr_341_5, addr_positional[5459:5456], addr_1364_6);

wire[27:0] addr_1365_6;

Selector_2 s1365_6(wires_341_5[1], addr_341_5, addr_positional[5463:5460], addr_1365_6);

wire[27:0] addr_1366_6;

Selector_2 s1366_6(wires_341_5[2], addr_341_5, addr_positional[5467:5464], addr_1366_6);

wire[27:0] addr_1367_6;

Selector_2 s1367_6(wires_341_5[3], addr_341_5, addr_positional[5471:5468], addr_1367_6);

wire[27:0] addr_1368_6;

Selector_2 s1368_6(wires_342_5[0], addr_342_5, addr_positional[5475:5472], addr_1368_6);

wire[27:0] addr_1369_6;

Selector_2 s1369_6(wires_342_5[1], addr_342_5, addr_positional[5479:5476], addr_1369_6);

wire[27:0] addr_1370_6;

Selector_2 s1370_6(wires_342_5[2], addr_342_5, addr_positional[5483:5480], addr_1370_6);

wire[27:0] addr_1371_6;

Selector_2 s1371_6(wires_342_5[3], addr_342_5, addr_positional[5487:5484], addr_1371_6);

wire[27:0] addr_1372_6;

Selector_2 s1372_6(wires_343_5[0], addr_343_5, addr_positional[5491:5488], addr_1372_6);

wire[27:0] addr_1373_6;

Selector_2 s1373_6(wires_343_5[1], addr_343_5, addr_positional[5495:5492], addr_1373_6);

wire[27:0] addr_1374_6;

Selector_2 s1374_6(wires_343_5[2], addr_343_5, addr_positional[5499:5496], addr_1374_6);

wire[27:0] addr_1375_6;

Selector_2 s1375_6(wires_343_5[3], addr_343_5, addr_positional[5503:5500], addr_1375_6);

wire[27:0] addr_1376_6;

Selector_2 s1376_6(wires_344_5[0], addr_344_5, addr_positional[5507:5504], addr_1376_6);

wire[27:0] addr_1377_6;

Selector_2 s1377_6(wires_344_5[1], addr_344_5, addr_positional[5511:5508], addr_1377_6);

wire[27:0] addr_1378_6;

Selector_2 s1378_6(wires_344_5[2], addr_344_5, addr_positional[5515:5512], addr_1378_6);

wire[27:0] addr_1379_6;

Selector_2 s1379_6(wires_344_5[3], addr_344_5, addr_positional[5519:5516], addr_1379_6);

wire[27:0] addr_1380_6;

Selector_2 s1380_6(wires_345_5[0], addr_345_5, addr_positional[5523:5520], addr_1380_6);

wire[27:0] addr_1381_6;

Selector_2 s1381_6(wires_345_5[1], addr_345_5, addr_positional[5527:5524], addr_1381_6);

wire[27:0] addr_1382_6;

Selector_2 s1382_6(wires_345_5[2], addr_345_5, addr_positional[5531:5528], addr_1382_6);

wire[27:0] addr_1383_6;

Selector_2 s1383_6(wires_345_5[3], addr_345_5, addr_positional[5535:5532], addr_1383_6);

wire[27:0] addr_1384_6;

Selector_2 s1384_6(wires_346_5[0], addr_346_5, addr_positional[5539:5536], addr_1384_6);

wire[27:0] addr_1385_6;

Selector_2 s1385_6(wires_346_5[1], addr_346_5, addr_positional[5543:5540], addr_1385_6);

wire[27:0] addr_1386_6;

Selector_2 s1386_6(wires_346_5[2], addr_346_5, addr_positional[5547:5544], addr_1386_6);

wire[27:0] addr_1387_6;

Selector_2 s1387_6(wires_346_5[3], addr_346_5, addr_positional[5551:5548], addr_1387_6);

wire[27:0] addr_1388_6;

Selector_2 s1388_6(wires_347_5[0], addr_347_5, addr_positional[5555:5552], addr_1388_6);

wire[27:0] addr_1389_6;

Selector_2 s1389_6(wires_347_5[1], addr_347_5, addr_positional[5559:5556], addr_1389_6);

wire[27:0] addr_1390_6;

Selector_2 s1390_6(wires_347_5[2], addr_347_5, addr_positional[5563:5560], addr_1390_6);

wire[27:0] addr_1391_6;

Selector_2 s1391_6(wires_347_5[3], addr_347_5, addr_positional[5567:5564], addr_1391_6);

wire[27:0] addr_1392_6;

Selector_2 s1392_6(wires_348_5[0], addr_348_5, addr_positional[5571:5568], addr_1392_6);

wire[27:0] addr_1393_6;

Selector_2 s1393_6(wires_348_5[1], addr_348_5, addr_positional[5575:5572], addr_1393_6);

wire[27:0] addr_1394_6;

Selector_2 s1394_6(wires_348_5[2], addr_348_5, addr_positional[5579:5576], addr_1394_6);

wire[27:0] addr_1395_6;

Selector_2 s1395_6(wires_348_5[3], addr_348_5, addr_positional[5583:5580], addr_1395_6);

wire[27:0] addr_1396_6;

Selector_2 s1396_6(wires_349_5[0], addr_349_5, addr_positional[5587:5584], addr_1396_6);

wire[27:0] addr_1397_6;

Selector_2 s1397_6(wires_349_5[1], addr_349_5, addr_positional[5591:5588], addr_1397_6);

wire[27:0] addr_1398_6;

Selector_2 s1398_6(wires_349_5[2], addr_349_5, addr_positional[5595:5592], addr_1398_6);

wire[27:0] addr_1399_6;

Selector_2 s1399_6(wires_349_5[3], addr_349_5, addr_positional[5599:5596], addr_1399_6);

wire[27:0] addr_1400_6;

Selector_2 s1400_6(wires_350_5[0], addr_350_5, addr_positional[5603:5600], addr_1400_6);

wire[27:0] addr_1401_6;

Selector_2 s1401_6(wires_350_5[1], addr_350_5, addr_positional[5607:5604], addr_1401_6);

wire[27:0] addr_1402_6;

Selector_2 s1402_6(wires_350_5[2], addr_350_5, addr_positional[5611:5608], addr_1402_6);

wire[27:0] addr_1403_6;

Selector_2 s1403_6(wires_350_5[3], addr_350_5, addr_positional[5615:5612], addr_1403_6);

wire[27:0] addr_1404_6;

Selector_2 s1404_6(wires_351_5[0], addr_351_5, addr_positional[5619:5616], addr_1404_6);

wire[27:0] addr_1405_6;

Selector_2 s1405_6(wires_351_5[1], addr_351_5, addr_positional[5623:5620], addr_1405_6);

wire[27:0] addr_1406_6;

Selector_2 s1406_6(wires_351_5[2], addr_351_5, addr_positional[5627:5624], addr_1406_6);

wire[27:0] addr_1407_6;

Selector_2 s1407_6(wires_351_5[3], addr_351_5, addr_positional[5631:5628], addr_1407_6);

wire[27:0] addr_1408_6;

Selector_2 s1408_6(wires_352_5[0], addr_352_5, addr_positional[5635:5632], addr_1408_6);

wire[27:0] addr_1409_6;

Selector_2 s1409_6(wires_352_5[1], addr_352_5, addr_positional[5639:5636], addr_1409_6);

wire[27:0] addr_1410_6;

Selector_2 s1410_6(wires_352_5[2], addr_352_5, addr_positional[5643:5640], addr_1410_6);

wire[27:0] addr_1411_6;

Selector_2 s1411_6(wires_352_5[3], addr_352_5, addr_positional[5647:5644], addr_1411_6);

wire[27:0] addr_1412_6;

Selector_2 s1412_6(wires_353_5[0], addr_353_5, addr_positional[5651:5648], addr_1412_6);

wire[27:0] addr_1413_6;

Selector_2 s1413_6(wires_353_5[1], addr_353_5, addr_positional[5655:5652], addr_1413_6);

wire[27:0] addr_1414_6;

Selector_2 s1414_6(wires_353_5[2], addr_353_5, addr_positional[5659:5656], addr_1414_6);

wire[27:0] addr_1415_6;

Selector_2 s1415_6(wires_353_5[3], addr_353_5, addr_positional[5663:5660], addr_1415_6);

wire[27:0] addr_1416_6;

Selector_2 s1416_6(wires_354_5[0], addr_354_5, addr_positional[5667:5664], addr_1416_6);

wire[27:0] addr_1417_6;

Selector_2 s1417_6(wires_354_5[1], addr_354_5, addr_positional[5671:5668], addr_1417_6);

wire[27:0] addr_1418_6;

Selector_2 s1418_6(wires_354_5[2], addr_354_5, addr_positional[5675:5672], addr_1418_6);

wire[27:0] addr_1419_6;

Selector_2 s1419_6(wires_354_5[3], addr_354_5, addr_positional[5679:5676], addr_1419_6);

wire[27:0] addr_1420_6;

Selector_2 s1420_6(wires_355_5[0], addr_355_5, addr_positional[5683:5680], addr_1420_6);

wire[27:0] addr_1421_6;

Selector_2 s1421_6(wires_355_5[1], addr_355_5, addr_positional[5687:5684], addr_1421_6);

wire[27:0] addr_1422_6;

Selector_2 s1422_6(wires_355_5[2], addr_355_5, addr_positional[5691:5688], addr_1422_6);

wire[27:0] addr_1423_6;

Selector_2 s1423_6(wires_355_5[3], addr_355_5, addr_positional[5695:5692], addr_1423_6);

wire[27:0] addr_1424_6;

Selector_2 s1424_6(wires_356_5[0], addr_356_5, addr_positional[5699:5696], addr_1424_6);

wire[27:0] addr_1425_6;

Selector_2 s1425_6(wires_356_5[1], addr_356_5, addr_positional[5703:5700], addr_1425_6);

wire[27:0] addr_1426_6;

Selector_2 s1426_6(wires_356_5[2], addr_356_5, addr_positional[5707:5704], addr_1426_6);

wire[27:0] addr_1427_6;

Selector_2 s1427_6(wires_356_5[3], addr_356_5, addr_positional[5711:5708], addr_1427_6);

wire[27:0] addr_1428_6;

Selector_2 s1428_6(wires_357_5[0], addr_357_5, addr_positional[5715:5712], addr_1428_6);

wire[27:0] addr_1429_6;

Selector_2 s1429_6(wires_357_5[1], addr_357_5, addr_positional[5719:5716], addr_1429_6);

wire[27:0] addr_1430_6;

Selector_2 s1430_6(wires_357_5[2], addr_357_5, addr_positional[5723:5720], addr_1430_6);

wire[27:0] addr_1431_6;

Selector_2 s1431_6(wires_357_5[3], addr_357_5, addr_positional[5727:5724], addr_1431_6);

wire[27:0] addr_1432_6;

Selector_2 s1432_6(wires_358_5[0], addr_358_5, addr_positional[5731:5728], addr_1432_6);

wire[27:0] addr_1433_6;

Selector_2 s1433_6(wires_358_5[1], addr_358_5, addr_positional[5735:5732], addr_1433_6);

wire[27:0] addr_1434_6;

Selector_2 s1434_6(wires_358_5[2], addr_358_5, addr_positional[5739:5736], addr_1434_6);

wire[27:0] addr_1435_6;

Selector_2 s1435_6(wires_358_5[3], addr_358_5, addr_positional[5743:5740], addr_1435_6);

wire[27:0] addr_1436_6;

Selector_2 s1436_6(wires_359_5[0], addr_359_5, addr_positional[5747:5744], addr_1436_6);

wire[27:0] addr_1437_6;

Selector_2 s1437_6(wires_359_5[1], addr_359_5, addr_positional[5751:5748], addr_1437_6);

wire[27:0] addr_1438_6;

Selector_2 s1438_6(wires_359_5[2], addr_359_5, addr_positional[5755:5752], addr_1438_6);

wire[27:0] addr_1439_6;

Selector_2 s1439_6(wires_359_5[3], addr_359_5, addr_positional[5759:5756], addr_1439_6);

wire[27:0] addr_1440_6;

Selector_2 s1440_6(wires_360_5[0], addr_360_5, addr_positional[5763:5760], addr_1440_6);

wire[27:0] addr_1441_6;

Selector_2 s1441_6(wires_360_5[1], addr_360_5, addr_positional[5767:5764], addr_1441_6);

wire[27:0] addr_1442_6;

Selector_2 s1442_6(wires_360_5[2], addr_360_5, addr_positional[5771:5768], addr_1442_6);

wire[27:0] addr_1443_6;

Selector_2 s1443_6(wires_360_5[3], addr_360_5, addr_positional[5775:5772], addr_1443_6);

wire[27:0] addr_1444_6;

Selector_2 s1444_6(wires_361_5[0], addr_361_5, addr_positional[5779:5776], addr_1444_6);

wire[27:0] addr_1445_6;

Selector_2 s1445_6(wires_361_5[1], addr_361_5, addr_positional[5783:5780], addr_1445_6);

wire[27:0] addr_1446_6;

Selector_2 s1446_6(wires_361_5[2], addr_361_5, addr_positional[5787:5784], addr_1446_6);

wire[27:0] addr_1447_6;

Selector_2 s1447_6(wires_361_5[3], addr_361_5, addr_positional[5791:5788], addr_1447_6);

wire[27:0] addr_1448_6;

Selector_2 s1448_6(wires_362_5[0], addr_362_5, addr_positional[5795:5792], addr_1448_6);

wire[27:0] addr_1449_6;

Selector_2 s1449_6(wires_362_5[1], addr_362_5, addr_positional[5799:5796], addr_1449_6);

wire[27:0] addr_1450_6;

Selector_2 s1450_6(wires_362_5[2], addr_362_5, addr_positional[5803:5800], addr_1450_6);

wire[27:0] addr_1451_6;

Selector_2 s1451_6(wires_362_5[3], addr_362_5, addr_positional[5807:5804], addr_1451_6);

wire[27:0] addr_1452_6;

Selector_2 s1452_6(wires_363_5[0], addr_363_5, addr_positional[5811:5808], addr_1452_6);

wire[27:0] addr_1453_6;

Selector_2 s1453_6(wires_363_5[1], addr_363_5, addr_positional[5815:5812], addr_1453_6);

wire[27:0] addr_1454_6;

Selector_2 s1454_6(wires_363_5[2], addr_363_5, addr_positional[5819:5816], addr_1454_6);

wire[27:0] addr_1455_6;

Selector_2 s1455_6(wires_363_5[3], addr_363_5, addr_positional[5823:5820], addr_1455_6);

wire[27:0] addr_1456_6;

Selector_2 s1456_6(wires_364_5[0], addr_364_5, addr_positional[5827:5824], addr_1456_6);

wire[27:0] addr_1457_6;

Selector_2 s1457_6(wires_364_5[1], addr_364_5, addr_positional[5831:5828], addr_1457_6);

wire[27:0] addr_1458_6;

Selector_2 s1458_6(wires_364_5[2], addr_364_5, addr_positional[5835:5832], addr_1458_6);

wire[27:0] addr_1459_6;

Selector_2 s1459_6(wires_364_5[3], addr_364_5, addr_positional[5839:5836], addr_1459_6);

wire[27:0] addr_1460_6;

Selector_2 s1460_6(wires_365_5[0], addr_365_5, addr_positional[5843:5840], addr_1460_6);

wire[27:0] addr_1461_6;

Selector_2 s1461_6(wires_365_5[1], addr_365_5, addr_positional[5847:5844], addr_1461_6);

wire[27:0] addr_1462_6;

Selector_2 s1462_6(wires_365_5[2], addr_365_5, addr_positional[5851:5848], addr_1462_6);

wire[27:0] addr_1463_6;

Selector_2 s1463_6(wires_365_5[3], addr_365_5, addr_positional[5855:5852], addr_1463_6);

wire[27:0] addr_1464_6;

Selector_2 s1464_6(wires_366_5[0], addr_366_5, addr_positional[5859:5856], addr_1464_6);

wire[27:0] addr_1465_6;

Selector_2 s1465_6(wires_366_5[1], addr_366_5, addr_positional[5863:5860], addr_1465_6);

wire[27:0] addr_1466_6;

Selector_2 s1466_6(wires_366_5[2], addr_366_5, addr_positional[5867:5864], addr_1466_6);

wire[27:0] addr_1467_6;

Selector_2 s1467_6(wires_366_5[3], addr_366_5, addr_positional[5871:5868], addr_1467_6);

wire[27:0] addr_1468_6;

Selector_2 s1468_6(wires_367_5[0], addr_367_5, addr_positional[5875:5872], addr_1468_6);

wire[27:0] addr_1469_6;

Selector_2 s1469_6(wires_367_5[1], addr_367_5, addr_positional[5879:5876], addr_1469_6);

wire[27:0] addr_1470_6;

Selector_2 s1470_6(wires_367_5[2], addr_367_5, addr_positional[5883:5880], addr_1470_6);

wire[27:0] addr_1471_6;

Selector_2 s1471_6(wires_367_5[3], addr_367_5, addr_positional[5887:5884], addr_1471_6);

wire[27:0] addr_1472_6;

Selector_2 s1472_6(wires_368_5[0], addr_368_5, addr_positional[5891:5888], addr_1472_6);

wire[27:0] addr_1473_6;

Selector_2 s1473_6(wires_368_5[1], addr_368_5, addr_positional[5895:5892], addr_1473_6);

wire[27:0] addr_1474_6;

Selector_2 s1474_6(wires_368_5[2], addr_368_5, addr_positional[5899:5896], addr_1474_6);

wire[27:0] addr_1475_6;

Selector_2 s1475_6(wires_368_5[3], addr_368_5, addr_positional[5903:5900], addr_1475_6);

wire[27:0] addr_1476_6;

Selector_2 s1476_6(wires_369_5[0], addr_369_5, addr_positional[5907:5904], addr_1476_6);

wire[27:0] addr_1477_6;

Selector_2 s1477_6(wires_369_5[1], addr_369_5, addr_positional[5911:5908], addr_1477_6);

wire[27:0] addr_1478_6;

Selector_2 s1478_6(wires_369_5[2], addr_369_5, addr_positional[5915:5912], addr_1478_6);

wire[27:0] addr_1479_6;

Selector_2 s1479_6(wires_369_5[3], addr_369_5, addr_positional[5919:5916], addr_1479_6);

wire[27:0] addr_1480_6;

Selector_2 s1480_6(wires_370_5[0], addr_370_5, addr_positional[5923:5920], addr_1480_6);

wire[27:0] addr_1481_6;

Selector_2 s1481_6(wires_370_5[1], addr_370_5, addr_positional[5927:5924], addr_1481_6);

wire[27:0] addr_1482_6;

Selector_2 s1482_6(wires_370_5[2], addr_370_5, addr_positional[5931:5928], addr_1482_6);

wire[27:0] addr_1483_6;

Selector_2 s1483_6(wires_370_5[3], addr_370_5, addr_positional[5935:5932], addr_1483_6);

wire[27:0] addr_1484_6;

Selector_2 s1484_6(wires_371_5[0], addr_371_5, addr_positional[5939:5936], addr_1484_6);

wire[27:0] addr_1485_6;

Selector_2 s1485_6(wires_371_5[1], addr_371_5, addr_positional[5943:5940], addr_1485_6);

wire[27:0] addr_1486_6;

Selector_2 s1486_6(wires_371_5[2], addr_371_5, addr_positional[5947:5944], addr_1486_6);

wire[27:0] addr_1487_6;

Selector_2 s1487_6(wires_371_5[3], addr_371_5, addr_positional[5951:5948], addr_1487_6);

wire[27:0] addr_1488_6;

Selector_2 s1488_6(wires_372_5[0], addr_372_5, addr_positional[5955:5952], addr_1488_6);

wire[27:0] addr_1489_6;

Selector_2 s1489_6(wires_372_5[1], addr_372_5, addr_positional[5959:5956], addr_1489_6);

wire[27:0] addr_1490_6;

Selector_2 s1490_6(wires_372_5[2], addr_372_5, addr_positional[5963:5960], addr_1490_6);

wire[27:0] addr_1491_6;

Selector_2 s1491_6(wires_372_5[3], addr_372_5, addr_positional[5967:5964], addr_1491_6);

wire[27:0] addr_1492_6;

Selector_2 s1492_6(wires_373_5[0], addr_373_5, addr_positional[5971:5968], addr_1492_6);

wire[27:0] addr_1493_6;

Selector_2 s1493_6(wires_373_5[1], addr_373_5, addr_positional[5975:5972], addr_1493_6);

wire[27:0] addr_1494_6;

Selector_2 s1494_6(wires_373_5[2], addr_373_5, addr_positional[5979:5976], addr_1494_6);

wire[27:0] addr_1495_6;

Selector_2 s1495_6(wires_373_5[3], addr_373_5, addr_positional[5983:5980], addr_1495_6);

wire[27:0] addr_1496_6;

Selector_2 s1496_6(wires_374_5[0], addr_374_5, addr_positional[5987:5984], addr_1496_6);

wire[27:0] addr_1497_6;

Selector_2 s1497_6(wires_374_5[1], addr_374_5, addr_positional[5991:5988], addr_1497_6);

wire[27:0] addr_1498_6;

Selector_2 s1498_6(wires_374_5[2], addr_374_5, addr_positional[5995:5992], addr_1498_6);

wire[27:0] addr_1499_6;

Selector_2 s1499_6(wires_374_5[3], addr_374_5, addr_positional[5999:5996], addr_1499_6);

wire[27:0] addr_1500_6;

Selector_2 s1500_6(wires_375_5[0], addr_375_5, addr_positional[6003:6000], addr_1500_6);

wire[27:0] addr_1501_6;

Selector_2 s1501_6(wires_375_5[1], addr_375_5, addr_positional[6007:6004], addr_1501_6);

wire[27:0] addr_1502_6;

Selector_2 s1502_6(wires_375_5[2], addr_375_5, addr_positional[6011:6008], addr_1502_6);

wire[27:0] addr_1503_6;

Selector_2 s1503_6(wires_375_5[3], addr_375_5, addr_positional[6015:6012], addr_1503_6);

wire[27:0] addr_1504_6;

Selector_2 s1504_6(wires_376_5[0], addr_376_5, addr_positional[6019:6016], addr_1504_6);

wire[27:0] addr_1505_6;

Selector_2 s1505_6(wires_376_5[1], addr_376_5, addr_positional[6023:6020], addr_1505_6);

wire[27:0] addr_1506_6;

Selector_2 s1506_6(wires_376_5[2], addr_376_5, addr_positional[6027:6024], addr_1506_6);

wire[27:0] addr_1507_6;

Selector_2 s1507_6(wires_376_5[3], addr_376_5, addr_positional[6031:6028], addr_1507_6);

wire[27:0] addr_1508_6;

Selector_2 s1508_6(wires_377_5[0], addr_377_5, addr_positional[6035:6032], addr_1508_6);

wire[27:0] addr_1509_6;

Selector_2 s1509_6(wires_377_5[1], addr_377_5, addr_positional[6039:6036], addr_1509_6);

wire[27:0] addr_1510_6;

Selector_2 s1510_6(wires_377_5[2], addr_377_5, addr_positional[6043:6040], addr_1510_6);

wire[27:0] addr_1511_6;

Selector_2 s1511_6(wires_377_5[3], addr_377_5, addr_positional[6047:6044], addr_1511_6);

wire[27:0] addr_1512_6;

Selector_2 s1512_6(wires_378_5[0], addr_378_5, addr_positional[6051:6048], addr_1512_6);

wire[27:0] addr_1513_6;

Selector_2 s1513_6(wires_378_5[1], addr_378_5, addr_positional[6055:6052], addr_1513_6);

wire[27:0] addr_1514_6;

Selector_2 s1514_6(wires_378_5[2], addr_378_5, addr_positional[6059:6056], addr_1514_6);

wire[27:0] addr_1515_6;

Selector_2 s1515_6(wires_378_5[3], addr_378_5, addr_positional[6063:6060], addr_1515_6);

wire[27:0] addr_1516_6;

Selector_2 s1516_6(wires_379_5[0], addr_379_5, addr_positional[6067:6064], addr_1516_6);

wire[27:0] addr_1517_6;

Selector_2 s1517_6(wires_379_5[1], addr_379_5, addr_positional[6071:6068], addr_1517_6);

wire[27:0] addr_1518_6;

Selector_2 s1518_6(wires_379_5[2], addr_379_5, addr_positional[6075:6072], addr_1518_6);

wire[27:0] addr_1519_6;

Selector_2 s1519_6(wires_379_5[3], addr_379_5, addr_positional[6079:6076], addr_1519_6);

wire[27:0] addr_1520_6;

Selector_2 s1520_6(wires_380_5[0], addr_380_5, addr_positional[6083:6080], addr_1520_6);

wire[27:0] addr_1521_6;

Selector_2 s1521_6(wires_380_5[1], addr_380_5, addr_positional[6087:6084], addr_1521_6);

wire[27:0] addr_1522_6;

Selector_2 s1522_6(wires_380_5[2], addr_380_5, addr_positional[6091:6088], addr_1522_6);

wire[27:0] addr_1523_6;

Selector_2 s1523_6(wires_380_5[3], addr_380_5, addr_positional[6095:6092], addr_1523_6);

wire[27:0] addr_1524_6;

Selector_2 s1524_6(wires_381_5[0], addr_381_5, addr_positional[6099:6096], addr_1524_6);

wire[27:0] addr_1525_6;

Selector_2 s1525_6(wires_381_5[1], addr_381_5, addr_positional[6103:6100], addr_1525_6);

wire[27:0] addr_1526_6;

Selector_2 s1526_6(wires_381_5[2], addr_381_5, addr_positional[6107:6104], addr_1526_6);

wire[27:0] addr_1527_6;

Selector_2 s1527_6(wires_381_5[3], addr_381_5, addr_positional[6111:6108], addr_1527_6);

wire[27:0] addr_1528_6;

Selector_2 s1528_6(wires_382_5[0], addr_382_5, addr_positional[6115:6112], addr_1528_6);

wire[27:0] addr_1529_6;

Selector_2 s1529_6(wires_382_5[1], addr_382_5, addr_positional[6119:6116], addr_1529_6);

wire[27:0] addr_1530_6;

Selector_2 s1530_6(wires_382_5[2], addr_382_5, addr_positional[6123:6120], addr_1530_6);

wire[27:0] addr_1531_6;

Selector_2 s1531_6(wires_382_5[3], addr_382_5, addr_positional[6127:6124], addr_1531_6);

wire[27:0] addr_1532_6;

Selector_2 s1532_6(wires_383_5[0], addr_383_5, addr_positional[6131:6128], addr_1532_6);

wire[27:0] addr_1533_6;

Selector_2 s1533_6(wires_383_5[1], addr_383_5, addr_positional[6135:6132], addr_1533_6);

wire[27:0] addr_1534_6;

Selector_2 s1534_6(wires_383_5[2], addr_383_5, addr_positional[6139:6136], addr_1534_6);

wire[27:0] addr_1535_6;

Selector_2 s1535_6(wires_383_5[3], addr_383_5, addr_positional[6143:6140], addr_1535_6);

wire[27:0] addr_1536_6;

Selector_2 s1536_6(wires_384_5[0], addr_384_5, addr_positional[6147:6144], addr_1536_6);

wire[27:0] addr_1537_6;

Selector_2 s1537_6(wires_384_5[1], addr_384_5, addr_positional[6151:6148], addr_1537_6);

wire[27:0] addr_1538_6;

Selector_2 s1538_6(wires_384_5[2], addr_384_5, addr_positional[6155:6152], addr_1538_6);

wire[27:0] addr_1539_6;

Selector_2 s1539_6(wires_384_5[3], addr_384_5, addr_positional[6159:6156], addr_1539_6);

wire[27:0] addr_1540_6;

Selector_2 s1540_6(wires_385_5[0], addr_385_5, addr_positional[6163:6160], addr_1540_6);

wire[27:0] addr_1541_6;

Selector_2 s1541_6(wires_385_5[1], addr_385_5, addr_positional[6167:6164], addr_1541_6);

wire[27:0] addr_1542_6;

Selector_2 s1542_6(wires_385_5[2], addr_385_5, addr_positional[6171:6168], addr_1542_6);

wire[27:0] addr_1543_6;

Selector_2 s1543_6(wires_385_5[3], addr_385_5, addr_positional[6175:6172], addr_1543_6);

wire[27:0] addr_1544_6;

Selector_2 s1544_6(wires_386_5[0], addr_386_5, addr_positional[6179:6176], addr_1544_6);

wire[27:0] addr_1545_6;

Selector_2 s1545_6(wires_386_5[1], addr_386_5, addr_positional[6183:6180], addr_1545_6);

wire[27:0] addr_1546_6;

Selector_2 s1546_6(wires_386_5[2], addr_386_5, addr_positional[6187:6184], addr_1546_6);

wire[27:0] addr_1547_6;

Selector_2 s1547_6(wires_386_5[3], addr_386_5, addr_positional[6191:6188], addr_1547_6);

wire[27:0] addr_1548_6;

Selector_2 s1548_6(wires_387_5[0], addr_387_5, addr_positional[6195:6192], addr_1548_6);

wire[27:0] addr_1549_6;

Selector_2 s1549_6(wires_387_5[1], addr_387_5, addr_positional[6199:6196], addr_1549_6);

wire[27:0] addr_1550_6;

Selector_2 s1550_6(wires_387_5[2], addr_387_5, addr_positional[6203:6200], addr_1550_6);

wire[27:0] addr_1551_6;

Selector_2 s1551_6(wires_387_5[3], addr_387_5, addr_positional[6207:6204], addr_1551_6);

wire[27:0] addr_1552_6;

Selector_2 s1552_6(wires_388_5[0], addr_388_5, addr_positional[6211:6208], addr_1552_6);

wire[27:0] addr_1553_6;

Selector_2 s1553_6(wires_388_5[1], addr_388_5, addr_positional[6215:6212], addr_1553_6);

wire[27:0] addr_1554_6;

Selector_2 s1554_6(wires_388_5[2], addr_388_5, addr_positional[6219:6216], addr_1554_6);

wire[27:0] addr_1555_6;

Selector_2 s1555_6(wires_388_5[3], addr_388_5, addr_positional[6223:6220], addr_1555_6);

wire[27:0] addr_1556_6;

Selector_2 s1556_6(wires_389_5[0], addr_389_5, addr_positional[6227:6224], addr_1556_6);

wire[27:0] addr_1557_6;

Selector_2 s1557_6(wires_389_5[1], addr_389_5, addr_positional[6231:6228], addr_1557_6);

wire[27:0] addr_1558_6;

Selector_2 s1558_6(wires_389_5[2], addr_389_5, addr_positional[6235:6232], addr_1558_6);

wire[27:0] addr_1559_6;

Selector_2 s1559_6(wires_389_5[3], addr_389_5, addr_positional[6239:6236], addr_1559_6);

wire[27:0] addr_1560_6;

Selector_2 s1560_6(wires_390_5[0], addr_390_5, addr_positional[6243:6240], addr_1560_6);

wire[27:0] addr_1561_6;

Selector_2 s1561_6(wires_390_5[1], addr_390_5, addr_positional[6247:6244], addr_1561_6);

wire[27:0] addr_1562_6;

Selector_2 s1562_6(wires_390_5[2], addr_390_5, addr_positional[6251:6248], addr_1562_6);

wire[27:0] addr_1563_6;

Selector_2 s1563_6(wires_390_5[3], addr_390_5, addr_positional[6255:6252], addr_1563_6);

wire[27:0] addr_1564_6;

Selector_2 s1564_6(wires_391_5[0], addr_391_5, addr_positional[6259:6256], addr_1564_6);

wire[27:0] addr_1565_6;

Selector_2 s1565_6(wires_391_5[1], addr_391_5, addr_positional[6263:6260], addr_1565_6);

wire[27:0] addr_1566_6;

Selector_2 s1566_6(wires_391_5[2], addr_391_5, addr_positional[6267:6264], addr_1566_6);

wire[27:0] addr_1567_6;

Selector_2 s1567_6(wires_391_5[3], addr_391_5, addr_positional[6271:6268], addr_1567_6);

wire[27:0] addr_1568_6;

Selector_2 s1568_6(wires_392_5[0], addr_392_5, addr_positional[6275:6272], addr_1568_6);

wire[27:0] addr_1569_6;

Selector_2 s1569_6(wires_392_5[1], addr_392_5, addr_positional[6279:6276], addr_1569_6);

wire[27:0] addr_1570_6;

Selector_2 s1570_6(wires_392_5[2], addr_392_5, addr_positional[6283:6280], addr_1570_6);

wire[27:0] addr_1571_6;

Selector_2 s1571_6(wires_392_5[3], addr_392_5, addr_positional[6287:6284], addr_1571_6);

wire[27:0] addr_1572_6;

Selector_2 s1572_6(wires_393_5[0], addr_393_5, addr_positional[6291:6288], addr_1572_6);

wire[27:0] addr_1573_6;

Selector_2 s1573_6(wires_393_5[1], addr_393_5, addr_positional[6295:6292], addr_1573_6);

wire[27:0] addr_1574_6;

Selector_2 s1574_6(wires_393_5[2], addr_393_5, addr_positional[6299:6296], addr_1574_6);

wire[27:0] addr_1575_6;

Selector_2 s1575_6(wires_393_5[3], addr_393_5, addr_positional[6303:6300], addr_1575_6);

wire[27:0] addr_1576_6;

Selector_2 s1576_6(wires_394_5[0], addr_394_5, addr_positional[6307:6304], addr_1576_6);

wire[27:0] addr_1577_6;

Selector_2 s1577_6(wires_394_5[1], addr_394_5, addr_positional[6311:6308], addr_1577_6);

wire[27:0] addr_1578_6;

Selector_2 s1578_6(wires_394_5[2], addr_394_5, addr_positional[6315:6312], addr_1578_6);

wire[27:0] addr_1579_6;

Selector_2 s1579_6(wires_394_5[3], addr_394_5, addr_positional[6319:6316], addr_1579_6);

wire[27:0] addr_1580_6;

Selector_2 s1580_6(wires_395_5[0], addr_395_5, addr_positional[6323:6320], addr_1580_6);

wire[27:0] addr_1581_6;

Selector_2 s1581_6(wires_395_5[1], addr_395_5, addr_positional[6327:6324], addr_1581_6);

wire[27:0] addr_1582_6;

Selector_2 s1582_6(wires_395_5[2], addr_395_5, addr_positional[6331:6328], addr_1582_6);

wire[27:0] addr_1583_6;

Selector_2 s1583_6(wires_395_5[3], addr_395_5, addr_positional[6335:6332], addr_1583_6);

wire[27:0] addr_1584_6;

Selector_2 s1584_6(wires_396_5[0], addr_396_5, addr_positional[6339:6336], addr_1584_6);

wire[27:0] addr_1585_6;

Selector_2 s1585_6(wires_396_5[1], addr_396_5, addr_positional[6343:6340], addr_1585_6);

wire[27:0] addr_1586_6;

Selector_2 s1586_6(wires_396_5[2], addr_396_5, addr_positional[6347:6344], addr_1586_6);

wire[27:0] addr_1587_6;

Selector_2 s1587_6(wires_396_5[3], addr_396_5, addr_positional[6351:6348], addr_1587_6);

wire[27:0] addr_1588_6;

Selector_2 s1588_6(wires_397_5[0], addr_397_5, addr_positional[6355:6352], addr_1588_6);

wire[27:0] addr_1589_6;

Selector_2 s1589_6(wires_397_5[1], addr_397_5, addr_positional[6359:6356], addr_1589_6);

wire[27:0] addr_1590_6;

Selector_2 s1590_6(wires_397_5[2], addr_397_5, addr_positional[6363:6360], addr_1590_6);

wire[27:0] addr_1591_6;

Selector_2 s1591_6(wires_397_5[3], addr_397_5, addr_positional[6367:6364], addr_1591_6);

wire[27:0] addr_1592_6;

Selector_2 s1592_6(wires_398_5[0], addr_398_5, addr_positional[6371:6368], addr_1592_6);

wire[27:0] addr_1593_6;

Selector_2 s1593_6(wires_398_5[1], addr_398_5, addr_positional[6375:6372], addr_1593_6);

wire[27:0] addr_1594_6;

Selector_2 s1594_6(wires_398_5[2], addr_398_5, addr_positional[6379:6376], addr_1594_6);

wire[27:0] addr_1595_6;

Selector_2 s1595_6(wires_398_5[3], addr_398_5, addr_positional[6383:6380], addr_1595_6);

wire[27:0] addr_1596_6;

Selector_2 s1596_6(wires_399_5[0], addr_399_5, addr_positional[6387:6384], addr_1596_6);

wire[27:0] addr_1597_6;

Selector_2 s1597_6(wires_399_5[1], addr_399_5, addr_positional[6391:6388], addr_1597_6);

wire[27:0] addr_1598_6;

Selector_2 s1598_6(wires_399_5[2], addr_399_5, addr_positional[6395:6392], addr_1598_6);

wire[27:0] addr_1599_6;

Selector_2 s1599_6(wires_399_5[3], addr_399_5, addr_positional[6399:6396], addr_1599_6);

wire[27:0] addr_1600_6;

Selector_2 s1600_6(wires_400_5[0], addr_400_5, addr_positional[6403:6400], addr_1600_6);

wire[27:0] addr_1601_6;

Selector_2 s1601_6(wires_400_5[1], addr_400_5, addr_positional[6407:6404], addr_1601_6);

wire[27:0] addr_1602_6;

Selector_2 s1602_6(wires_400_5[2], addr_400_5, addr_positional[6411:6408], addr_1602_6);

wire[27:0] addr_1603_6;

Selector_2 s1603_6(wires_400_5[3], addr_400_5, addr_positional[6415:6412], addr_1603_6);

wire[27:0] addr_1604_6;

Selector_2 s1604_6(wires_401_5[0], addr_401_5, addr_positional[6419:6416], addr_1604_6);

wire[27:0] addr_1605_6;

Selector_2 s1605_6(wires_401_5[1], addr_401_5, addr_positional[6423:6420], addr_1605_6);

wire[27:0] addr_1606_6;

Selector_2 s1606_6(wires_401_5[2], addr_401_5, addr_positional[6427:6424], addr_1606_6);

wire[27:0] addr_1607_6;

Selector_2 s1607_6(wires_401_5[3], addr_401_5, addr_positional[6431:6428], addr_1607_6);

wire[27:0] addr_1608_6;

Selector_2 s1608_6(wires_402_5[0], addr_402_5, addr_positional[6435:6432], addr_1608_6);

wire[27:0] addr_1609_6;

Selector_2 s1609_6(wires_402_5[1], addr_402_5, addr_positional[6439:6436], addr_1609_6);

wire[27:0] addr_1610_6;

Selector_2 s1610_6(wires_402_5[2], addr_402_5, addr_positional[6443:6440], addr_1610_6);

wire[27:0] addr_1611_6;

Selector_2 s1611_6(wires_402_5[3], addr_402_5, addr_positional[6447:6444], addr_1611_6);

wire[27:0] addr_1612_6;

Selector_2 s1612_6(wires_403_5[0], addr_403_5, addr_positional[6451:6448], addr_1612_6);

wire[27:0] addr_1613_6;

Selector_2 s1613_6(wires_403_5[1], addr_403_5, addr_positional[6455:6452], addr_1613_6);

wire[27:0] addr_1614_6;

Selector_2 s1614_6(wires_403_5[2], addr_403_5, addr_positional[6459:6456], addr_1614_6);

wire[27:0] addr_1615_6;

Selector_2 s1615_6(wires_403_5[3], addr_403_5, addr_positional[6463:6460], addr_1615_6);

wire[27:0] addr_1616_6;

Selector_2 s1616_6(wires_404_5[0], addr_404_5, addr_positional[6467:6464], addr_1616_6);

wire[27:0] addr_1617_6;

Selector_2 s1617_6(wires_404_5[1], addr_404_5, addr_positional[6471:6468], addr_1617_6);

wire[27:0] addr_1618_6;

Selector_2 s1618_6(wires_404_5[2], addr_404_5, addr_positional[6475:6472], addr_1618_6);

wire[27:0] addr_1619_6;

Selector_2 s1619_6(wires_404_5[3], addr_404_5, addr_positional[6479:6476], addr_1619_6);

wire[27:0] addr_1620_6;

Selector_2 s1620_6(wires_405_5[0], addr_405_5, addr_positional[6483:6480], addr_1620_6);

wire[27:0] addr_1621_6;

Selector_2 s1621_6(wires_405_5[1], addr_405_5, addr_positional[6487:6484], addr_1621_6);

wire[27:0] addr_1622_6;

Selector_2 s1622_6(wires_405_5[2], addr_405_5, addr_positional[6491:6488], addr_1622_6);

wire[27:0] addr_1623_6;

Selector_2 s1623_6(wires_405_5[3], addr_405_5, addr_positional[6495:6492], addr_1623_6);

wire[27:0] addr_1624_6;

Selector_2 s1624_6(wires_406_5[0], addr_406_5, addr_positional[6499:6496], addr_1624_6);

wire[27:0] addr_1625_6;

Selector_2 s1625_6(wires_406_5[1], addr_406_5, addr_positional[6503:6500], addr_1625_6);

wire[27:0] addr_1626_6;

Selector_2 s1626_6(wires_406_5[2], addr_406_5, addr_positional[6507:6504], addr_1626_6);

wire[27:0] addr_1627_6;

Selector_2 s1627_6(wires_406_5[3], addr_406_5, addr_positional[6511:6508], addr_1627_6);

wire[27:0] addr_1628_6;

Selector_2 s1628_6(wires_407_5[0], addr_407_5, addr_positional[6515:6512], addr_1628_6);

wire[27:0] addr_1629_6;

Selector_2 s1629_6(wires_407_5[1], addr_407_5, addr_positional[6519:6516], addr_1629_6);

wire[27:0] addr_1630_6;

Selector_2 s1630_6(wires_407_5[2], addr_407_5, addr_positional[6523:6520], addr_1630_6);

wire[27:0] addr_1631_6;

Selector_2 s1631_6(wires_407_5[3], addr_407_5, addr_positional[6527:6524], addr_1631_6);

wire[27:0] addr_1632_6;

Selector_2 s1632_6(wires_408_5[0], addr_408_5, addr_positional[6531:6528], addr_1632_6);

wire[27:0] addr_1633_6;

Selector_2 s1633_6(wires_408_5[1], addr_408_5, addr_positional[6535:6532], addr_1633_6);

wire[27:0] addr_1634_6;

Selector_2 s1634_6(wires_408_5[2], addr_408_5, addr_positional[6539:6536], addr_1634_6);

wire[27:0] addr_1635_6;

Selector_2 s1635_6(wires_408_5[3], addr_408_5, addr_positional[6543:6540], addr_1635_6);

wire[27:0] addr_1636_6;

Selector_2 s1636_6(wires_409_5[0], addr_409_5, addr_positional[6547:6544], addr_1636_6);

wire[27:0] addr_1637_6;

Selector_2 s1637_6(wires_409_5[1], addr_409_5, addr_positional[6551:6548], addr_1637_6);

wire[27:0] addr_1638_6;

Selector_2 s1638_6(wires_409_5[2], addr_409_5, addr_positional[6555:6552], addr_1638_6);

wire[27:0] addr_1639_6;

Selector_2 s1639_6(wires_409_5[3], addr_409_5, addr_positional[6559:6556], addr_1639_6);

wire[27:0] addr_1640_6;

Selector_2 s1640_6(wires_410_5[0], addr_410_5, addr_positional[6563:6560], addr_1640_6);

wire[27:0] addr_1641_6;

Selector_2 s1641_6(wires_410_5[1], addr_410_5, addr_positional[6567:6564], addr_1641_6);

wire[27:0] addr_1642_6;

Selector_2 s1642_6(wires_410_5[2], addr_410_5, addr_positional[6571:6568], addr_1642_6);

wire[27:0] addr_1643_6;

Selector_2 s1643_6(wires_410_5[3], addr_410_5, addr_positional[6575:6572], addr_1643_6);

wire[27:0] addr_1644_6;

Selector_2 s1644_6(wires_411_5[0], addr_411_5, addr_positional[6579:6576], addr_1644_6);

wire[27:0] addr_1645_6;

Selector_2 s1645_6(wires_411_5[1], addr_411_5, addr_positional[6583:6580], addr_1645_6);

wire[27:0] addr_1646_6;

Selector_2 s1646_6(wires_411_5[2], addr_411_5, addr_positional[6587:6584], addr_1646_6);

wire[27:0] addr_1647_6;

Selector_2 s1647_6(wires_411_5[3], addr_411_5, addr_positional[6591:6588], addr_1647_6);

wire[27:0] addr_1648_6;

Selector_2 s1648_6(wires_412_5[0], addr_412_5, addr_positional[6595:6592], addr_1648_6);

wire[27:0] addr_1649_6;

Selector_2 s1649_6(wires_412_5[1], addr_412_5, addr_positional[6599:6596], addr_1649_6);

wire[27:0] addr_1650_6;

Selector_2 s1650_6(wires_412_5[2], addr_412_5, addr_positional[6603:6600], addr_1650_6);

wire[27:0] addr_1651_6;

Selector_2 s1651_6(wires_412_5[3], addr_412_5, addr_positional[6607:6604], addr_1651_6);

wire[27:0] addr_1652_6;

Selector_2 s1652_6(wires_413_5[0], addr_413_5, addr_positional[6611:6608], addr_1652_6);

wire[27:0] addr_1653_6;

Selector_2 s1653_6(wires_413_5[1], addr_413_5, addr_positional[6615:6612], addr_1653_6);

wire[27:0] addr_1654_6;

Selector_2 s1654_6(wires_413_5[2], addr_413_5, addr_positional[6619:6616], addr_1654_6);

wire[27:0] addr_1655_6;

Selector_2 s1655_6(wires_413_5[3], addr_413_5, addr_positional[6623:6620], addr_1655_6);

wire[27:0] addr_1656_6;

Selector_2 s1656_6(wires_414_5[0], addr_414_5, addr_positional[6627:6624], addr_1656_6);

wire[27:0] addr_1657_6;

Selector_2 s1657_6(wires_414_5[1], addr_414_5, addr_positional[6631:6628], addr_1657_6);

wire[27:0] addr_1658_6;

Selector_2 s1658_6(wires_414_5[2], addr_414_5, addr_positional[6635:6632], addr_1658_6);

wire[27:0] addr_1659_6;

Selector_2 s1659_6(wires_414_5[3], addr_414_5, addr_positional[6639:6636], addr_1659_6);

wire[27:0] addr_1660_6;

Selector_2 s1660_6(wires_415_5[0], addr_415_5, addr_positional[6643:6640], addr_1660_6);

wire[27:0] addr_1661_6;

Selector_2 s1661_6(wires_415_5[1], addr_415_5, addr_positional[6647:6644], addr_1661_6);

wire[27:0] addr_1662_6;

Selector_2 s1662_6(wires_415_5[2], addr_415_5, addr_positional[6651:6648], addr_1662_6);

wire[27:0] addr_1663_6;

Selector_2 s1663_6(wires_415_5[3], addr_415_5, addr_positional[6655:6652], addr_1663_6);

wire[27:0] addr_1664_6;

Selector_2 s1664_6(wires_416_5[0], addr_416_5, addr_positional[6659:6656], addr_1664_6);

wire[27:0] addr_1665_6;

Selector_2 s1665_6(wires_416_5[1], addr_416_5, addr_positional[6663:6660], addr_1665_6);

wire[27:0] addr_1666_6;

Selector_2 s1666_6(wires_416_5[2], addr_416_5, addr_positional[6667:6664], addr_1666_6);

wire[27:0] addr_1667_6;

Selector_2 s1667_6(wires_416_5[3], addr_416_5, addr_positional[6671:6668], addr_1667_6);

wire[27:0] addr_1668_6;

Selector_2 s1668_6(wires_417_5[0], addr_417_5, addr_positional[6675:6672], addr_1668_6);

wire[27:0] addr_1669_6;

Selector_2 s1669_6(wires_417_5[1], addr_417_5, addr_positional[6679:6676], addr_1669_6);

wire[27:0] addr_1670_6;

Selector_2 s1670_6(wires_417_5[2], addr_417_5, addr_positional[6683:6680], addr_1670_6);

wire[27:0] addr_1671_6;

Selector_2 s1671_6(wires_417_5[3], addr_417_5, addr_positional[6687:6684], addr_1671_6);

wire[27:0] addr_1672_6;

Selector_2 s1672_6(wires_418_5[0], addr_418_5, addr_positional[6691:6688], addr_1672_6);

wire[27:0] addr_1673_6;

Selector_2 s1673_6(wires_418_5[1], addr_418_5, addr_positional[6695:6692], addr_1673_6);

wire[27:0] addr_1674_6;

Selector_2 s1674_6(wires_418_5[2], addr_418_5, addr_positional[6699:6696], addr_1674_6);

wire[27:0] addr_1675_6;

Selector_2 s1675_6(wires_418_5[3], addr_418_5, addr_positional[6703:6700], addr_1675_6);

wire[27:0] addr_1676_6;

Selector_2 s1676_6(wires_419_5[0], addr_419_5, addr_positional[6707:6704], addr_1676_6);

wire[27:0] addr_1677_6;

Selector_2 s1677_6(wires_419_5[1], addr_419_5, addr_positional[6711:6708], addr_1677_6);

wire[27:0] addr_1678_6;

Selector_2 s1678_6(wires_419_5[2], addr_419_5, addr_positional[6715:6712], addr_1678_6);

wire[27:0] addr_1679_6;

Selector_2 s1679_6(wires_419_5[3], addr_419_5, addr_positional[6719:6716], addr_1679_6);

wire[27:0] addr_1680_6;

Selector_2 s1680_6(wires_420_5[0], addr_420_5, addr_positional[6723:6720], addr_1680_6);

wire[27:0] addr_1681_6;

Selector_2 s1681_6(wires_420_5[1], addr_420_5, addr_positional[6727:6724], addr_1681_6);

wire[27:0] addr_1682_6;

Selector_2 s1682_6(wires_420_5[2], addr_420_5, addr_positional[6731:6728], addr_1682_6);

wire[27:0] addr_1683_6;

Selector_2 s1683_6(wires_420_5[3], addr_420_5, addr_positional[6735:6732], addr_1683_6);

wire[27:0] addr_1684_6;

Selector_2 s1684_6(wires_421_5[0], addr_421_5, addr_positional[6739:6736], addr_1684_6);

wire[27:0] addr_1685_6;

Selector_2 s1685_6(wires_421_5[1], addr_421_5, addr_positional[6743:6740], addr_1685_6);

wire[27:0] addr_1686_6;

Selector_2 s1686_6(wires_421_5[2], addr_421_5, addr_positional[6747:6744], addr_1686_6);

wire[27:0] addr_1687_6;

Selector_2 s1687_6(wires_421_5[3], addr_421_5, addr_positional[6751:6748], addr_1687_6);

wire[27:0] addr_1688_6;

Selector_2 s1688_6(wires_422_5[0], addr_422_5, addr_positional[6755:6752], addr_1688_6);

wire[27:0] addr_1689_6;

Selector_2 s1689_6(wires_422_5[1], addr_422_5, addr_positional[6759:6756], addr_1689_6);

wire[27:0] addr_1690_6;

Selector_2 s1690_6(wires_422_5[2], addr_422_5, addr_positional[6763:6760], addr_1690_6);

wire[27:0] addr_1691_6;

Selector_2 s1691_6(wires_422_5[3], addr_422_5, addr_positional[6767:6764], addr_1691_6);

wire[27:0] addr_1692_6;

Selector_2 s1692_6(wires_423_5[0], addr_423_5, addr_positional[6771:6768], addr_1692_6);

wire[27:0] addr_1693_6;

Selector_2 s1693_6(wires_423_5[1], addr_423_5, addr_positional[6775:6772], addr_1693_6);

wire[27:0] addr_1694_6;

Selector_2 s1694_6(wires_423_5[2], addr_423_5, addr_positional[6779:6776], addr_1694_6);

wire[27:0] addr_1695_6;

Selector_2 s1695_6(wires_423_5[3], addr_423_5, addr_positional[6783:6780], addr_1695_6);

wire[27:0] addr_1696_6;

Selector_2 s1696_6(wires_424_5[0], addr_424_5, addr_positional[6787:6784], addr_1696_6);

wire[27:0] addr_1697_6;

Selector_2 s1697_6(wires_424_5[1], addr_424_5, addr_positional[6791:6788], addr_1697_6);

wire[27:0] addr_1698_6;

Selector_2 s1698_6(wires_424_5[2], addr_424_5, addr_positional[6795:6792], addr_1698_6);

wire[27:0] addr_1699_6;

Selector_2 s1699_6(wires_424_5[3], addr_424_5, addr_positional[6799:6796], addr_1699_6);

wire[27:0] addr_1700_6;

Selector_2 s1700_6(wires_425_5[0], addr_425_5, addr_positional[6803:6800], addr_1700_6);

wire[27:0] addr_1701_6;

Selector_2 s1701_6(wires_425_5[1], addr_425_5, addr_positional[6807:6804], addr_1701_6);

wire[27:0] addr_1702_6;

Selector_2 s1702_6(wires_425_5[2], addr_425_5, addr_positional[6811:6808], addr_1702_6);

wire[27:0] addr_1703_6;

Selector_2 s1703_6(wires_425_5[3], addr_425_5, addr_positional[6815:6812], addr_1703_6);

wire[27:0] addr_1704_6;

Selector_2 s1704_6(wires_426_5[0], addr_426_5, addr_positional[6819:6816], addr_1704_6);

wire[27:0] addr_1705_6;

Selector_2 s1705_6(wires_426_5[1], addr_426_5, addr_positional[6823:6820], addr_1705_6);

wire[27:0] addr_1706_6;

Selector_2 s1706_6(wires_426_5[2], addr_426_5, addr_positional[6827:6824], addr_1706_6);

wire[27:0] addr_1707_6;

Selector_2 s1707_6(wires_426_5[3], addr_426_5, addr_positional[6831:6828], addr_1707_6);

wire[27:0] addr_1708_6;

Selector_2 s1708_6(wires_427_5[0], addr_427_5, addr_positional[6835:6832], addr_1708_6);

wire[27:0] addr_1709_6;

Selector_2 s1709_6(wires_427_5[1], addr_427_5, addr_positional[6839:6836], addr_1709_6);

wire[27:0] addr_1710_6;

Selector_2 s1710_6(wires_427_5[2], addr_427_5, addr_positional[6843:6840], addr_1710_6);

wire[27:0] addr_1711_6;

Selector_2 s1711_6(wires_427_5[3], addr_427_5, addr_positional[6847:6844], addr_1711_6);

wire[27:0] addr_1712_6;

Selector_2 s1712_6(wires_428_5[0], addr_428_5, addr_positional[6851:6848], addr_1712_6);

wire[27:0] addr_1713_6;

Selector_2 s1713_6(wires_428_5[1], addr_428_5, addr_positional[6855:6852], addr_1713_6);

wire[27:0] addr_1714_6;

Selector_2 s1714_6(wires_428_5[2], addr_428_5, addr_positional[6859:6856], addr_1714_6);

wire[27:0] addr_1715_6;

Selector_2 s1715_6(wires_428_5[3], addr_428_5, addr_positional[6863:6860], addr_1715_6);

wire[27:0] addr_1716_6;

Selector_2 s1716_6(wires_429_5[0], addr_429_5, addr_positional[6867:6864], addr_1716_6);

wire[27:0] addr_1717_6;

Selector_2 s1717_6(wires_429_5[1], addr_429_5, addr_positional[6871:6868], addr_1717_6);

wire[27:0] addr_1718_6;

Selector_2 s1718_6(wires_429_5[2], addr_429_5, addr_positional[6875:6872], addr_1718_6);

wire[27:0] addr_1719_6;

Selector_2 s1719_6(wires_429_5[3], addr_429_5, addr_positional[6879:6876], addr_1719_6);

wire[27:0] addr_1720_6;

Selector_2 s1720_6(wires_430_5[0], addr_430_5, addr_positional[6883:6880], addr_1720_6);

wire[27:0] addr_1721_6;

Selector_2 s1721_6(wires_430_5[1], addr_430_5, addr_positional[6887:6884], addr_1721_6);

wire[27:0] addr_1722_6;

Selector_2 s1722_6(wires_430_5[2], addr_430_5, addr_positional[6891:6888], addr_1722_6);

wire[27:0] addr_1723_6;

Selector_2 s1723_6(wires_430_5[3], addr_430_5, addr_positional[6895:6892], addr_1723_6);

wire[27:0] addr_1724_6;

Selector_2 s1724_6(wires_431_5[0], addr_431_5, addr_positional[6899:6896], addr_1724_6);

wire[27:0] addr_1725_6;

Selector_2 s1725_6(wires_431_5[1], addr_431_5, addr_positional[6903:6900], addr_1725_6);

wire[27:0] addr_1726_6;

Selector_2 s1726_6(wires_431_5[2], addr_431_5, addr_positional[6907:6904], addr_1726_6);

wire[27:0] addr_1727_6;

Selector_2 s1727_6(wires_431_5[3], addr_431_5, addr_positional[6911:6908], addr_1727_6);

wire[27:0] addr_1728_6;

Selector_2 s1728_6(wires_432_5[0], addr_432_5, addr_positional[6915:6912], addr_1728_6);

wire[27:0] addr_1729_6;

Selector_2 s1729_6(wires_432_5[1], addr_432_5, addr_positional[6919:6916], addr_1729_6);

wire[27:0] addr_1730_6;

Selector_2 s1730_6(wires_432_5[2], addr_432_5, addr_positional[6923:6920], addr_1730_6);

wire[27:0] addr_1731_6;

Selector_2 s1731_6(wires_432_5[3], addr_432_5, addr_positional[6927:6924], addr_1731_6);

wire[27:0] addr_1732_6;

Selector_2 s1732_6(wires_433_5[0], addr_433_5, addr_positional[6931:6928], addr_1732_6);

wire[27:0] addr_1733_6;

Selector_2 s1733_6(wires_433_5[1], addr_433_5, addr_positional[6935:6932], addr_1733_6);

wire[27:0] addr_1734_6;

Selector_2 s1734_6(wires_433_5[2], addr_433_5, addr_positional[6939:6936], addr_1734_6);

wire[27:0] addr_1735_6;

Selector_2 s1735_6(wires_433_5[3], addr_433_5, addr_positional[6943:6940], addr_1735_6);

wire[27:0] addr_1736_6;

Selector_2 s1736_6(wires_434_5[0], addr_434_5, addr_positional[6947:6944], addr_1736_6);

wire[27:0] addr_1737_6;

Selector_2 s1737_6(wires_434_5[1], addr_434_5, addr_positional[6951:6948], addr_1737_6);

wire[27:0] addr_1738_6;

Selector_2 s1738_6(wires_434_5[2], addr_434_5, addr_positional[6955:6952], addr_1738_6);

wire[27:0] addr_1739_6;

Selector_2 s1739_6(wires_434_5[3], addr_434_5, addr_positional[6959:6956], addr_1739_6);

wire[27:0] addr_1740_6;

Selector_2 s1740_6(wires_435_5[0], addr_435_5, addr_positional[6963:6960], addr_1740_6);

wire[27:0] addr_1741_6;

Selector_2 s1741_6(wires_435_5[1], addr_435_5, addr_positional[6967:6964], addr_1741_6);

wire[27:0] addr_1742_6;

Selector_2 s1742_6(wires_435_5[2], addr_435_5, addr_positional[6971:6968], addr_1742_6);

wire[27:0] addr_1743_6;

Selector_2 s1743_6(wires_435_5[3], addr_435_5, addr_positional[6975:6972], addr_1743_6);

wire[27:0] addr_1744_6;

Selector_2 s1744_6(wires_436_5[0], addr_436_5, addr_positional[6979:6976], addr_1744_6);

wire[27:0] addr_1745_6;

Selector_2 s1745_6(wires_436_5[1], addr_436_5, addr_positional[6983:6980], addr_1745_6);

wire[27:0] addr_1746_6;

Selector_2 s1746_6(wires_436_5[2], addr_436_5, addr_positional[6987:6984], addr_1746_6);

wire[27:0] addr_1747_6;

Selector_2 s1747_6(wires_436_5[3], addr_436_5, addr_positional[6991:6988], addr_1747_6);

wire[27:0] addr_1748_6;

Selector_2 s1748_6(wires_437_5[0], addr_437_5, addr_positional[6995:6992], addr_1748_6);

wire[27:0] addr_1749_6;

Selector_2 s1749_6(wires_437_5[1], addr_437_5, addr_positional[6999:6996], addr_1749_6);

wire[27:0] addr_1750_6;

Selector_2 s1750_6(wires_437_5[2], addr_437_5, addr_positional[7003:7000], addr_1750_6);

wire[27:0] addr_1751_6;

Selector_2 s1751_6(wires_437_5[3], addr_437_5, addr_positional[7007:7004], addr_1751_6);

wire[27:0] addr_1752_6;

Selector_2 s1752_6(wires_438_5[0], addr_438_5, addr_positional[7011:7008], addr_1752_6);

wire[27:0] addr_1753_6;

Selector_2 s1753_6(wires_438_5[1], addr_438_5, addr_positional[7015:7012], addr_1753_6);

wire[27:0] addr_1754_6;

Selector_2 s1754_6(wires_438_5[2], addr_438_5, addr_positional[7019:7016], addr_1754_6);

wire[27:0] addr_1755_6;

Selector_2 s1755_6(wires_438_5[3], addr_438_5, addr_positional[7023:7020], addr_1755_6);

wire[27:0] addr_1756_6;

Selector_2 s1756_6(wires_439_5[0], addr_439_5, addr_positional[7027:7024], addr_1756_6);

wire[27:0] addr_1757_6;

Selector_2 s1757_6(wires_439_5[1], addr_439_5, addr_positional[7031:7028], addr_1757_6);

wire[27:0] addr_1758_6;

Selector_2 s1758_6(wires_439_5[2], addr_439_5, addr_positional[7035:7032], addr_1758_6);

wire[27:0] addr_1759_6;

Selector_2 s1759_6(wires_439_5[3], addr_439_5, addr_positional[7039:7036], addr_1759_6);

wire[27:0] addr_1760_6;

Selector_2 s1760_6(wires_440_5[0], addr_440_5, addr_positional[7043:7040], addr_1760_6);

wire[27:0] addr_1761_6;

Selector_2 s1761_6(wires_440_5[1], addr_440_5, addr_positional[7047:7044], addr_1761_6);

wire[27:0] addr_1762_6;

Selector_2 s1762_6(wires_440_5[2], addr_440_5, addr_positional[7051:7048], addr_1762_6);

wire[27:0] addr_1763_6;

Selector_2 s1763_6(wires_440_5[3], addr_440_5, addr_positional[7055:7052], addr_1763_6);

wire[27:0] addr_1764_6;

Selector_2 s1764_6(wires_441_5[0], addr_441_5, addr_positional[7059:7056], addr_1764_6);

wire[27:0] addr_1765_6;

Selector_2 s1765_6(wires_441_5[1], addr_441_5, addr_positional[7063:7060], addr_1765_6);

wire[27:0] addr_1766_6;

Selector_2 s1766_6(wires_441_5[2], addr_441_5, addr_positional[7067:7064], addr_1766_6);

wire[27:0] addr_1767_6;

Selector_2 s1767_6(wires_441_5[3], addr_441_5, addr_positional[7071:7068], addr_1767_6);

wire[27:0] addr_1768_6;

Selector_2 s1768_6(wires_442_5[0], addr_442_5, addr_positional[7075:7072], addr_1768_6);

wire[27:0] addr_1769_6;

Selector_2 s1769_6(wires_442_5[1], addr_442_5, addr_positional[7079:7076], addr_1769_6);

wire[27:0] addr_1770_6;

Selector_2 s1770_6(wires_442_5[2], addr_442_5, addr_positional[7083:7080], addr_1770_6);

wire[27:0] addr_1771_6;

Selector_2 s1771_6(wires_442_5[3], addr_442_5, addr_positional[7087:7084], addr_1771_6);

wire[27:0] addr_1772_6;

Selector_2 s1772_6(wires_443_5[0], addr_443_5, addr_positional[7091:7088], addr_1772_6);

wire[27:0] addr_1773_6;

Selector_2 s1773_6(wires_443_5[1], addr_443_5, addr_positional[7095:7092], addr_1773_6);

wire[27:0] addr_1774_6;

Selector_2 s1774_6(wires_443_5[2], addr_443_5, addr_positional[7099:7096], addr_1774_6);

wire[27:0] addr_1775_6;

Selector_2 s1775_6(wires_443_5[3], addr_443_5, addr_positional[7103:7100], addr_1775_6);

wire[27:0] addr_1776_6;

Selector_2 s1776_6(wires_444_5[0], addr_444_5, addr_positional[7107:7104], addr_1776_6);

wire[27:0] addr_1777_6;

Selector_2 s1777_6(wires_444_5[1], addr_444_5, addr_positional[7111:7108], addr_1777_6);

wire[27:0] addr_1778_6;

Selector_2 s1778_6(wires_444_5[2], addr_444_5, addr_positional[7115:7112], addr_1778_6);

wire[27:0] addr_1779_6;

Selector_2 s1779_6(wires_444_5[3], addr_444_5, addr_positional[7119:7116], addr_1779_6);

wire[27:0] addr_1780_6;

Selector_2 s1780_6(wires_445_5[0], addr_445_5, addr_positional[7123:7120], addr_1780_6);

wire[27:0] addr_1781_6;

Selector_2 s1781_6(wires_445_5[1], addr_445_5, addr_positional[7127:7124], addr_1781_6);

wire[27:0] addr_1782_6;

Selector_2 s1782_6(wires_445_5[2], addr_445_5, addr_positional[7131:7128], addr_1782_6);

wire[27:0] addr_1783_6;

Selector_2 s1783_6(wires_445_5[3], addr_445_5, addr_positional[7135:7132], addr_1783_6);

wire[27:0] addr_1784_6;

Selector_2 s1784_6(wires_446_5[0], addr_446_5, addr_positional[7139:7136], addr_1784_6);

wire[27:0] addr_1785_6;

Selector_2 s1785_6(wires_446_5[1], addr_446_5, addr_positional[7143:7140], addr_1785_6);

wire[27:0] addr_1786_6;

Selector_2 s1786_6(wires_446_5[2], addr_446_5, addr_positional[7147:7144], addr_1786_6);

wire[27:0] addr_1787_6;

Selector_2 s1787_6(wires_446_5[3], addr_446_5, addr_positional[7151:7148], addr_1787_6);

wire[27:0] addr_1788_6;

Selector_2 s1788_6(wires_447_5[0], addr_447_5, addr_positional[7155:7152], addr_1788_6);

wire[27:0] addr_1789_6;

Selector_2 s1789_6(wires_447_5[1], addr_447_5, addr_positional[7159:7156], addr_1789_6);

wire[27:0] addr_1790_6;

Selector_2 s1790_6(wires_447_5[2], addr_447_5, addr_positional[7163:7160], addr_1790_6);

wire[27:0] addr_1791_6;

Selector_2 s1791_6(wires_447_5[3], addr_447_5, addr_positional[7167:7164], addr_1791_6);

wire[27:0] addr_1792_6;

Selector_2 s1792_6(wires_448_5[0], addr_448_5, addr_positional[7171:7168], addr_1792_6);

wire[27:0] addr_1793_6;

Selector_2 s1793_6(wires_448_5[1], addr_448_5, addr_positional[7175:7172], addr_1793_6);

wire[27:0] addr_1794_6;

Selector_2 s1794_6(wires_448_5[2], addr_448_5, addr_positional[7179:7176], addr_1794_6);

wire[27:0] addr_1795_6;

Selector_2 s1795_6(wires_448_5[3], addr_448_5, addr_positional[7183:7180], addr_1795_6);

wire[27:0] addr_1796_6;

Selector_2 s1796_6(wires_449_5[0], addr_449_5, addr_positional[7187:7184], addr_1796_6);

wire[27:0] addr_1797_6;

Selector_2 s1797_6(wires_449_5[1], addr_449_5, addr_positional[7191:7188], addr_1797_6);

wire[27:0] addr_1798_6;

Selector_2 s1798_6(wires_449_5[2], addr_449_5, addr_positional[7195:7192], addr_1798_6);

wire[27:0] addr_1799_6;

Selector_2 s1799_6(wires_449_5[3], addr_449_5, addr_positional[7199:7196], addr_1799_6);

wire[27:0] addr_1800_6;

Selector_2 s1800_6(wires_450_5[0], addr_450_5, addr_positional[7203:7200], addr_1800_6);

wire[27:0] addr_1801_6;

Selector_2 s1801_6(wires_450_5[1], addr_450_5, addr_positional[7207:7204], addr_1801_6);

wire[27:0] addr_1802_6;

Selector_2 s1802_6(wires_450_5[2], addr_450_5, addr_positional[7211:7208], addr_1802_6);

wire[27:0] addr_1803_6;

Selector_2 s1803_6(wires_450_5[3], addr_450_5, addr_positional[7215:7212], addr_1803_6);

wire[27:0] addr_1804_6;

Selector_2 s1804_6(wires_451_5[0], addr_451_5, addr_positional[7219:7216], addr_1804_6);

wire[27:0] addr_1805_6;

Selector_2 s1805_6(wires_451_5[1], addr_451_5, addr_positional[7223:7220], addr_1805_6);

wire[27:0] addr_1806_6;

Selector_2 s1806_6(wires_451_5[2], addr_451_5, addr_positional[7227:7224], addr_1806_6);

wire[27:0] addr_1807_6;

Selector_2 s1807_6(wires_451_5[3], addr_451_5, addr_positional[7231:7228], addr_1807_6);

wire[27:0] addr_1808_6;

Selector_2 s1808_6(wires_452_5[0], addr_452_5, addr_positional[7235:7232], addr_1808_6);

wire[27:0] addr_1809_6;

Selector_2 s1809_6(wires_452_5[1], addr_452_5, addr_positional[7239:7236], addr_1809_6);

wire[27:0] addr_1810_6;

Selector_2 s1810_6(wires_452_5[2], addr_452_5, addr_positional[7243:7240], addr_1810_6);

wire[27:0] addr_1811_6;

Selector_2 s1811_6(wires_452_5[3], addr_452_5, addr_positional[7247:7244], addr_1811_6);

wire[27:0] addr_1812_6;

Selector_2 s1812_6(wires_453_5[0], addr_453_5, addr_positional[7251:7248], addr_1812_6);

wire[27:0] addr_1813_6;

Selector_2 s1813_6(wires_453_5[1], addr_453_5, addr_positional[7255:7252], addr_1813_6);

wire[27:0] addr_1814_6;

Selector_2 s1814_6(wires_453_5[2], addr_453_5, addr_positional[7259:7256], addr_1814_6);

wire[27:0] addr_1815_6;

Selector_2 s1815_6(wires_453_5[3], addr_453_5, addr_positional[7263:7260], addr_1815_6);

wire[27:0] addr_1816_6;

Selector_2 s1816_6(wires_454_5[0], addr_454_5, addr_positional[7267:7264], addr_1816_6);

wire[27:0] addr_1817_6;

Selector_2 s1817_6(wires_454_5[1], addr_454_5, addr_positional[7271:7268], addr_1817_6);

wire[27:0] addr_1818_6;

Selector_2 s1818_6(wires_454_5[2], addr_454_5, addr_positional[7275:7272], addr_1818_6);

wire[27:0] addr_1819_6;

Selector_2 s1819_6(wires_454_5[3], addr_454_5, addr_positional[7279:7276], addr_1819_6);

wire[27:0] addr_1820_6;

Selector_2 s1820_6(wires_455_5[0], addr_455_5, addr_positional[7283:7280], addr_1820_6);

wire[27:0] addr_1821_6;

Selector_2 s1821_6(wires_455_5[1], addr_455_5, addr_positional[7287:7284], addr_1821_6);

wire[27:0] addr_1822_6;

Selector_2 s1822_6(wires_455_5[2], addr_455_5, addr_positional[7291:7288], addr_1822_6);

wire[27:0] addr_1823_6;

Selector_2 s1823_6(wires_455_5[3], addr_455_5, addr_positional[7295:7292], addr_1823_6);

wire[27:0] addr_1824_6;

Selector_2 s1824_6(wires_456_5[0], addr_456_5, addr_positional[7299:7296], addr_1824_6);

wire[27:0] addr_1825_6;

Selector_2 s1825_6(wires_456_5[1], addr_456_5, addr_positional[7303:7300], addr_1825_6);

wire[27:0] addr_1826_6;

Selector_2 s1826_6(wires_456_5[2], addr_456_5, addr_positional[7307:7304], addr_1826_6);

wire[27:0] addr_1827_6;

Selector_2 s1827_6(wires_456_5[3], addr_456_5, addr_positional[7311:7308], addr_1827_6);

wire[27:0] addr_1828_6;

Selector_2 s1828_6(wires_457_5[0], addr_457_5, addr_positional[7315:7312], addr_1828_6);

wire[27:0] addr_1829_6;

Selector_2 s1829_6(wires_457_5[1], addr_457_5, addr_positional[7319:7316], addr_1829_6);

wire[27:0] addr_1830_6;

Selector_2 s1830_6(wires_457_5[2], addr_457_5, addr_positional[7323:7320], addr_1830_6);

wire[27:0] addr_1831_6;

Selector_2 s1831_6(wires_457_5[3], addr_457_5, addr_positional[7327:7324], addr_1831_6);

wire[27:0] addr_1832_6;

Selector_2 s1832_6(wires_458_5[0], addr_458_5, addr_positional[7331:7328], addr_1832_6);

wire[27:0] addr_1833_6;

Selector_2 s1833_6(wires_458_5[1], addr_458_5, addr_positional[7335:7332], addr_1833_6);

wire[27:0] addr_1834_6;

Selector_2 s1834_6(wires_458_5[2], addr_458_5, addr_positional[7339:7336], addr_1834_6);

wire[27:0] addr_1835_6;

Selector_2 s1835_6(wires_458_5[3], addr_458_5, addr_positional[7343:7340], addr_1835_6);

wire[27:0] addr_1836_6;

Selector_2 s1836_6(wires_459_5[0], addr_459_5, addr_positional[7347:7344], addr_1836_6);

wire[27:0] addr_1837_6;

Selector_2 s1837_6(wires_459_5[1], addr_459_5, addr_positional[7351:7348], addr_1837_6);

wire[27:0] addr_1838_6;

Selector_2 s1838_6(wires_459_5[2], addr_459_5, addr_positional[7355:7352], addr_1838_6);

wire[27:0] addr_1839_6;

Selector_2 s1839_6(wires_459_5[3], addr_459_5, addr_positional[7359:7356], addr_1839_6);

wire[27:0] addr_1840_6;

Selector_2 s1840_6(wires_460_5[0], addr_460_5, addr_positional[7363:7360], addr_1840_6);

wire[27:0] addr_1841_6;

Selector_2 s1841_6(wires_460_5[1], addr_460_5, addr_positional[7367:7364], addr_1841_6);

wire[27:0] addr_1842_6;

Selector_2 s1842_6(wires_460_5[2], addr_460_5, addr_positional[7371:7368], addr_1842_6);

wire[27:0] addr_1843_6;

Selector_2 s1843_6(wires_460_5[3], addr_460_5, addr_positional[7375:7372], addr_1843_6);

wire[27:0] addr_1844_6;

Selector_2 s1844_6(wires_461_5[0], addr_461_5, addr_positional[7379:7376], addr_1844_6);

wire[27:0] addr_1845_6;

Selector_2 s1845_6(wires_461_5[1], addr_461_5, addr_positional[7383:7380], addr_1845_6);

wire[27:0] addr_1846_6;

Selector_2 s1846_6(wires_461_5[2], addr_461_5, addr_positional[7387:7384], addr_1846_6);

wire[27:0] addr_1847_6;

Selector_2 s1847_6(wires_461_5[3], addr_461_5, addr_positional[7391:7388], addr_1847_6);

wire[27:0] addr_1848_6;

Selector_2 s1848_6(wires_462_5[0], addr_462_5, addr_positional[7395:7392], addr_1848_6);

wire[27:0] addr_1849_6;

Selector_2 s1849_6(wires_462_5[1], addr_462_5, addr_positional[7399:7396], addr_1849_6);

wire[27:0] addr_1850_6;

Selector_2 s1850_6(wires_462_5[2], addr_462_5, addr_positional[7403:7400], addr_1850_6);

wire[27:0] addr_1851_6;

Selector_2 s1851_6(wires_462_5[3], addr_462_5, addr_positional[7407:7404], addr_1851_6);

wire[27:0] addr_1852_6;

Selector_2 s1852_6(wires_463_5[0], addr_463_5, addr_positional[7411:7408], addr_1852_6);

wire[27:0] addr_1853_6;

Selector_2 s1853_6(wires_463_5[1], addr_463_5, addr_positional[7415:7412], addr_1853_6);

wire[27:0] addr_1854_6;

Selector_2 s1854_6(wires_463_5[2], addr_463_5, addr_positional[7419:7416], addr_1854_6);

wire[27:0] addr_1855_6;

Selector_2 s1855_6(wires_463_5[3], addr_463_5, addr_positional[7423:7420], addr_1855_6);

wire[27:0] addr_1856_6;

Selector_2 s1856_6(wires_464_5[0], addr_464_5, addr_positional[7427:7424], addr_1856_6);

wire[27:0] addr_1857_6;

Selector_2 s1857_6(wires_464_5[1], addr_464_5, addr_positional[7431:7428], addr_1857_6);

wire[27:0] addr_1858_6;

Selector_2 s1858_6(wires_464_5[2], addr_464_5, addr_positional[7435:7432], addr_1858_6);

wire[27:0] addr_1859_6;

Selector_2 s1859_6(wires_464_5[3], addr_464_5, addr_positional[7439:7436], addr_1859_6);

wire[27:0] addr_1860_6;

Selector_2 s1860_6(wires_465_5[0], addr_465_5, addr_positional[7443:7440], addr_1860_6);

wire[27:0] addr_1861_6;

Selector_2 s1861_6(wires_465_5[1], addr_465_5, addr_positional[7447:7444], addr_1861_6);

wire[27:0] addr_1862_6;

Selector_2 s1862_6(wires_465_5[2], addr_465_5, addr_positional[7451:7448], addr_1862_6);

wire[27:0] addr_1863_6;

Selector_2 s1863_6(wires_465_5[3], addr_465_5, addr_positional[7455:7452], addr_1863_6);

wire[27:0] addr_1864_6;

Selector_2 s1864_6(wires_466_5[0], addr_466_5, addr_positional[7459:7456], addr_1864_6);

wire[27:0] addr_1865_6;

Selector_2 s1865_6(wires_466_5[1], addr_466_5, addr_positional[7463:7460], addr_1865_6);

wire[27:0] addr_1866_6;

Selector_2 s1866_6(wires_466_5[2], addr_466_5, addr_positional[7467:7464], addr_1866_6);

wire[27:0] addr_1867_6;

Selector_2 s1867_6(wires_466_5[3], addr_466_5, addr_positional[7471:7468], addr_1867_6);

wire[27:0] addr_1868_6;

Selector_2 s1868_6(wires_467_5[0], addr_467_5, addr_positional[7475:7472], addr_1868_6);

wire[27:0] addr_1869_6;

Selector_2 s1869_6(wires_467_5[1], addr_467_5, addr_positional[7479:7476], addr_1869_6);

wire[27:0] addr_1870_6;

Selector_2 s1870_6(wires_467_5[2], addr_467_5, addr_positional[7483:7480], addr_1870_6);

wire[27:0] addr_1871_6;

Selector_2 s1871_6(wires_467_5[3], addr_467_5, addr_positional[7487:7484], addr_1871_6);

wire[27:0] addr_1872_6;

Selector_2 s1872_6(wires_468_5[0], addr_468_5, addr_positional[7491:7488], addr_1872_6);

wire[27:0] addr_1873_6;

Selector_2 s1873_6(wires_468_5[1], addr_468_5, addr_positional[7495:7492], addr_1873_6);

wire[27:0] addr_1874_6;

Selector_2 s1874_6(wires_468_5[2], addr_468_5, addr_positional[7499:7496], addr_1874_6);

wire[27:0] addr_1875_6;

Selector_2 s1875_6(wires_468_5[3], addr_468_5, addr_positional[7503:7500], addr_1875_6);

wire[27:0] addr_1876_6;

Selector_2 s1876_6(wires_469_5[0], addr_469_5, addr_positional[7507:7504], addr_1876_6);

wire[27:0] addr_1877_6;

Selector_2 s1877_6(wires_469_5[1], addr_469_5, addr_positional[7511:7508], addr_1877_6);

wire[27:0] addr_1878_6;

Selector_2 s1878_6(wires_469_5[2], addr_469_5, addr_positional[7515:7512], addr_1878_6);

wire[27:0] addr_1879_6;

Selector_2 s1879_6(wires_469_5[3], addr_469_5, addr_positional[7519:7516], addr_1879_6);

wire[27:0] addr_1880_6;

Selector_2 s1880_6(wires_470_5[0], addr_470_5, addr_positional[7523:7520], addr_1880_6);

wire[27:0] addr_1881_6;

Selector_2 s1881_6(wires_470_5[1], addr_470_5, addr_positional[7527:7524], addr_1881_6);

wire[27:0] addr_1882_6;

Selector_2 s1882_6(wires_470_5[2], addr_470_5, addr_positional[7531:7528], addr_1882_6);

wire[27:0] addr_1883_6;

Selector_2 s1883_6(wires_470_5[3], addr_470_5, addr_positional[7535:7532], addr_1883_6);

wire[27:0] addr_1884_6;

Selector_2 s1884_6(wires_471_5[0], addr_471_5, addr_positional[7539:7536], addr_1884_6);

wire[27:0] addr_1885_6;

Selector_2 s1885_6(wires_471_5[1], addr_471_5, addr_positional[7543:7540], addr_1885_6);

wire[27:0] addr_1886_6;

Selector_2 s1886_6(wires_471_5[2], addr_471_5, addr_positional[7547:7544], addr_1886_6);

wire[27:0] addr_1887_6;

Selector_2 s1887_6(wires_471_5[3], addr_471_5, addr_positional[7551:7548], addr_1887_6);

wire[27:0] addr_1888_6;

Selector_2 s1888_6(wires_472_5[0], addr_472_5, addr_positional[7555:7552], addr_1888_6);

wire[27:0] addr_1889_6;

Selector_2 s1889_6(wires_472_5[1], addr_472_5, addr_positional[7559:7556], addr_1889_6);

wire[27:0] addr_1890_6;

Selector_2 s1890_6(wires_472_5[2], addr_472_5, addr_positional[7563:7560], addr_1890_6);

wire[27:0] addr_1891_6;

Selector_2 s1891_6(wires_472_5[3], addr_472_5, addr_positional[7567:7564], addr_1891_6);

wire[27:0] addr_1892_6;

Selector_2 s1892_6(wires_473_5[0], addr_473_5, addr_positional[7571:7568], addr_1892_6);

wire[27:0] addr_1893_6;

Selector_2 s1893_6(wires_473_5[1], addr_473_5, addr_positional[7575:7572], addr_1893_6);

wire[27:0] addr_1894_6;

Selector_2 s1894_6(wires_473_5[2], addr_473_5, addr_positional[7579:7576], addr_1894_6);

wire[27:0] addr_1895_6;

Selector_2 s1895_6(wires_473_5[3], addr_473_5, addr_positional[7583:7580], addr_1895_6);

wire[27:0] addr_1896_6;

Selector_2 s1896_6(wires_474_5[0], addr_474_5, addr_positional[7587:7584], addr_1896_6);

wire[27:0] addr_1897_6;

Selector_2 s1897_6(wires_474_5[1], addr_474_5, addr_positional[7591:7588], addr_1897_6);

wire[27:0] addr_1898_6;

Selector_2 s1898_6(wires_474_5[2], addr_474_5, addr_positional[7595:7592], addr_1898_6);

wire[27:0] addr_1899_6;

Selector_2 s1899_6(wires_474_5[3], addr_474_5, addr_positional[7599:7596], addr_1899_6);

wire[27:0] addr_1900_6;

Selector_2 s1900_6(wires_475_5[0], addr_475_5, addr_positional[7603:7600], addr_1900_6);

wire[27:0] addr_1901_6;

Selector_2 s1901_6(wires_475_5[1], addr_475_5, addr_positional[7607:7604], addr_1901_6);

wire[27:0] addr_1902_6;

Selector_2 s1902_6(wires_475_5[2], addr_475_5, addr_positional[7611:7608], addr_1902_6);

wire[27:0] addr_1903_6;

Selector_2 s1903_6(wires_475_5[3], addr_475_5, addr_positional[7615:7612], addr_1903_6);

wire[27:0] addr_1904_6;

Selector_2 s1904_6(wires_476_5[0], addr_476_5, addr_positional[7619:7616], addr_1904_6);

wire[27:0] addr_1905_6;

Selector_2 s1905_6(wires_476_5[1], addr_476_5, addr_positional[7623:7620], addr_1905_6);

wire[27:0] addr_1906_6;

Selector_2 s1906_6(wires_476_5[2], addr_476_5, addr_positional[7627:7624], addr_1906_6);

wire[27:0] addr_1907_6;

Selector_2 s1907_6(wires_476_5[3], addr_476_5, addr_positional[7631:7628], addr_1907_6);

wire[27:0] addr_1908_6;

Selector_2 s1908_6(wires_477_5[0], addr_477_5, addr_positional[7635:7632], addr_1908_6);

wire[27:0] addr_1909_6;

Selector_2 s1909_6(wires_477_5[1], addr_477_5, addr_positional[7639:7636], addr_1909_6);

wire[27:0] addr_1910_6;

Selector_2 s1910_6(wires_477_5[2], addr_477_5, addr_positional[7643:7640], addr_1910_6);

wire[27:0] addr_1911_6;

Selector_2 s1911_6(wires_477_5[3], addr_477_5, addr_positional[7647:7644], addr_1911_6);

wire[27:0] addr_1912_6;

Selector_2 s1912_6(wires_478_5[0], addr_478_5, addr_positional[7651:7648], addr_1912_6);

wire[27:0] addr_1913_6;

Selector_2 s1913_6(wires_478_5[1], addr_478_5, addr_positional[7655:7652], addr_1913_6);

wire[27:0] addr_1914_6;

Selector_2 s1914_6(wires_478_5[2], addr_478_5, addr_positional[7659:7656], addr_1914_6);

wire[27:0] addr_1915_6;

Selector_2 s1915_6(wires_478_5[3], addr_478_5, addr_positional[7663:7660], addr_1915_6);

wire[27:0] addr_1916_6;

Selector_2 s1916_6(wires_479_5[0], addr_479_5, addr_positional[7667:7664], addr_1916_6);

wire[27:0] addr_1917_6;

Selector_2 s1917_6(wires_479_5[1], addr_479_5, addr_positional[7671:7668], addr_1917_6);

wire[27:0] addr_1918_6;

Selector_2 s1918_6(wires_479_5[2], addr_479_5, addr_positional[7675:7672], addr_1918_6);

wire[27:0] addr_1919_6;

Selector_2 s1919_6(wires_479_5[3], addr_479_5, addr_positional[7679:7676], addr_1919_6);

wire[27:0] addr_1920_6;

Selector_2 s1920_6(wires_480_5[0], addr_480_5, addr_positional[7683:7680], addr_1920_6);

wire[27:0] addr_1921_6;

Selector_2 s1921_6(wires_480_5[1], addr_480_5, addr_positional[7687:7684], addr_1921_6);

wire[27:0] addr_1922_6;

Selector_2 s1922_6(wires_480_5[2], addr_480_5, addr_positional[7691:7688], addr_1922_6);

wire[27:0] addr_1923_6;

Selector_2 s1923_6(wires_480_5[3], addr_480_5, addr_positional[7695:7692], addr_1923_6);

wire[27:0] addr_1924_6;

Selector_2 s1924_6(wires_481_5[0], addr_481_5, addr_positional[7699:7696], addr_1924_6);

wire[27:0] addr_1925_6;

Selector_2 s1925_6(wires_481_5[1], addr_481_5, addr_positional[7703:7700], addr_1925_6);

wire[27:0] addr_1926_6;

Selector_2 s1926_6(wires_481_5[2], addr_481_5, addr_positional[7707:7704], addr_1926_6);

wire[27:0] addr_1927_6;

Selector_2 s1927_6(wires_481_5[3], addr_481_5, addr_positional[7711:7708], addr_1927_6);

wire[27:0] addr_1928_6;

Selector_2 s1928_6(wires_482_5[0], addr_482_5, addr_positional[7715:7712], addr_1928_6);

wire[27:0] addr_1929_6;

Selector_2 s1929_6(wires_482_5[1], addr_482_5, addr_positional[7719:7716], addr_1929_6);

wire[27:0] addr_1930_6;

Selector_2 s1930_6(wires_482_5[2], addr_482_5, addr_positional[7723:7720], addr_1930_6);

wire[27:0] addr_1931_6;

Selector_2 s1931_6(wires_482_5[3], addr_482_5, addr_positional[7727:7724], addr_1931_6);

wire[27:0] addr_1932_6;

Selector_2 s1932_6(wires_483_5[0], addr_483_5, addr_positional[7731:7728], addr_1932_6);

wire[27:0] addr_1933_6;

Selector_2 s1933_6(wires_483_5[1], addr_483_5, addr_positional[7735:7732], addr_1933_6);

wire[27:0] addr_1934_6;

Selector_2 s1934_6(wires_483_5[2], addr_483_5, addr_positional[7739:7736], addr_1934_6);

wire[27:0] addr_1935_6;

Selector_2 s1935_6(wires_483_5[3], addr_483_5, addr_positional[7743:7740], addr_1935_6);

wire[27:0] addr_1936_6;

Selector_2 s1936_6(wires_484_5[0], addr_484_5, addr_positional[7747:7744], addr_1936_6);

wire[27:0] addr_1937_6;

Selector_2 s1937_6(wires_484_5[1], addr_484_5, addr_positional[7751:7748], addr_1937_6);

wire[27:0] addr_1938_6;

Selector_2 s1938_6(wires_484_5[2], addr_484_5, addr_positional[7755:7752], addr_1938_6);

wire[27:0] addr_1939_6;

Selector_2 s1939_6(wires_484_5[3], addr_484_5, addr_positional[7759:7756], addr_1939_6);

wire[27:0] addr_1940_6;

Selector_2 s1940_6(wires_485_5[0], addr_485_5, addr_positional[7763:7760], addr_1940_6);

wire[27:0] addr_1941_6;

Selector_2 s1941_6(wires_485_5[1], addr_485_5, addr_positional[7767:7764], addr_1941_6);

wire[27:0] addr_1942_6;

Selector_2 s1942_6(wires_485_5[2], addr_485_5, addr_positional[7771:7768], addr_1942_6);

wire[27:0] addr_1943_6;

Selector_2 s1943_6(wires_485_5[3], addr_485_5, addr_positional[7775:7772], addr_1943_6);

wire[27:0] addr_1944_6;

Selector_2 s1944_6(wires_486_5[0], addr_486_5, addr_positional[7779:7776], addr_1944_6);

wire[27:0] addr_1945_6;

Selector_2 s1945_6(wires_486_5[1], addr_486_5, addr_positional[7783:7780], addr_1945_6);

wire[27:0] addr_1946_6;

Selector_2 s1946_6(wires_486_5[2], addr_486_5, addr_positional[7787:7784], addr_1946_6);

wire[27:0] addr_1947_6;

Selector_2 s1947_6(wires_486_5[3], addr_486_5, addr_positional[7791:7788], addr_1947_6);

wire[27:0] addr_1948_6;

Selector_2 s1948_6(wires_487_5[0], addr_487_5, addr_positional[7795:7792], addr_1948_6);

wire[27:0] addr_1949_6;

Selector_2 s1949_6(wires_487_5[1], addr_487_5, addr_positional[7799:7796], addr_1949_6);

wire[27:0] addr_1950_6;

Selector_2 s1950_6(wires_487_5[2], addr_487_5, addr_positional[7803:7800], addr_1950_6);

wire[27:0] addr_1951_6;

Selector_2 s1951_6(wires_487_5[3], addr_487_5, addr_positional[7807:7804], addr_1951_6);

wire[27:0] addr_1952_6;

Selector_2 s1952_6(wires_488_5[0], addr_488_5, addr_positional[7811:7808], addr_1952_6);

wire[27:0] addr_1953_6;

Selector_2 s1953_6(wires_488_5[1], addr_488_5, addr_positional[7815:7812], addr_1953_6);

wire[27:0] addr_1954_6;

Selector_2 s1954_6(wires_488_5[2], addr_488_5, addr_positional[7819:7816], addr_1954_6);

wire[27:0] addr_1955_6;

Selector_2 s1955_6(wires_488_5[3], addr_488_5, addr_positional[7823:7820], addr_1955_6);

wire[27:0] addr_1956_6;

Selector_2 s1956_6(wires_489_5[0], addr_489_5, addr_positional[7827:7824], addr_1956_6);

wire[27:0] addr_1957_6;

Selector_2 s1957_6(wires_489_5[1], addr_489_5, addr_positional[7831:7828], addr_1957_6);

wire[27:0] addr_1958_6;

Selector_2 s1958_6(wires_489_5[2], addr_489_5, addr_positional[7835:7832], addr_1958_6);

wire[27:0] addr_1959_6;

Selector_2 s1959_6(wires_489_5[3], addr_489_5, addr_positional[7839:7836], addr_1959_6);

wire[27:0] addr_1960_6;

Selector_2 s1960_6(wires_490_5[0], addr_490_5, addr_positional[7843:7840], addr_1960_6);

wire[27:0] addr_1961_6;

Selector_2 s1961_6(wires_490_5[1], addr_490_5, addr_positional[7847:7844], addr_1961_6);

wire[27:0] addr_1962_6;

Selector_2 s1962_6(wires_490_5[2], addr_490_5, addr_positional[7851:7848], addr_1962_6);

wire[27:0] addr_1963_6;

Selector_2 s1963_6(wires_490_5[3], addr_490_5, addr_positional[7855:7852], addr_1963_6);

wire[27:0] addr_1964_6;

Selector_2 s1964_6(wires_491_5[0], addr_491_5, addr_positional[7859:7856], addr_1964_6);

wire[27:0] addr_1965_6;

Selector_2 s1965_6(wires_491_5[1], addr_491_5, addr_positional[7863:7860], addr_1965_6);

wire[27:0] addr_1966_6;

Selector_2 s1966_6(wires_491_5[2], addr_491_5, addr_positional[7867:7864], addr_1966_6);

wire[27:0] addr_1967_6;

Selector_2 s1967_6(wires_491_5[3], addr_491_5, addr_positional[7871:7868], addr_1967_6);

wire[27:0] addr_1968_6;

Selector_2 s1968_6(wires_492_5[0], addr_492_5, addr_positional[7875:7872], addr_1968_6);

wire[27:0] addr_1969_6;

Selector_2 s1969_6(wires_492_5[1], addr_492_5, addr_positional[7879:7876], addr_1969_6);

wire[27:0] addr_1970_6;

Selector_2 s1970_6(wires_492_5[2], addr_492_5, addr_positional[7883:7880], addr_1970_6);

wire[27:0] addr_1971_6;

Selector_2 s1971_6(wires_492_5[3], addr_492_5, addr_positional[7887:7884], addr_1971_6);

wire[27:0] addr_1972_6;

Selector_2 s1972_6(wires_493_5[0], addr_493_5, addr_positional[7891:7888], addr_1972_6);

wire[27:0] addr_1973_6;

Selector_2 s1973_6(wires_493_5[1], addr_493_5, addr_positional[7895:7892], addr_1973_6);

wire[27:0] addr_1974_6;

Selector_2 s1974_6(wires_493_5[2], addr_493_5, addr_positional[7899:7896], addr_1974_6);

wire[27:0] addr_1975_6;

Selector_2 s1975_6(wires_493_5[3], addr_493_5, addr_positional[7903:7900], addr_1975_6);

wire[27:0] addr_1976_6;

Selector_2 s1976_6(wires_494_5[0], addr_494_5, addr_positional[7907:7904], addr_1976_6);

wire[27:0] addr_1977_6;

Selector_2 s1977_6(wires_494_5[1], addr_494_5, addr_positional[7911:7908], addr_1977_6);

wire[27:0] addr_1978_6;

Selector_2 s1978_6(wires_494_5[2], addr_494_5, addr_positional[7915:7912], addr_1978_6);

wire[27:0] addr_1979_6;

Selector_2 s1979_6(wires_494_5[3], addr_494_5, addr_positional[7919:7916], addr_1979_6);

wire[27:0] addr_1980_6;

Selector_2 s1980_6(wires_495_5[0], addr_495_5, addr_positional[7923:7920], addr_1980_6);

wire[27:0] addr_1981_6;

Selector_2 s1981_6(wires_495_5[1], addr_495_5, addr_positional[7927:7924], addr_1981_6);

wire[27:0] addr_1982_6;

Selector_2 s1982_6(wires_495_5[2], addr_495_5, addr_positional[7931:7928], addr_1982_6);

wire[27:0] addr_1983_6;

Selector_2 s1983_6(wires_495_5[3], addr_495_5, addr_positional[7935:7932], addr_1983_6);

wire[27:0] addr_1984_6;

Selector_2 s1984_6(wires_496_5[0], addr_496_5, addr_positional[7939:7936], addr_1984_6);

wire[27:0] addr_1985_6;

Selector_2 s1985_6(wires_496_5[1], addr_496_5, addr_positional[7943:7940], addr_1985_6);

wire[27:0] addr_1986_6;

Selector_2 s1986_6(wires_496_5[2], addr_496_5, addr_positional[7947:7944], addr_1986_6);

wire[27:0] addr_1987_6;

Selector_2 s1987_6(wires_496_5[3], addr_496_5, addr_positional[7951:7948], addr_1987_6);

wire[27:0] addr_1988_6;

Selector_2 s1988_6(wires_497_5[0], addr_497_5, addr_positional[7955:7952], addr_1988_6);

wire[27:0] addr_1989_6;

Selector_2 s1989_6(wires_497_5[1], addr_497_5, addr_positional[7959:7956], addr_1989_6);

wire[27:0] addr_1990_6;

Selector_2 s1990_6(wires_497_5[2], addr_497_5, addr_positional[7963:7960], addr_1990_6);

wire[27:0] addr_1991_6;

Selector_2 s1991_6(wires_497_5[3], addr_497_5, addr_positional[7967:7964], addr_1991_6);

wire[27:0] addr_1992_6;

Selector_2 s1992_6(wires_498_5[0], addr_498_5, addr_positional[7971:7968], addr_1992_6);

wire[27:0] addr_1993_6;

Selector_2 s1993_6(wires_498_5[1], addr_498_5, addr_positional[7975:7972], addr_1993_6);

wire[27:0] addr_1994_6;

Selector_2 s1994_6(wires_498_5[2], addr_498_5, addr_positional[7979:7976], addr_1994_6);

wire[27:0] addr_1995_6;

Selector_2 s1995_6(wires_498_5[3], addr_498_5, addr_positional[7983:7980], addr_1995_6);

wire[27:0] addr_1996_6;

Selector_2 s1996_6(wires_499_5[0], addr_499_5, addr_positional[7987:7984], addr_1996_6);

wire[27:0] addr_1997_6;

Selector_2 s1997_6(wires_499_5[1], addr_499_5, addr_positional[7991:7988], addr_1997_6);

wire[27:0] addr_1998_6;

Selector_2 s1998_6(wires_499_5[2], addr_499_5, addr_positional[7995:7992], addr_1998_6);

wire[27:0] addr_1999_6;

Selector_2 s1999_6(wires_499_5[3], addr_499_5, addr_positional[7999:7996], addr_1999_6);

wire[27:0] addr_2000_6;

Selector_2 s2000_6(wires_500_5[0], addr_500_5, addr_positional[8003:8000], addr_2000_6);

wire[27:0] addr_2001_6;

Selector_2 s2001_6(wires_500_5[1], addr_500_5, addr_positional[8007:8004], addr_2001_6);

wire[27:0] addr_2002_6;

Selector_2 s2002_6(wires_500_5[2], addr_500_5, addr_positional[8011:8008], addr_2002_6);

wire[27:0] addr_2003_6;

Selector_2 s2003_6(wires_500_5[3], addr_500_5, addr_positional[8015:8012], addr_2003_6);

wire[27:0] addr_2004_6;

Selector_2 s2004_6(wires_501_5[0], addr_501_5, addr_positional[8019:8016], addr_2004_6);

wire[27:0] addr_2005_6;

Selector_2 s2005_6(wires_501_5[1], addr_501_5, addr_positional[8023:8020], addr_2005_6);

wire[27:0] addr_2006_6;

Selector_2 s2006_6(wires_501_5[2], addr_501_5, addr_positional[8027:8024], addr_2006_6);

wire[27:0] addr_2007_6;

Selector_2 s2007_6(wires_501_5[3], addr_501_5, addr_positional[8031:8028], addr_2007_6);

wire[27:0] addr_2008_6;

Selector_2 s2008_6(wires_502_5[0], addr_502_5, addr_positional[8035:8032], addr_2008_6);

wire[27:0] addr_2009_6;

Selector_2 s2009_6(wires_502_5[1], addr_502_5, addr_positional[8039:8036], addr_2009_6);

wire[27:0] addr_2010_6;

Selector_2 s2010_6(wires_502_5[2], addr_502_5, addr_positional[8043:8040], addr_2010_6);

wire[27:0] addr_2011_6;

Selector_2 s2011_6(wires_502_5[3], addr_502_5, addr_positional[8047:8044], addr_2011_6);

wire[27:0] addr_2012_6;

Selector_2 s2012_6(wires_503_5[0], addr_503_5, addr_positional[8051:8048], addr_2012_6);

wire[27:0] addr_2013_6;

Selector_2 s2013_6(wires_503_5[1], addr_503_5, addr_positional[8055:8052], addr_2013_6);

wire[27:0] addr_2014_6;

Selector_2 s2014_6(wires_503_5[2], addr_503_5, addr_positional[8059:8056], addr_2014_6);

wire[27:0] addr_2015_6;

Selector_2 s2015_6(wires_503_5[3], addr_503_5, addr_positional[8063:8060], addr_2015_6);

wire[27:0] addr_2016_6;

Selector_2 s2016_6(wires_504_5[0], addr_504_5, addr_positional[8067:8064], addr_2016_6);

wire[27:0] addr_2017_6;

Selector_2 s2017_6(wires_504_5[1], addr_504_5, addr_positional[8071:8068], addr_2017_6);

wire[27:0] addr_2018_6;

Selector_2 s2018_6(wires_504_5[2], addr_504_5, addr_positional[8075:8072], addr_2018_6);

wire[27:0] addr_2019_6;

Selector_2 s2019_6(wires_504_5[3], addr_504_5, addr_positional[8079:8076], addr_2019_6);

wire[27:0] addr_2020_6;

Selector_2 s2020_6(wires_505_5[0], addr_505_5, addr_positional[8083:8080], addr_2020_6);

wire[27:0] addr_2021_6;

Selector_2 s2021_6(wires_505_5[1], addr_505_5, addr_positional[8087:8084], addr_2021_6);

wire[27:0] addr_2022_6;

Selector_2 s2022_6(wires_505_5[2], addr_505_5, addr_positional[8091:8088], addr_2022_6);

wire[27:0] addr_2023_6;

Selector_2 s2023_6(wires_505_5[3], addr_505_5, addr_positional[8095:8092], addr_2023_6);

wire[27:0] addr_2024_6;

Selector_2 s2024_6(wires_506_5[0], addr_506_5, addr_positional[8099:8096], addr_2024_6);

wire[27:0] addr_2025_6;

Selector_2 s2025_6(wires_506_5[1], addr_506_5, addr_positional[8103:8100], addr_2025_6);

wire[27:0] addr_2026_6;

Selector_2 s2026_6(wires_506_5[2], addr_506_5, addr_positional[8107:8104], addr_2026_6);

wire[27:0] addr_2027_6;

Selector_2 s2027_6(wires_506_5[3], addr_506_5, addr_positional[8111:8108], addr_2027_6);

wire[27:0] addr_2028_6;

Selector_2 s2028_6(wires_507_5[0], addr_507_5, addr_positional[8115:8112], addr_2028_6);

wire[27:0] addr_2029_6;

Selector_2 s2029_6(wires_507_5[1], addr_507_5, addr_positional[8119:8116], addr_2029_6);

wire[27:0] addr_2030_6;

Selector_2 s2030_6(wires_507_5[2], addr_507_5, addr_positional[8123:8120], addr_2030_6);

wire[27:0] addr_2031_6;

Selector_2 s2031_6(wires_507_5[3], addr_507_5, addr_positional[8127:8124], addr_2031_6);

wire[27:0] addr_2032_6;

Selector_2 s2032_6(wires_508_5[0], addr_508_5, addr_positional[8131:8128], addr_2032_6);

wire[27:0] addr_2033_6;

Selector_2 s2033_6(wires_508_5[1], addr_508_5, addr_positional[8135:8132], addr_2033_6);

wire[27:0] addr_2034_6;

Selector_2 s2034_6(wires_508_5[2], addr_508_5, addr_positional[8139:8136], addr_2034_6);

wire[27:0] addr_2035_6;

Selector_2 s2035_6(wires_508_5[3], addr_508_5, addr_positional[8143:8140], addr_2035_6);

wire[27:0] addr_2036_6;

Selector_2 s2036_6(wires_509_5[0], addr_509_5, addr_positional[8147:8144], addr_2036_6);

wire[27:0] addr_2037_6;

Selector_2 s2037_6(wires_509_5[1], addr_509_5, addr_positional[8151:8148], addr_2037_6);

wire[27:0] addr_2038_6;

Selector_2 s2038_6(wires_509_5[2], addr_509_5, addr_positional[8155:8152], addr_2038_6);

wire[27:0] addr_2039_6;

Selector_2 s2039_6(wires_509_5[3], addr_509_5, addr_positional[8159:8156], addr_2039_6);

wire[27:0] addr_2040_6;

Selector_2 s2040_6(wires_510_5[0], addr_510_5, addr_positional[8163:8160], addr_2040_6);

wire[27:0] addr_2041_6;

Selector_2 s2041_6(wires_510_5[1], addr_510_5, addr_positional[8167:8164], addr_2041_6);

wire[27:0] addr_2042_6;

Selector_2 s2042_6(wires_510_5[2], addr_510_5, addr_positional[8171:8168], addr_2042_6);

wire[27:0] addr_2043_6;

Selector_2 s2043_6(wires_510_5[3], addr_510_5, addr_positional[8175:8172], addr_2043_6);

wire[27:0] addr_2044_6;

Selector_2 s2044_6(wires_511_5[0], addr_511_5, addr_positional[8179:8176], addr_2044_6);

wire[27:0] addr_2045_6;

Selector_2 s2045_6(wires_511_5[1], addr_511_5, addr_positional[8183:8180], addr_2045_6);

wire[27:0] addr_2046_6;

Selector_2 s2046_6(wires_511_5[2], addr_511_5, addr_positional[8187:8184], addr_2046_6);

wire[27:0] addr_2047_6;

Selector_2 s2047_6(wires_511_5[3], addr_511_5, addr_positional[8191:8188], addr_2047_6);

wire[27:0] addr_2048_6;

Selector_2 s2048_6(wires_512_5[0], addr_512_5, addr_positional[8195:8192], addr_2048_6);

wire[27:0] addr_2049_6;

Selector_2 s2049_6(wires_512_5[1], addr_512_5, addr_positional[8199:8196], addr_2049_6);

wire[27:0] addr_2050_6;

Selector_2 s2050_6(wires_512_5[2], addr_512_5, addr_positional[8203:8200], addr_2050_6);

wire[27:0] addr_2051_6;

Selector_2 s2051_6(wires_512_5[3], addr_512_5, addr_positional[8207:8204], addr_2051_6);

wire[27:0] addr_2052_6;

Selector_2 s2052_6(wires_513_5[0], addr_513_5, addr_positional[8211:8208], addr_2052_6);

wire[27:0] addr_2053_6;

Selector_2 s2053_6(wires_513_5[1], addr_513_5, addr_positional[8215:8212], addr_2053_6);

wire[27:0] addr_2054_6;

Selector_2 s2054_6(wires_513_5[2], addr_513_5, addr_positional[8219:8216], addr_2054_6);

wire[27:0] addr_2055_6;

Selector_2 s2055_6(wires_513_5[3], addr_513_5, addr_positional[8223:8220], addr_2055_6);

wire[27:0] addr_2056_6;

Selector_2 s2056_6(wires_514_5[0], addr_514_5, addr_positional[8227:8224], addr_2056_6);

wire[27:0] addr_2057_6;

Selector_2 s2057_6(wires_514_5[1], addr_514_5, addr_positional[8231:8228], addr_2057_6);

wire[27:0] addr_2058_6;

Selector_2 s2058_6(wires_514_5[2], addr_514_5, addr_positional[8235:8232], addr_2058_6);

wire[27:0] addr_2059_6;

Selector_2 s2059_6(wires_514_5[3], addr_514_5, addr_positional[8239:8236], addr_2059_6);

wire[27:0] addr_2060_6;

Selector_2 s2060_6(wires_515_5[0], addr_515_5, addr_positional[8243:8240], addr_2060_6);

wire[27:0] addr_2061_6;

Selector_2 s2061_6(wires_515_5[1], addr_515_5, addr_positional[8247:8244], addr_2061_6);

wire[27:0] addr_2062_6;

Selector_2 s2062_6(wires_515_5[2], addr_515_5, addr_positional[8251:8248], addr_2062_6);

wire[27:0] addr_2063_6;

Selector_2 s2063_6(wires_515_5[3], addr_515_5, addr_positional[8255:8252], addr_2063_6);

wire[27:0] addr_2064_6;

Selector_2 s2064_6(wires_516_5[0], addr_516_5, addr_positional[8259:8256], addr_2064_6);

wire[27:0] addr_2065_6;

Selector_2 s2065_6(wires_516_5[1], addr_516_5, addr_positional[8263:8260], addr_2065_6);

wire[27:0] addr_2066_6;

Selector_2 s2066_6(wires_516_5[2], addr_516_5, addr_positional[8267:8264], addr_2066_6);

wire[27:0] addr_2067_6;

Selector_2 s2067_6(wires_516_5[3], addr_516_5, addr_positional[8271:8268], addr_2067_6);

wire[27:0] addr_2068_6;

Selector_2 s2068_6(wires_517_5[0], addr_517_5, addr_positional[8275:8272], addr_2068_6);

wire[27:0] addr_2069_6;

Selector_2 s2069_6(wires_517_5[1], addr_517_5, addr_positional[8279:8276], addr_2069_6);

wire[27:0] addr_2070_6;

Selector_2 s2070_6(wires_517_5[2], addr_517_5, addr_positional[8283:8280], addr_2070_6);

wire[27:0] addr_2071_6;

Selector_2 s2071_6(wires_517_5[3], addr_517_5, addr_positional[8287:8284], addr_2071_6);

wire[27:0] addr_2072_6;

Selector_2 s2072_6(wires_518_5[0], addr_518_5, addr_positional[8291:8288], addr_2072_6);

wire[27:0] addr_2073_6;

Selector_2 s2073_6(wires_518_5[1], addr_518_5, addr_positional[8295:8292], addr_2073_6);

wire[27:0] addr_2074_6;

Selector_2 s2074_6(wires_518_5[2], addr_518_5, addr_positional[8299:8296], addr_2074_6);

wire[27:0] addr_2075_6;

Selector_2 s2075_6(wires_518_5[3], addr_518_5, addr_positional[8303:8300], addr_2075_6);

wire[27:0] addr_2076_6;

Selector_2 s2076_6(wires_519_5[0], addr_519_5, addr_positional[8307:8304], addr_2076_6);

wire[27:0] addr_2077_6;

Selector_2 s2077_6(wires_519_5[1], addr_519_5, addr_positional[8311:8308], addr_2077_6);

wire[27:0] addr_2078_6;

Selector_2 s2078_6(wires_519_5[2], addr_519_5, addr_positional[8315:8312], addr_2078_6);

wire[27:0] addr_2079_6;

Selector_2 s2079_6(wires_519_5[3], addr_519_5, addr_positional[8319:8316], addr_2079_6);

wire[27:0] addr_2080_6;

Selector_2 s2080_6(wires_520_5[0], addr_520_5, addr_positional[8323:8320], addr_2080_6);

wire[27:0] addr_2081_6;

Selector_2 s2081_6(wires_520_5[1], addr_520_5, addr_positional[8327:8324], addr_2081_6);

wire[27:0] addr_2082_6;

Selector_2 s2082_6(wires_520_5[2], addr_520_5, addr_positional[8331:8328], addr_2082_6);

wire[27:0] addr_2083_6;

Selector_2 s2083_6(wires_520_5[3], addr_520_5, addr_positional[8335:8332], addr_2083_6);

wire[27:0] addr_2084_6;

Selector_2 s2084_6(wires_521_5[0], addr_521_5, addr_positional[8339:8336], addr_2084_6);

wire[27:0] addr_2085_6;

Selector_2 s2085_6(wires_521_5[1], addr_521_5, addr_positional[8343:8340], addr_2085_6);

wire[27:0] addr_2086_6;

Selector_2 s2086_6(wires_521_5[2], addr_521_5, addr_positional[8347:8344], addr_2086_6);

wire[27:0] addr_2087_6;

Selector_2 s2087_6(wires_521_5[3], addr_521_5, addr_positional[8351:8348], addr_2087_6);

wire[27:0] addr_2088_6;

Selector_2 s2088_6(wires_522_5[0], addr_522_5, addr_positional[8355:8352], addr_2088_6);

wire[27:0] addr_2089_6;

Selector_2 s2089_6(wires_522_5[1], addr_522_5, addr_positional[8359:8356], addr_2089_6);

wire[27:0] addr_2090_6;

Selector_2 s2090_6(wires_522_5[2], addr_522_5, addr_positional[8363:8360], addr_2090_6);

wire[27:0] addr_2091_6;

Selector_2 s2091_6(wires_522_5[3], addr_522_5, addr_positional[8367:8364], addr_2091_6);

wire[27:0] addr_2092_6;

Selector_2 s2092_6(wires_523_5[0], addr_523_5, addr_positional[8371:8368], addr_2092_6);

wire[27:0] addr_2093_6;

Selector_2 s2093_6(wires_523_5[1], addr_523_5, addr_positional[8375:8372], addr_2093_6);

wire[27:0] addr_2094_6;

Selector_2 s2094_6(wires_523_5[2], addr_523_5, addr_positional[8379:8376], addr_2094_6);

wire[27:0] addr_2095_6;

Selector_2 s2095_6(wires_523_5[3], addr_523_5, addr_positional[8383:8380], addr_2095_6);

wire[27:0] addr_2096_6;

Selector_2 s2096_6(wires_524_5[0], addr_524_5, addr_positional[8387:8384], addr_2096_6);

wire[27:0] addr_2097_6;

Selector_2 s2097_6(wires_524_5[1], addr_524_5, addr_positional[8391:8388], addr_2097_6);

wire[27:0] addr_2098_6;

Selector_2 s2098_6(wires_524_5[2], addr_524_5, addr_positional[8395:8392], addr_2098_6);

wire[27:0] addr_2099_6;

Selector_2 s2099_6(wires_524_5[3], addr_524_5, addr_positional[8399:8396], addr_2099_6);

wire[27:0] addr_2100_6;

Selector_2 s2100_6(wires_525_5[0], addr_525_5, addr_positional[8403:8400], addr_2100_6);

wire[27:0] addr_2101_6;

Selector_2 s2101_6(wires_525_5[1], addr_525_5, addr_positional[8407:8404], addr_2101_6);

wire[27:0] addr_2102_6;

Selector_2 s2102_6(wires_525_5[2], addr_525_5, addr_positional[8411:8408], addr_2102_6);

wire[27:0] addr_2103_6;

Selector_2 s2103_6(wires_525_5[3], addr_525_5, addr_positional[8415:8412], addr_2103_6);

wire[27:0] addr_2104_6;

Selector_2 s2104_6(wires_526_5[0], addr_526_5, addr_positional[8419:8416], addr_2104_6);

wire[27:0] addr_2105_6;

Selector_2 s2105_6(wires_526_5[1], addr_526_5, addr_positional[8423:8420], addr_2105_6);

wire[27:0] addr_2106_6;

Selector_2 s2106_6(wires_526_5[2], addr_526_5, addr_positional[8427:8424], addr_2106_6);

wire[27:0] addr_2107_6;

Selector_2 s2107_6(wires_526_5[3], addr_526_5, addr_positional[8431:8428], addr_2107_6);

wire[27:0] addr_2108_6;

Selector_2 s2108_6(wires_527_5[0], addr_527_5, addr_positional[8435:8432], addr_2108_6);

wire[27:0] addr_2109_6;

Selector_2 s2109_6(wires_527_5[1], addr_527_5, addr_positional[8439:8436], addr_2109_6);

wire[27:0] addr_2110_6;

Selector_2 s2110_6(wires_527_5[2], addr_527_5, addr_positional[8443:8440], addr_2110_6);

wire[27:0] addr_2111_6;

Selector_2 s2111_6(wires_527_5[3], addr_527_5, addr_positional[8447:8444], addr_2111_6);

wire[27:0] addr_2112_6;

Selector_2 s2112_6(wires_528_5[0], addr_528_5, addr_positional[8451:8448], addr_2112_6);

wire[27:0] addr_2113_6;

Selector_2 s2113_6(wires_528_5[1], addr_528_5, addr_positional[8455:8452], addr_2113_6);

wire[27:0] addr_2114_6;

Selector_2 s2114_6(wires_528_5[2], addr_528_5, addr_positional[8459:8456], addr_2114_6);

wire[27:0] addr_2115_6;

Selector_2 s2115_6(wires_528_5[3], addr_528_5, addr_positional[8463:8460], addr_2115_6);

wire[27:0] addr_2116_6;

Selector_2 s2116_6(wires_529_5[0], addr_529_5, addr_positional[8467:8464], addr_2116_6);

wire[27:0] addr_2117_6;

Selector_2 s2117_6(wires_529_5[1], addr_529_5, addr_positional[8471:8468], addr_2117_6);

wire[27:0] addr_2118_6;

Selector_2 s2118_6(wires_529_5[2], addr_529_5, addr_positional[8475:8472], addr_2118_6);

wire[27:0] addr_2119_6;

Selector_2 s2119_6(wires_529_5[3], addr_529_5, addr_positional[8479:8476], addr_2119_6);

wire[27:0] addr_2120_6;

Selector_2 s2120_6(wires_530_5[0], addr_530_5, addr_positional[8483:8480], addr_2120_6);

wire[27:0] addr_2121_6;

Selector_2 s2121_6(wires_530_5[1], addr_530_5, addr_positional[8487:8484], addr_2121_6);

wire[27:0] addr_2122_6;

Selector_2 s2122_6(wires_530_5[2], addr_530_5, addr_positional[8491:8488], addr_2122_6);

wire[27:0] addr_2123_6;

Selector_2 s2123_6(wires_530_5[3], addr_530_5, addr_positional[8495:8492], addr_2123_6);

wire[27:0] addr_2124_6;

Selector_2 s2124_6(wires_531_5[0], addr_531_5, addr_positional[8499:8496], addr_2124_6);

wire[27:0] addr_2125_6;

Selector_2 s2125_6(wires_531_5[1], addr_531_5, addr_positional[8503:8500], addr_2125_6);

wire[27:0] addr_2126_6;

Selector_2 s2126_6(wires_531_5[2], addr_531_5, addr_positional[8507:8504], addr_2126_6);

wire[27:0] addr_2127_6;

Selector_2 s2127_6(wires_531_5[3], addr_531_5, addr_positional[8511:8508], addr_2127_6);

wire[27:0] addr_2128_6;

Selector_2 s2128_6(wires_532_5[0], addr_532_5, addr_positional[8515:8512], addr_2128_6);

wire[27:0] addr_2129_6;

Selector_2 s2129_6(wires_532_5[1], addr_532_5, addr_positional[8519:8516], addr_2129_6);

wire[27:0] addr_2130_6;

Selector_2 s2130_6(wires_532_5[2], addr_532_5, addr_positional[8523:8520], addr_2130_6);

wire[27:0] addr_2131_6;

Selector_2 s2131_6(wires_532_5[3], addr_532_5, addr_positional[8527:8524], addr_2131_6);

wire[27:0] addr_2132_6;

Selector_2 s2132_6(wires_533_5[0], addr_533_5, addr_positional[8531:8528], addr_2132_6);

wire[27:0] addr_2133_6;

Selector_2 s2133_6(wires_533_5[1], addr_533_5, addr_positional[8535:8532], addr_2133_6);

wire[27:0] addr_2134_6;

Selector_2 s2134_6(wires_533_5[2], addr_533_5, addr_positional[8539:8536], addr_2134_6);

wire[27:0] addr_2135_6;

Selector_2 s2135_6(wires_533_5[3], addr_533_5, addr_positional[8543:8540], addr_2135_6);

wire[27:0] addr_2136_6;

Selector_2 s2136_6(wires_534_5[0], addr_534_5, addr_positional[8547:8544], addr_2136_6);

wire[27:0] addr_2137_6;

Selector_2 s2137_6(wires_534_5[1], addr_534_5, addr_positional[8551:8548], addr_2137_6);

wire[27:0] addr_2138_6;

Selector_2 s2138_6(wires_534_5[2], addr_534_5, addr_positional[8555:8552], addr_2138_6);

wire[27:0] addr_2139_6;

Selector_2 s2139_6(wires_534_5[3], addr_534_5, addr_positional[8559:8556], addr_2139_6);

wire[27:0] addr_2140_6;

Selector_2 s2140_6(wires_535_5[0], addr_535_5, addr_positional[8563:8560], addr_2140_6);

wire[27:0] addr_2141_6;

Selector_2 s2141_6(wires_535_5[1], addr_535_5, addr_positional[8567:8564], addr_2141_6);

wire[27:0] addr_2142_6;

Selector_2 s2142_6(wires_535_5[2], addr_535_5, addr_positional[8571:8568], addr_2142_6);

wire[27:0] addr_2143_6;

Selector_2 s2143_6(wires_535_5[3], addr_535_5, addr_positional[8575:8572], addr_2143_6);

wire[27:0] addr_2144_6;

Selector_2 s2144_6(wires_536_5[0], addr_536_5, addr_positional[8579:8576], addr_2144_6);

wire[27:0] addr_2145_6;

Selector_2 s2145_6(wires_536_5[1], addr_536_5, addr_positional[8583:8580], addr_2145_6);

wire[27:0] addr_2146_6;

Selector_2 s2146_6(wires_536_5[2], addr_536_5, addr_positional[8587:8584], addr_2146_6);

wire[27:0] addr_2147_6;

Selector_2 s2147_6(wires_536_5[3], addr_536_5, addr_positional[8591:8588], addr_2147_6);

wire[27:0] addr_2148_6;

Selector_2 s2148_6(wires_537_5[0], addr_537_5, addr_positional[8595:8592], addr_2148_6);

wire[27:0] addr_2149_6;

Selector_2 s2149_6(wires_537_5[1], addr_537_5, addr_positional[8599:8596], addr_2149_6);

wire[27:0] addr_2150_6;

Selector_2 s2150_6(wires_537_5[2], addr_537_5, addr_positional[8603:8600], addr_2150_6);

wire[27:0] addr_2151_6;

Selector_2 s2151_6(wires_537_5[3], addr_537_5, addr_positional[8607:8604], addr_2151_6);

wire[27:0] addr_2152_6;

Selector_2 s2152_6(wires_538_5[0], addr_538_5, addr_positional[8611:8608], addr_2152_6);

wire[27:0] addr_2153_6;

Selector_2 s2153_6(wires_538_5[1], addr_538_5, addr_positional[8615:8612], addr_2153_6);

wire[27:0] addr_2154_6;

Selector_2 s2154_6(wires_538_5[2], addr_538_5, addr_positional[8619:8616], addr_2154_6);

wire[27:0] addr_2155_6;

Selector_2 s2155_6(wires_538_5[3], addr_538_5, addr_positional[8623:8620], addr_2155_6);

wire[27:0] addr_2156_6;

Selector_2 s2156_6(wires_539_5[0], addr_539_5, addr_positional[8627:8624], addr_2156_6);

wire[27:0] addr_2157_6;

Selector_2 s2157_6(wires_539_5[1], addr_539_5, addr_positional[8631:8628], addr_2157_6);

wire[27:0] addr_2158_6;

Selector_2 s2158_6(wires_539_5[2], addr_539_5, addr_positional[8635:8632], addr_2158_6);

wire[27:0] addr_2159_6;

Selector_2 s2159_6(wires_539_5[3], addr_539_5, addr_positional[8639:8636], addr_2159_6);

wire[27:0] addr_2160_6;

Selector_2 s2160_6(wires_540_5[0], addr_540_5, addr_positional[8643:8640], addr_2160_6);

wire[27:0] addr_2161_6;

Selector_2 s2161_6(wires_540_5[1], addr_540_5, addr_positional[8647:8644], addr_2161_6);

wire[27:0] addr_2162_6;

Selector_2 s2162_6(wires_540_5[2], addr_540_5, addr_positional[8651:8648], addr_2162_6);

wire[27:0] addr_2163_6;

Selector_2 s2163_6(wires_540_5[3], addr_540_5, addr_positional[8655:8652], addr_2163_6);

wire[27:0] addr_2164_6;

Selector_2 s2164_6(wires_541_5[0], addr_541_5, addr_positional[8659:8656], addr_2164_6);

wire[27:0] addr_2165_6;

Selector_2 s2165_6(wires_541_5[1], addr_541_5, addr_positional[8663:8660], addr_2165_6);

wire[27:0] addr_2166_6;

Selector_2 s2166_6(wires_541_5[2], addr_541_5, addr_positional[8667:8664], addr_2166_6);

wire[27:0] addr_2167_6;

Selector_2 s2167_6(wires_541_5[3], addr_541_5, addr_positional[8671:8668], addr_2167_6);

wire[27:0] addr_2168_6;

Selector_2 s2168_6(wires_542_5[0], addr_542_5, addr_positional[8675:8672], addr_2168_6);

wire[27:0] addr_2169_6;

Selector_2 s2169_6(wires_542_5[1], addr_542_5, addr_positional[8679:8676], addr_2169_6);

wire[27:0] addr_2170_6;

Selector_2 s2170_6(wires_542_5[2], addr_542_5, addr_positional[8683:8680], addr_2170_6);

wire[27:0] addr_2171_6;

Selector_2 s2171_6(wires_542_5[3], addr_542_5, addr_positional[8687:8684], addr_2171_6);

wire[27:0] addr_2172_6;

Selector_2 s2172_6(wires_543_5[0], addr_543_5, addr_positional[8691:8688], addr_2172_6);

wire[27:0] addr_2173_6;

Selector_2 s2173_6(wires_543_5[1], addr_543_5, addr_positional[8695:8692], addr_2173_6);

wire[27:0] addr_2174_6;

Selector_2 s2174_6(wires_543_5[2], addr_543_5, addr_positional[8699:8696], addr_2174_6);

wire[27:0] addr_2175_6;

Selector_2 s2175_6(wires_543_5[3], addr_543_5, addr_positional[8703:8700], addr_2175_6);

wire[27:0] addr_2176_6;

Selector_2 s2176_6(wires_544_5[0], addr_544_5, addr_positional[8707:8704], addr_2176_6);

wire[27:0] addr_2177_6;

Selector_2 s2177_6(wires_544_5[1], addr_544_5, addr_positional[8711:8708], addr_2177_6);

wire[27:0] addr_2178_6;

Selector_2 s2178_6(wires_544_5[2], addr_544_5, addr_positional[8715:8712], addr_2178_6);

wire[27:0] addr_2179_6;

Selector_2 s2179_6(wires_544_5[3], addr_544_5, addr_positional[8719:8716], addr_2179_6);

wire[27:0] addr_2180_6;

Selector_2 s2180_6(wires_545_5[0], addr_545_5, addr_positional[8723:8720], addr_2180_6);

wire[27:0] addr_2181_6;

Selector_2 s2181_6(wires_545_5[1], addr_545_5, addr_positional[8727:8724], addr_2181_6);

wire[27:0] addr_2182_6;

Selector_2 s2182_6(wires_545_5[2], addr_545_5, addr_positional[8731:8728], addr_2182_6);

wire[27:0] addr_2183_6;

Selector_2 s2183_6(wires_545_5[3], addr_545_5, addr_positional[8735:8732], addr_2183_6);

wire[27:0] addr_2184_6;

Selector_2 s2184_6(wires_546_5[0], addr_546_5, addr_positional[8739:8736], addr_2184_6);

wire[27:0] addr_2185_6;

Selector_2 s2185_6(wires_546_5[1], addr_546_5, addr_positional[8743:8740], addr_2185_6);

wire[27:0] addr_2186_6;

Selector_2 s2186_6(wires_546_5[2], addr_546_5, addr_positional[8747:8744], addr_2186_6);

wire[27:0] addr_2187_6;

Selector_2 s2187_6(wires_546_5[3], addr_546_5, addr_positional[8751:8748], addr_2187_6);

wire[27:0] addr_2188_6;

Selector_2 s2188_6(wires_547_5[0], addr_547_5, addr_positional[8755:8752], addr_2188_6);

wire[27:0] addr_2189_6;

Selector_2 s2189_6(wires_547_5[1], addr_547_5, addr_positional[8759:8756], addr_2189_6);

wire[27:0] addr_2190_6;

Selector_2 s2190_6(wires_547_5[2], addr_547_5, addr_positional[8763:8760], addr_2190_6);

wire[27:0] addr_2191_6;

Selector_2 s2191_6(wires_547_5[3], addr_547_5, addr_positional[8767:8764], addr_2191_6);

wire[27:0] addr_2192_6;

Selector_2 s2192_6(wires_548_5[0], addr_548_5, addr_positional[8771:8768], addr_2192_6);

wire[27:0] addr_2193_6;

Selector_2 s2193_6(wires_548_5[1], addr_548_5, addr_positional[8775:8772], addr_2193_6);

wire[27:0] addr_2194_6;

Selector_2 s2194_6(wires_548_5[2], addr_548_5, addr_positional[8779:8776], addr_2194_6);

wire[27:0] addr_2195_6;

Selector_2 s2195_6(wires_548_5[3], addr_548_5, addr_positional[8783:8780], addr_2195_6);

wire[27:0] addr_2196_6;

Selector_2 s2196_6(wires_549_5[0], addr_549_5, addr_positional[8787:8784], addr_2196_6);

wire[27:0] addr_2197_6;

Selector_2 s2197_6(wires_549_5[1], addr_549_5, addr_positional[8791:8788], addr_2197_6);

wire[27:0] addr_2198_6;

Selector_2 s2198_6(wires_549_5[2], addr_549_5, addr_positional[8795:8792], addr_2198_6);

wire[27:0] addr_2199_6;

Selector_2 s2199_6(wires_549_5[3], addr_549_5, addr_positional[8799:8796], addr_2199_6);

wire[27:0] addr_2200_6;

Selector_2 s2200_6(wires_550_5[0], addr_550_5, addr_positional[8803:8800], addr_2200_6);

wire[27:0] addr_2201_6;

Selector_2 s2201_6(wires_550_5[1], addr_550_5, addr_positional[8807:8804], addr_2201_6);

wire[27:0] addr_2202_6;

Selector_2 s2202_6(wires_550_5[2], addr_550_5, addr_positional[8811:8808], addr_2202_6);

wire[27:0] addr_2203_6;

Selector_2 s2203_6(wires_550_5[3], addr_550_5, addr_positional[8815:8812], addr_2203_6);

wire[27:0] addr_2204_6;

Selector_2 s2204_6(wires_551_5[0], addr_551_5, addr_positional[8819:8816], addr_2204_6);

wire[27:0] addr_2205_6;

Selector_2 s2205_6(wires_551_5[1], addr_551_5, addr_positional[8823:8820], addr_2205_6);

wire[27:0] addr_2206_6;

Selector_2 s2206_6(wires_551_5[2], addr_551_5, addr_positional[8827:8824], addr_2206_6);

wire[27:0] addr_2207_6;

Selector_2 s2207_6(wires_551_5[3], addr_551_5, addr_positional[8831:8828], addr_2207_6);

wire[27:0] addr_2208_6;

Selector_2 s2208_6(wires_552_5[0], addr_552_5, addr_positional[8835:8832], addr_2208_6);

wire[27:0] addr_2209_6;

Selector_2 s2209_6(wires_552_5[1], addr_552_5, addr_positional[8839:8836], addr_2209_6);

wire[27:0] addr_2210_6;

Selector_2 s2210_6(wires_552_5[2], addr_552_5, addr_positional[8843:8840], addr_2210_6);

wire[27:0] addr_2211_6;

Selector_2 s2211_6(wires_552_5[3], addr_552_5, addr_positional[8847:8844], addr_2211_6);

wire[27:0] addr_2212_6;

Selector_2 s2212_6(wires_553_5[0], addr_553_5, addr_positional[8851:8848], addr_2212_6);

wire[27:0] addr_2213_6;

Selector_2 s2213_6(wires_553_5[1], addr_553_5, addr_positional[8855:8852], addr_2213_6);

wire[27:0] addr_2214_6;

Selector_2 s2214_6(wires_553_5[2], addr_553_5, addr_positional[8859:8856], addr_2214_6);

wire[27:0] addr_2215_6;

Selector_2 s2215_6(wires_553_5[3], addr_553_5, addr_positional[8863:8860], addr_2215_6);

wire[27:0] addr_2216_6;

Selector_2 s2216_6(wires_554_5[0], addr_554_5, addr_positional[8867:8864], addr_2216_6);

wire[27:0] addr_2217_6;

Selector_2 s2217_6(wires_554_5[1], addr_554_5, addr_positional[8871:8868], addr_2217_6);

wire[27:0] addr_2218_6;

Selector_2 s2218_6(wires_554_5[2], addr_554_5, addr_positional[8875:8872], addr_2218_6);

wire[27:0] addr_2219_6;

Selector_2 s2219_6(wires_554_5[3], addr_554_5, addr_positional[8879:8876], addr_2219_6);

wire[27:0] addr_2220_6;

Selector_2 s2220_6(wires_555_5[0], addr_555_5, addr_positional[8883:8880], addr_2220_6);

wire[27:0] addr_2221_6;

Selector_2 s2221_6(wires_555_5[1], addr_555_5, addr_positional[8887:8884], addr_2221_6);

wire[27:0] addr_2222_6;

Selector_2 s2222_6(wires_555_5[2], addr_555_5, addr_positional[8891:8888], addr_2222_6);

wire[27:0] addr_2223_6;

Selector_2 s2223_6(wires_555_5[3], addr_555_5, addr_positional[8895:8892], addr_2223_6);

wire[27:0] addr_2224_6;

Selector_2 s2224_6(wires_556_5[0], addr_556_5, addr_positional[8899:8896], addr_2224_6);

wire[27:0] addr_2225_6;

Selector_2 s2225_6(wires_556_5[1], addr_556_5, addr_positional[8903:8900], addr_2225_6);

wire[27:0] addr_2226_6;

Selector_2 s2226_6(wires_556_5[2], addr_556_5, addr_positional[8907:8904], addr_2226_6);

wire[27:0] addr_2227_6;

Selector_2 s2227_6(wires_556_5[3], addr_556_5, addr_positional[8911:8908], addr_2227_6);

wire[27:0] addr_2228_6;

Selector_2 s2228_6(wires_557_5[0], addr_557_5, addr_positional[8915:8912], addr_2228_6);

wire[27:0] addr_2229_6;

Selector_2 s2229_6(wires_557_5[1], addr_557_5, addr_positional[8919:8916], addr_2229_6);

wire[27:0] addr_2230_6;

Selector_2 s2230_6(wires_557_5[2], addr_557_5, addr_positional[8923:8920], addr_2230_6);

wire[27:0] addr_2231_6;

Selector_2 s2231_6(wires_557_5[3], addr_557_5, addr_positional[8927:8924], addr_2231_6);

wire[27:0] addr_2232_6;

Selector_2 s2232_6(wires_558_5[0], addr_558_5, addr_positional[8931:8928], addr_2232_6);

wire[27:0] addr_2233_6;

Selector_2 s2233_6(wires_558_5[1], addr_558_5, addr_positional[8935:8932], addr_2233_6);

wire[27:0] addr_2234_6;

Selector_2 s2234_6(wires_558_5[2], addr_558_5, addr_positional[8939:8936], addr_2234_6);

wire[27:0] addr_2235_6;

Selector_2 s2235_6(wires_558_5[3], addr_558_5, addr_positional[8943:8940], addr_2235_6);

wire[27:0] addr_2236_6;

Selector_2 s2236_6(wires_559_5[0], addr_559_5, addr_positional[8947:8944], addr_2236_6);

wire[27:0] addr_2237_6;

Selector_2 s2237_6(wires_559_5[1], addr_559_5, addr_positional[8951:8948], addr_2237_6);

wire[27:0] addr_2238_6;

Selector_2 s2238_6(wires_559_5[2], addr_559_5, addr_positional[8955:8952], addr_2238_6);

wire[27:0] addr_2239_6;

Selector_2 s2239_6(wires_559_5[3], addr_559_5, addr_positional[8959:8956], addr_2239_6);

wire[27:0] addr_2240_6;

Selector_2 s2240_6(wires_560_5[0], addr_560_5, addr_positional[8963:8960], addr_2240_6);

wire[27:0] addr_2241_6;

Selector_2 s2241_6(wires_560_5[1], addr_560_5, addr_positional[8967:8964], addr_2241_6);

wire[27:0] addr_2242_6;

Selector_2 s2242_6(wires_560_5[2], addr_560_5, addr_positional[8971:8968], addr_2242_6);

wire[27:0] addr_2243_6;

Selector_2 s2243_6(wires_560_5[3], addr_560_5, addr_positional[8975:8972], addr_2243_6);

wire[27:0] addr_2244_6;

Selector_2 s2244_6(wires_561_5[0], addr_561_5, addr_positional[8979:8976], addr_2244_6);

wire[27:0] addr_2245_6;

Selector_2 s2245_6(wires_561_5[1], addr_561_5, addr_positional[8983:8980], addr_2245_6);

wire[27:0] addr_2246_6;

Selector_2 s2246_6(wires_561_5[2], addr_561_5, addr_positional[8987:8984], addr_2246_6);

wire[27:0] addr_2247_6;

Selector_2 s2247_6(wires_561_5[3], addr_561_5, addr_positional[8991:8988], addr_2247_6);

wire[27:0] addr_2248_6;

Selector_2 s2248_6(wires_562_5[0], addr_562_5, addr_positional[8995:8992], addr_2248_6);

wire[27:0] addr_2249_6;

Selector_2 s2249_6(wires_562_5[1], addr_562_5, addr_positional[8999:8996], addr_2249_6);

wire[27:0] addr_2250_6;

Selector_2 s2250_6(wires_562_5[2], addr_562_5, addr_positional[9003:9000], addr_2250_6);

wire[27:0] addr_2251_6;

Selector_2 s2251_6(wires_562_5[3], addr_562_5, addr_positional[9007:9004], addr_2251_6);

wire[27:0] addr_2252_6;

Selector_2 s2252_6(wires_563_5[0], addr_563_5, addr_positional[9011:9008], addr_2252_6);

wire[27:0] addr_2253_6;

Selector_2 s2253_6(wires_563_5[1], addr_563_5, addr_positional[9015:9012], addr_2253_6);

wire[27:0] addr_2254_6;

Selector_2 s2254_6(wires_563_5[2], addr_563_5, addr_positional[9019:9016], addr_2254_6);

wire[27:0] addr_2255_6;

Selector_2 s2255_6(wires_563_5[3], addr_563_5, addr_positional[9023:9020], addr_2255_6);

wire[27:0] addr_2256_6;

Selector_2 s2256_6(wires_564_5[0], addr_564_5, addr_positional[9027:9024], addr_2256_6);

wire[27:0] addr_2257_6;

Selector_2 s2257_6(wires_564_5[1], addr_564_5, addr_positional[9031:9028], addr_2257_6);

wire[27:0] addr_2258_6;

Selector_2 s2258_6(wires_564_5[2], addr_564_5, addr_positional[9035:9032], addr_2258_6);

wire[27:0] addr_2259_6;

Selector_2 s2259_6(wires_564_5[3], addr_564_5, addr_positional[9039:9036], addr_2259_6);

wire[27:0] addr_2260_6;

Selector_2 s2260_6(wires_565_5[0], addr_565_5, addr_positional[9043:9040], addr_2260_6);

wire[27:0] addr_2261_6;

Selector_2 s2261_6(wires_565_5[1], addr_565_5, addr_positional[9047:9044], addr_2261_6);

wire[27:0] addr_2262_6;

Selector_2 s2262_6(wires_565_5[2], addr_565_5, addr_positional[9051:9048], addr_2262_6);

wire[27:0] addr_2263_6;

Selector_2 s2263_6(wires_565_5[3], addr_565_5, addr_positional[9055:9052], addr_2263_6);

wire[27:0] addr_2264_6;

Selector_2 s2264_6(wires_566_5[0], addr_566_5, addr_positional[9059:9056], addr_2264_6);

wire[27:0] addr_2265_6;

Selector_2 s2265_6(wires_566_5[1], addr_566_5, addr_positional[9063:9060], addr_2265_6);

wire[27:0] addr_2266_6;

Selector_2 s2266_6(wires_566_5[2], addr_566_5, addr_positional[9067:9064], addr_2266_6);

wire[27:0] addr_2267_6;

Selector_2 s2267_6(wires_566_5[3], addr_566_5, addr_positional[9071:9068], addr_2267_6);

wire[27:0] addr_2268_6;

Selector_2 s2268_6(wires_567_5[0], addr_567_5, addr_positional[9075:9072], addr_2268_6);

wire[27:0] addr_2269_6;

Selector_2 s2269_6(wires_567_5[1], addr_567_5, addr_positional[9079:9076], addr_2269_6);

wire[27:0] addr_2270_6;

Selector_2 s2270_6(wires_567_5[2], addr_567_5, addr_positional[9083:9080], addr_2270_6);

wire[27:0] addr_2271_6;

Selector_2 s2271_6(wires_567_5[3], addr_567_5, addr_positional[9087:9084], addr_2271_6);

wire[27:0] addr_2272_6;

Selector_2 s2272_6(wires_568_5[0], addr_568_5, addr_positional[9091:9088], addr_2272_6);

wire[27:0] addr_2273_6;

Selector_2 s2273_6(wires_568_5[1], addr_568_5, addr_positional[9095:9092], addr_2273_6);

wire[27:0] addr_2274_6;

Selector_2 s2274_6(wires_568_5[2], addr_568_5, addr_positional[9099:9096], addr_2274_6);

wire[27:0] addr_2275_6;

Selector_2 s2275_6(wires_568_5[3], addr_568_5, addr_positional[9103:9100], addr_2275_6);

wire[27:0] addr_2276_6;

Selector_2 s2276_6(wires_569_5[0], addr_569_5, addr_positional[9107:9104], addr_2276_6);

wire[27:0] addr_2277_6;

Selector_2 s2277_6(wires_569_5[1], addr_569_5, addr_positional[9111:9108], addr_2277_6);

wire[27:0] addr_2278_6;

Selector_2 s2278_6(wires_569_5[2], addr_569_5, addr_positional[9115:9112], addr_2278_6);

wire[27:0] addr_2279_6;

Selector_2 s2279_6(wires_569_5[3], addr_569_5, addr_positional[9119:9116], addr_2279_6);

wire[27:0] addr_2280_6;

Selector_2 s2280_6(wires_570_5[0], addr_570_5, addr_positional[9123:9120], addr_2280_6);

wire[27:0] addr_2281_6;

Selector_2 s2281_6(wires_570_5[1], addr_570_5, addr_positional[9127:9124], addr_2281_6);

wire[27:0] addr_2282_6;

Selector_2 s2282_6(wires_570_5[2], addr_570_5, addr_positional[9131:9128], addr_2282_6);

wire[27:0] addr_2283_6;

Selector_2 s2283_6(wires_570_5[3], addr_570_5, addr_positional[9135:9132], addr_2283_6);

wire[27:0] addr_2284_6;

Selector_2 s2284_6(wires_571_5[0], addr_571_5, addr_positional[9139:9136], addr_2284_6);

wire[27:0] addr_2285_6;

Selector_2 s2285_6(wires_571_5[1], addr_571_5, addr_positional[9143:9140], addr_2285_6);

wire[27:0] addr_2286_6;

Selector_2 s2286_6(wires_571_5[2], addr_571_5, addr_positional[9147:9144], addr_2286_6);

wire[27:0] addr_2287_6;

Selector_2 s2287_6(wires_571_5[3], addr_571_5, addr_positional[9151:9148], addr_2287_6);

wire[27:0] addr_2288_6;

Selector_2 s2288_6(wires_572_5[0], addr_572_5, addr_positional[9155:9152], addr_2288_6);

wire[27:0] addr_2289_6;

Selector_2 s2289_6(wires_572_5[1], addr_572_5, addr_positional[9159:9156], addr_2289_6);

wire[27:0] addr_2290_6;

Selector_2 s2290_6(wires_572_5[2], addr_572_5, addr_positional[9163:9160], addr_2290_6);

wire[27:0] addr_2291_6;

Selector_2 s2291_6(wires_572_5[3], addr_572_5, addr_positional[9167:9164], addr_2291_6);

wire[27:0] addr_2292_6;

Selector_2 s2292_6(wires_573_5[0], addr_573_5, addr_positional[9171:9168], addr_2292_6);

wire[27:0] addr_2293_6;

Selector_2 s2293_6(wires_573_5[1], addr_573_5, addr_positional[9175:9172], addr_2293_6);

wire[27:0] addr_2294_6;

Selector_2 s2294_6(wires_573_5[2], addr_573_5, addr_positional[9179:9176], addr_2294_6);

wire[27:0] addr_2295_6;

Selector_2 s2295_6(wires_573_5[3], addr_573_5, addr_positional[9183:9180], addr_2295_6);

wire[27:0] addr_2296_6;

Selector_2 s2296_6(wires_574_5[0], addr_574_5, addr_positional[9187:9184], addr_2296_6);

wire[27:0] addr_2297_6;

Selector_2 s2297_6(wires_574_5[1], addr_574_5, addr_positional[9191:9188], addr_2297_6);

wire[27:0] addr_2298_6;

Selector_2 s2298_6(wires_574_5[2], addr_574_5, addr_positional[9195:9192], addr_2298_6);

wire[27:0] addr_2299_6;

Selector_2 s2299_6(wires_574_5[3], addr_574_5, addr_positional[9199:9196], addr_2299_6);

wire[27:0] addr_2300_6;

Selector_2 s2300_6(wires_575_5[0], addr_575_5, addr_positional[9203:9200], addr_2300_6);

wire[27:0] addr_2301_6;

Selector_2 s2301_6(wires_575_5[1], addr_575_5, addr_positional[9207:9204], addr_2301_6);

wire[27:0] addr_2302_6;

Selector_2 s2302_6(wires_575_5[2], addr_575_5, addr_positional[9211:9208], addr_2302_6);

wire[27:0] addr_2303_6;

Selector_2 s2303_6(wires_575_5[3], addr_575_5, addr_positional[9215:9212], addr_2303_6);

wire[27:0] addr_2304_6;

Selector_2 s2304_6(wires_576_5[0], addr_576_5, addr_positional[9219:9216], addr_2304_6);

wire[27:0] addr_2305_6;

Selector_2 s2305_6(wires_576_5[1], addr_576_5, addr_positional[9223:9220], addr_2305_6);

wire[27:0] addr_2306_6;

Selector_2 s2306_6(wires_576_5[2], addr_576_5, addr_positional[9227:9224], addr_2306_6);

wire[27:0] addr_2307_6;

Selector_2 s2307_6(wires_576_5[3], addr_576_5, addr_positional[9231:9228], addr_2307_6);

wire[27:0] addr_2308_6;

Selector_2 s2308_6(wires_577_5[0], addr_577_5, addr_positional[9235:9232], addr_2308_6);

wire[27:0] addr_2309_6;

Selector_2 s2309_6(wires_577_5[1], addr_577_5, addr_positional[9239:9236], addr_2309_6);

wire[27:0] addr_2310_6;

Selector_2 s2310_6(wires_577_5[2], addr_577_5, addr_positional[9243:9240], addr_2310_6);

wire[27:0] addr_2311_6;

Selector_2 s2311_6(wires_577_5[3], addr_577_5, addr_positional[9247:9244], addr_2311_6);

wire[27:0] addr_2312_6;

Selector_2 s2312_6(wires_578_5[0], addr_578_5, addr_positional[9251:9248], addr_2312_6);

wire[27:0] addr_2313_6;

Selector_2 s2313_6(wires_578_5[1], addr_578_5, addr_positional[9255:9252], addr_2313_6);

wire[27:0] addr_2314_6;

Selector_2 s2314_6(wires_578_5[2], addr_578_5, addr_positional[9259:9256], addr_2314_6);

wire[27:0] addr_2315_6;

Selector_2 s2315_6(wires_578_5[3], addr_578_5, addr_positional[9263:9260], addr_2315_6);

wire[27:0] addr_2316_6;

Selector_2 s2316_6(wires_579_5[0], addr_579_5, addr_positional[9267:9264], addr_2316_6);

wire[27:0] addr_2317_6;

Selector_2 s2317_6(wires_579_5[1], addr_579_5, addr_positional[9271:9268], addr_2317_6);

wire[27:0] addr_2318_6;

Selector_2 s2318_6(wires_579_5[2], addr_579_5, addr_positional[9275:9272], addr_2318_6);

wire[27:0] addr_2319_6;

Selector_2 s2319_6(wires_579_5[3], addr_579_5, addr_positional[9279:9276], addr_2319_6);

wire[27:0] addr_2320_6;

Selector_2 s2320_6(wires_580_5[0], addr_580_5, addr_positional[9283:9280], addr_2320_6);

wire[27:0] addr_2321_6;

Selector_2 s2321_6(wires_580_5[1], addr_580_5, addr_positional[9287:9284], addr_2321_6);

wire[27:0] addr_2322_6;

Selector_2 s2322_6(wires_580_5[2], addr_580_5, addr_positional[9291:9288], addr_2322_6);

wire[27:0] addr_2323_6;

Selector_2 s2323_6(wires_580_5[3], addr_580_5, addr_positional[9295:9292], addr_2323_6);

wire[27:0] addr_2324_6;

Selector_2 s2324_6(wires_581_5[0], addr_581_5, addr_positional[9299:9296], addr_2324_6);

wire[27:0] addr_2325_6;

Selector_2 s2325_6(wires_581_5[1], addr_581_5, addr_positional[9303:9300], addr_2325_6);

wire[27:0] addr_2326_6;

Selector_2 s2326_6(wires_581_5[2], addr_581_5, addr_positional[9307:9304], addr_2326_6);

wire[27:0] addr_2327_6;

Selector_2 s2327_6(wires_581_5[3], addr_581_5, addr_positional[9311:9308], addr_2327_6);

wire[27:0] addr_2328_6;

Selector_2 s2328_6(wires_582_5[0], addr_582_5, addr_positional[9315:9312], addr_2328_6);

wire[27:0] addr_2329_6;

Selector_2 s2329_6(wires_582_5[1], addr_582_5, addr_positional[9319:9316], addr_2329_6);

wire[27:0] addr_2330_6;

Selector_2 s2330_6(wires_582_5[2], addr_582_5, addr_positional[9323:9320], addr_2330_6);

wire[27:0] addr_2331_6;

Selector_2 s2331_6(wires_582_5[3], addr_582_5, addr_positional[9327:9324], addr_2331_6);

wire[27:0] addr_2332_6;

Selector_2 s2332_6(wires_583_5[0], addr_583_5, addr_positional[9331:9328], addr_2332_6);

wire[27:0] addr_2333_6;

Selector_2 s2333_6(wires_583_5[1], addr_583_5, addr_positional[9335:9332], addr_2333_6);

wire[27:0] addr_2334_6;

Selector_2 s2334_6(wires_583_5[2], addr_583_5, addr_positional[9339:9336], addr_2334_6);

wire[27:0] addr_2335_6;

Selector_2 s2335_6(wires_583_5[3], addr_583_5, addr_positional[9343:9340], addr_2335_6);

wire[27:0] addr_2336_6;

Selector_2 s2336_6(wires_584_5[0], addr_584_5, addr_positional[9347:9344], addr_2336_6);

wire[27:0] addr_2337_6;

Selector_2 s2337_6(wires_584_5[1], addr_584_5, addr_positional[9351:9348], addr_2337_6);

wire[27:0] addr_2338_6;

Selector_2 s2338_6(wires_584_5[2], addr_584_5, addr_positional[9355:9352], addr_2338_6);

wire[27:0] addr_2339_6;

Selector_2 s2339_6(wires_584_5[3], addr_584_5, addr_positional[9359:9356], addr_2339_6);

wire[27:0] addr_2340_6;

Selector_2 s2340_6(wires_585_5[0], addr_585_5, addr_positional[9363:9360], addr_2340_6);

wire[27:0] addr_2341_6;

Selector_2 s2341_6(wires_585_5[1], addr_585_5, addr_positional[9367:9364], addr_2341_6);

wire[27:0] addr_2342_6;

Selector_2 s2342_6(wires_585_5[2], addr_585_5, addr_positional[9371:9368], addr_2342_6);

wire[27:0] addr_2343_6;

Selector_2 s2343_6(wires_585_5[3], addr_585_5, addr_positional[9375:9372], addr_2343_6);

wire[27:0] addr_2344_6;

Selector_2 s2344_6(wires_586_5[0], addr_586_5, addr_positional[9379:9376], addr_2344_6);

wire[27:0] addr_2345_6;

Selector_2 s2345_6(wires_586_5[1], addr_586_5, addr_positional[9383:9380], addr_2345_6);

wire[27:0] addr_2346_6;

Selector_2 s2346_6(wires_586_5[2], addr_586_5, addr_positional[9387:9384], addr_2346_6);

wire[27:0] addr_2347_6;

Selector_2 s2347_6(wires_586_5[3], addr_586_5, addr_positional[9391:9388], addr_2347_6);

wire[27:0] addr_2348_6;

Selector_2 s2348_6(wires_587_5[0], addr_587_5, addr_positional[9395:9392], addr_2348_6);

wire[27:0] addr_2349_6;

Selector_2 s2349_6(wires_587_5[1], addr_587_5, addr_positional[9399:9396], addr_2349_6);

wire[27:0] addr_2350_6;

Selector_2 s2350_6(wires_587_5[2], addr_587_5, addr_positional[9403:9400], addr_2350_6);

wire[27:0] addr_2351_6;

Selector_2 s2351_6(wires_587_5[3], addr_587_5, addr_positional[9407:9404], addr_2351_6);

wire[27:0] addr_2352_6;

Selector_2 s2352_6(wires_588_5[0], addr_588_5, addr_positional[9411:9408], addr_2352_6);

wire[27:0] addr_2353_6;

Selector_2 s2353_6(wires_588_5[1], addr_588_5, addr_positional[9415:9412], addr_2353_6);

wire[27:0] addr_2354_6;

Selector_2 s2354_6(wires_588_5[2], addr_588_5, addr_positional[9419:9416], addr_2354_6);

wire[27:0] addr_2355_6;

Selector_2 s2355_6(wires_588_5[3], addr_588_5, addr_positional[9423:9420], addr_2355_6);

wire[27:0] addr_2356_6;

Selector_2 s2356_6(wires_589_5[0], addr_589_5, addr_positional[9427:9424], addr_2356_6);

wire[27:0] addr_2357_6;

Selector_2 s2357_6(wires_589_5[1], addr_589_5, addr_positional[9431:9428], addr_2357_6);

wire[27:0] addr_2358_6;

Selector_2 s2358_6(wires_589_5[2], addr_589_5, addr_positional[9435:9432], addr_2358_6);

wire[27:0] addr_2359_6;

Selector_2 s2359_6(wires_589_5[3], addr_589_5, addr_positional[9439:9436], addr_2359_6);

wire[27:0] addr_2360_6;

Selector_2 s2360_6(wires_590_5[0], addr_590_5, addr_positional[9443:9440], addr_2360_6);

wire[27:0] addr_2361_6;

Selector_2 s2361_6(wires_590_5[1], addr_590_5, addr_positional[9447:9444], addr_2361_6);

wire[27:0] addr_2362_6;

Selector_2 s2362_6(wires_590_5[2], addr_590_5, addr_positional[9451:9448], addr_2362_6);

wire[27:0] addr_2363_6;

Selector_2 s2363_6(wires_590_5[3], addr_590_5, addr_positional[9455:9452], addr_2363_6);

wire[27:0] addr_2364_6;

Selector_2 s2364_6(wires_591_5[0], addr_591_5, addr_positional[9459:9456], addr_2364_6);

wire[27:0] addr_2365_6;

Selector_2 s2365_6(wires_591_5[1], addr_591_5, addr_positional[9463:9460], addr_2365_6);

wire[27:0] addr_2366_6;

Selector_2 s2366_6(wires_591_5[2], addr_591_5, addr_positional[9467:9464], addr_2366_6);

wire[27:0] addr_2367_6;

Selector_2 s2367_6(wires_591_5[3], addr_591_5, addr_positional[9471:9468], addr_2367_6);

wire[27:0] addr_2368_6;

Selector_2 s2368_6(wires_592_5[0], addr_592_5, addr_positional[9475:9472], addr_2368_6);

wire[27:0] addr_2369_6;

Selector_2 s2369_6(wires_592_5[1], addr_592_5, addr_positional[9479:9476], addr_2369_6);

wire[27:0] addr_2370_6;

Selector_2 s2370_6(wires_592_5[2], addr_592_5, addr_positional[9483:9480], addr_2370_6);

wire[27:0] addr_2371_6;

Selector_2 s2371_6(wires_592_5[3], addr_592_5, addr_positional[9487:9484], addr_2371_6);

wire[27:0] addr_2372_6;

Selector_2 s2372_6(wires_593_5[0], addr_593_5, addr_positional[9491:9488], addr_2372_6);

wire[27:0] addr_2373_6;

Selector_2 s2373_6(wires_593_5[1], addr_593_5, addr_positional[9495:9492], addr_2373_6);

wire[27:0] addr_2374_6;

Selector_2 s2374_6(wires_593_5[2], addr_593_5, addr_positional[9499:9496], addr_2374_6);

wire[27:0] addr_2375_6;

Selector_2 s2375_6(wires_593_5[3], addr_593_5, addr_positional[9503:9500], addr_2375_6);

wire[27:0] addr_2376_6;

Selector_2 s2376_6(wires_594_5[0], addr_594_5, addr_positional[9507:9504], addr_2376_6);

wire[27:0] addr_2377_6;

Selector_2 s2377_6(wires_594_5[1], addr_594_5, addr_positional[9511:9508], addr_2377_6);

wire[27:0] addr_2378_6;

Selector_2 s2378_6(wires_594_5[2], addr_594_5, addr_positional[9515:9512], addr_2378_6);

wire[27:0] addr_2379_6;

Selector_2 s2379_6(wires_594_5[3], addr_594_5, addr_positional[9519:9516], addr_2379_6);

wire[27:0] addr_2380_6;

Selector_2 s2380_6(wires_595_5[0], addr_595_5, addr_positional[9523:9520], addr_2380_6);

wire[27:0] addr_2381_6;

Selector_2 s2381_6(wires_595_5[1], addr_595_5, addr_positional[9527:9524], addr_2381_6);

wire[27:0] addr_2382_6;

Selector_2 s2382_6(wires_595_5[2], addr_595_5, addr_positional[9531:9528], addr_2382_6);

wire[27:0] addr_2383_6;

Selector_2 s2383_6(wires_595_5[3], addr_595_5, addr_positional[9535:9532], addr_2383_6);

wire[27:0] addr_2384_6;

Selector_2 s2384_6(wires_596_5[0], addr_596_5, addr_positional[9539:9536], addr_2384_6);

wire[27:0] addr_2385_6;

Selector_2 s2385_6(wires_596_5[1], addr_596_5, addr_positional[9543:9540], addr_2385_6);

wire[27:0] addr_2386_6;

Selector_2 s2386_6(wires_596_5[2], addr_596_5, addr_positional[9547:9544], addr_2386_6);

wire[27:0] addr_2387_6;

Selector_2 s2387_6(wires_596_5[3], addr_596_5, addr_positional[9551:9548], addr_2387_6);

wire[27:0] addr_2388_6;

Selector_2 s2388_6(wires_597_5[0], addr_597_5, addr_positional[9555:9552], addr_2388_6);

wire[27:0] addr_2389_6;

Selector_2 s2389_6(wires_597_5[1], addr_597_5, addr_positional[9559:9556], addr_2389_6);

wire[27:0] addr_2390_6;

Selector_2 s2390_6(wires_597_5[2], addr_597_5, addr_positional[9563:9560], addr_2390_6);

wire[27:0] addr_2391_6;

Selector_2 s2391_6(wires_597_5[3], addr_597_5, addr_positional[9567:9564], addr_2391_6);

wire[27:0] addr_2392_6;

Selector_2 s2392_6(wires_598_5[0], addr_598_5, addr_positional[9571:9568], addr_2392_6);

wire[27:0] addr_2393_6;

Selector_2 s2393_6(wires_598_5[1], addr_598_5, addr_positional[9575:9572], addr_2393_6);

wire[27:0] addr_2394_6;

Selector_2 s2394_6(wires_598_5[2], addr_598_5, addr_positional[9579:9576], addr_2394_6);

wire[27:0] addr_2395_6;

Selector_2 s2395_6(wires_598_5[3], addr_598_5, addr_positional[9583:9580], addr_2395_6);

wire[27:0] addr_2396_6;

Selector_2 s2396_6(wires_599_5[0], addr_599_5, addr_positional[9587:9584], addr_2396_6);

wire[27:0] addr_2397_6;

Selector_2 s2397_6(wires_599_5[1], addr_599_5, addr_positional[9591:9588], addr_2397_6);

wire[27:0] addr_2398_6;

Selector_2 s2398_6(wires_599_5[2], addr_599_5, addr_positional[9595:9592], addr_2398_6);

wire[27:0] addr_2399_6;

Selector_2 s2399_6(wires_599_5[3], addr_599_5, addr_positional[9599:9596], addr_2399_6);

wire[27:0] addr_2400_6;

Selector_2 s2400_6(wires_600_5[0], addr_600_5, addr_positional[9603:9600], addr_2400_6);

wire[27:0] addr_2401_6;

Selector_2 s2401_6(wires_600_5[1], addr_600_5, addr_positional[9607:9604], addr_2401_6);

wire[27:0] addr_2402_6;

Selector_2 s2402_6(wires_600_5[2], addr_600_5, addr_positional[9611:9608], addr_2402_6);

wire[27:0] addr_2403_6;

Selector_2 s2403_6(wires_600_5[3], addr_600_5, addr_positional[9615:9612], addr_2403_6);

wire[27:0] addr_2404_6;

Selector_2 s2404_6(wires_601_5[0], addr_601_5, addr_positional[9619:9616], addr_2404_6);

wire[27:0] addr_2405_6;

Selector_2 s2405_6(wires_601_5[1], addr_601_5, addr_positional[9623:9620], addr_2405_6);

wire[27:0] addr_2406_6;

Selector_2 s2406_6(wires_601_5[2], addr_601_5, addr_positional[9627:9624], addr_2406_6);

wire[27:0] addr_2407_6;

Selector_2 s2407_6(wires_601_5[3], addr_601_5, addr_positional[9631:9628], addr_2407_6);

wire[27:0] addr_2408_6;

Selector_2 s2408_6(wires_602_5[0], addr_602_5, addr_positional[9635:9632], addr_2408_6);

wire[27:0] addr_2409_6;

Selector_2 s2409_6(wires_602_5[1], addr_602_5, addr_positional[9639:9636], addr_2409_6);

wire[27:0] addr_2410_6;

Selector_2 s2410_6(wires_602_5[2], addr_602_5, addr_positional[9643:9640], addr_2410_6);

wire[27:0] addr_2411_6;

Selector_2 s2411_6(wires_602_5[3], addr_602_5, addr_positional[9647:9644], addr_2411_6);

wire[27:0] addr_2412_6;

Selector_2 s2412_6(wires_603_5[0], addr_603_5, addr_positional[9651:9648], addr_2412_6);

wire[27:0] addr_2413_6;

Selector_2 s2413_6(wires_603_5[1], addr_603_5, addr_positional[9655:9652], addr_2413_6);

wire[27:0] addr_2414_6;

Selector_2 s2414_6(wires_603_5[2], addr_603_5, addr_positional[9659:9656], addr_2414_6);

wire[27:0] addr_2415_6;

Selector_2 s2415_6(wires_603_5[3], addr_603_5, addr_positional[9663:9660], addr_2415_6);

wire[27:0] addr_2416_6;

Selector_2 s2416_6(wires_604_5[0], addr_604_5, addr_positional[9667:9664], addr_2416_6);

wire[27:0] addr_2417_6;

Selector_2 s2417_6(wires_604_5[1], addr_604_5, addr_positional[9671:9668], addr_2417_6);

wire[27:0] addr_2418_6;

Selector_2 s2418_6(wires_604_5[2], addr_604_5, addr_positional[9675:9672], addr_2418_6);

wire[27:0] addr_2419_6;

Selector_2 s2419_6(wires_604_5[3], addr_604_5, addr_positional[9679:9676], addr_2419_6);

wire[27:0] addr_2420_6;

Selector_2 s2420_6(wires_605_5[0], addr_605_5, addr_positional[9683:9680], addr_2420_6);

wire[27:0] addr_2421_6;

Selector_2 s2421_6(wires_605_5[1], addr_605_5, addr_positional[9687:9684], addr_2421_6);

wire[27:0] addr_2422_6;

Selector_2 s2422_6(wires_605_5[2], addr_605_5, addr_positional[9691:9688], addr_2422_6);

wire[27:0] addr_2423_6;

Selector_2 s2423_6(wires_605_5[3], addr_605_5, addr_positional[9695:9692], addr_2423_6);

wire[27:0] addr_2424_6;

Selector_2 s2424_6(wires_606_5[0], addr_606_5, addr_positional[9699:9696], addr_2424_6);

wire[27:0] addr_2425_6;

Selector_2 s2425_6(wires_606_5[1], addr_606_5, addr_positional[9703:9700], addr_2425_6);

wire[27:0] addr_2426_6;

Selector_2 s2426_6(wires_606_5[2], addr_606_5, addr_positional[9707:9704], addr_2426_6);

wire[27:0] addr_2427_6;

Selector_2 s2427_6(wires_606_5[3], addr_606_5, addr_positional[9711:9708], addr_2427_6);

wire[27:0] addr_2428_6;

Selector_2 s2428_6(wires_607_5[0], addr_607_5, addr_positional[9715:9712], addr_2428_6);

wire[27:0] addr_2429_6;

Selector_2 s2429_6(wires_607_5[1], addr_607_5, addr_positional[9719:9716], addr_2429_6);

wire[27:0] addr_2430_6;

Selector_2 s2430_6(wires_607_5[2], addr_607_5, addr_positional[9723:9720], addr_2430_6);

wire[27:0] addr_2431_6;

Selector_2 s2431_6(wires_607_5[3], addr_607_5, addr_positional[9727:9724], addr_2431_6);

wire[27:0] addr_2432_6;

Selector_2 s2432_6(wires_608_5[0], addr_608_5, addr_positional[9731:9728], addr_2432_6);

wire[27:0] addr_2433_6;

Selector_2 s2433_6(wires_608_5[1], addr_608_5, addr_positional[9735:9732], addr_2433_6);

wire[27:0] addr_2434_6;

Selector_2 s2434_6(wires_608_5[2], addr_608_5, addr_positional[9739:9736], addr_2434_6);

wire[27:0] addr_2435_6;

Selector_2 s2435_6(wires_608_5[3], addr_608_5, addr_positional[9743:9740], addr_2435_6);

wire[27:0] addr_2436_6;

Selector_2 s2436_6(wires_609_5[0], addr_609_5, addr_positional[9747:9744], addr_2436_6);

wire[27:0] addr_2437_6;

Selector_2 s2437_6(wires_609_5[1], addr_609_5, addr_positional[9751:9748], addr_2437_6);

wire[27:0] addr_2438_6;

Selector_2 s2438_6(wires_609_5[2], addr_609_5, addr_positional[9755:9752], addr_2438_6);

wire[27:0] addr_2439_6;

Selector_2 s2439_6(wires_609_5[3], addr_609_5, addr_positional[9759:9756], addr_2439_6);

wire[27:0] addr_2440_6;

Selector_2 s2440_6(wires_610_5[0], addr_610_5, addr_positional[9763:9760], addr_2440_6);

wire[27:0] addr_2441_6;

Selector_2 s2441_6(wires_610_5[1], addr_610_5, addr_positional[9767:9764], addr_2441_6);

wire[27:0] addr_2442_6;

Selector_2 s2442_6(wires_610_5[2], addr_610_5, addr_positional[9771:9768], addr_2442_6);

wire[27:0] addr_2443_6;

Selector_2 s2443_6(wires_610_5[3], addr_610_5, addr_positional[9775:9772], addr_2443_6);

wire[27:0] addr_2444_6;

Selector_2 s2444_6(wires_611_5[0], addr_611_5, addr_positional[9779:9776], addr_2444_6);

wire[27:0] addr_2445_6;

Selector_2 s2445_6(wires_611_5[1], addr_611_5, addr_positional[9783:9780], addr_2445_6);

wire[27:0] addr_2446_6;

Selector_2 s2446_6(wires_611_5[2], addr_611_5, addr_positional[9787:9784], addr_2446_6);

wire[27:0] addr_2447_6;

Selector_2 s2447_6(wires_611_5[3], addr_611_5, addr_positional[9791:9788], addr_2447_6);

wire[27:0] addr_2448_6;

Selector_2 s2448_6(wires_612_5[0], addr_612_5, addr_positional[9795:9792], addr_2448_6);

wire[27:0] addr_2449_6;

Selector_2 s2449_6(wires_612_5[1], addr_612_5, addr_positional[9799:9796], addr_2449_6);

wire[27:0] addr_2450_6;

Selector_2 s2450_6(wires_612_5[2], addr_612_5, addr_positional[9803:9800], addr_2450_6);

wire[27:0] addr_2451_6;

Selector_2 s2451_6(wires_612_5[3], addr_612_5, addr_positional[9807:9804], addr_2451_6);

wire[27:0] addr_2452_6;

Selector_2 s2452_6(wires_613_5[0], addr_613_5, addr_positional[9811:9808], addr_2452_6);

wire[27:0] addr_2453_6;

Selector_2 s2453_6(wires_613_5[1], addr_613_5, addr_positional[9815:9812], addr_2453_6);

wire[27:0] addr_2454_6;

Selector_2 s2454_6(wires_613_5[2], addr_613_5, addr_positional[9819:9816], addr_2454_6);

wire[27:0] addr_2455_6;

Selector_2 s2455_6(wires_613_5[3], addr_613_5, addr_positional[9823:9820], addr_2455_6);

wire[27:0] addr_2456_6;

Selector_2 s2456_6(wires_614_5[0], addr_614_5, addr_positional[9827:9824], addr_2456_6);

wire[27:0] addr_2457_6;

Selector_2 s2457_6(wires_614_5[1], addr_614_5, addr_positional[9831:9828], addr_2457_6);

wire[27:0] addr_2458_6;

Selector_2 s2458_6(wires_614_5[2], addr_614_5, addr_positional[9835:9832], addr_2458_6);

wire[27:0] addr_2459_6;

Selector_2 s2459_6(wires_614_5[3], addr_614_5, addr_positional[9839:9836], addr_2459_6);

wire[27:0] addr_2460_6;

Selector_2 s2460_6(wires_615_5[0], addr_615_5, addr_positional[9843:9840], addr_2460_6);

wire[27:0] addr_2461_6;

Selector_2 s2461_6(wires_615_5[1], addr_615_5, addr_positional[9847:9844], addr_2461_6);

wire[27:0] addr_2462_6;

Selector_2 s2462_6(wires_615_5[2], addr_615_5, addr_positional[9851:9848], addr_2462_6);

wire[27:0] addr_2463_6;

Selector_2 s2463_6(wires_615_5[3], addr_615_5, addr_positional[9855:9852], addr_2463_6);

wire[27:0] addr_2464_6;

Selector_2 s2464_6(wires_616_5[0], addr_616_5, addr_positional[9859:9856], addr_2464_6);

wire[27:0] addr_2465_6;

Selector_2 s2465_6(wires_616_5[1], addr_616_5, addr_positional[9863:9860], addr_2465_6);

wire[27:0] addr_2466_6;

Selector_2 s2466_6(wires_616_5[2], addr_616_5, addr_positional[9867:9864], addr_2466_6);

wire[27:0] addr_2467_6;

Selector_2 s2467_6(wires_616_5[3], addr_616_5, addr_positional[9871:9868], addr_2467_6);

wire[27:0] addr_2468_6;

Selector_2 s2468_6(wires_617_5[0], addr_617_5, addr_positional[9875:9872], addr_2468_6);

wire[27:0] addr_2469_6;

Selector_2 s2469_6(wires_617_5[1], addr_617_5, addr_positional[9879:9876], addr_2469_6);

wire[27:0] addr_2470_6;

Selector_2 s2470_6(wires_617_5[2], addr_617_5, addr_positional[9883:9880], addr_2470_6);

wire[27:0] addr_2471_6;

Selector_2 s2471_6(wires_617_5[3], addr_617_5, addr_positional[9887:9884], addr_2471_6);

wire[27:0] addr_2472_6;

Selector_2 s2472_6(wires_618_5[0], addr_618_5, addr_positional[9891:9888], addr_2472_6);

wire[27:0] addr_2473_6;

Selector_2 s2473_6(wires_618_5[1], addr_618_5, addr_positional[9895:9892], addr_2473_6);

wire[27:0] addr_2474_6;

Selector_2 s2474_6(wires_618_5[2], addr_618_5, addr_positional[9899:9896], addr_2474_6);

wire[27:0] addr_2475_6;

Selector_2 s2475_6(wires_618_5[3], addr_618_5, addr_positional[9903:9900], addr_2475_6);

wire[27:0] addr_2476_6;

Selector_2 s2476_6(wires_619_5[0], addr_619_5, addr_positional[9907:9904], addr_2476_6);

wire[27:0] addr_2477_6;

Selector_2 s2477_6(wires_619_5[1], addr_619_5, addr_positional[9911:9908], addr_2477_6);

wire[27:0] addr_2478_6;

Selector_2 s2478_6(wires_619_5[2], addr_619_5, addr_positional[9915:9912], addr_2478_6);

wire[27:0] addr_2479_6;

Selector_2 s2479_6(wires_619_5[3], addr_619_5, addr_positional[9919:9916], addr_2479_6);

wire[27:0] addr_2480_6;

Selector_2 s2480_6(wires_620_5[0], addr_620_5, addr_positional[9923:9920], addr_2480_6);

wire[27:0] addr_2481_6;

Selector_2 s2481_6(wires_620_5[1], addr_620_5, addr_positional[9927:9924], addr_2481_6);

wire[27:0] addr_2482_6;

Selector_2 s2482_6(wires_620_5[2], addr_620_5, addr_positional[9931:9928], addr_2482_6);

wire[27:0] addr_2483_6;

Selector_2 s2483_6(wires_620_5[3], addr_620_5, addr_positional[9935:9932], addr_2483_6);

wire[27:0] addr_2484_6;

Selector_2 s2484_6(wires_621_5[0], addr_621_5, addr_positional[9939:9936], addr_2484_6);

wire[27:0] addr_2485_6;

Selector_2 s2485_6(wires_621_5[1], addr_621_5, addr_positional[9943:9940], addr_2485_6);

wire[27:0] addr_2486_6;

Selector_2 s2486_6(wires_621_5[2], addr_621_5, addr_positional[9947:9944], addr_2486_6);

wire[27:0] addr_2487_6;

Selector_2 s2487_6(wires_621_5[3], addr_621_5, addr_positional[9951:9948], addr_2487_6);

wire[27:0] addr_2488_6;

Selector_2 s2488_6(wires_622_5[0], addr_622_5, addr_positional[9955:9952], addr_2488_6);

wire[27:0] addr_2489_6;

Selector_2 s2489_6(wires_622_5[1], addr_622_5, addr_positional[9959:9956], addr_2489_6);

wire[27:0] addr_2490_6;

Selector_2 s2490_6(wires_622_5[2], addr_622_5, addr_positional[9963:9960], addr_2490_6);

wire[27:0] addr_2491_6;

Selector_2 s2491_6(wires_622_5[3], addr_622_5, addr_positional[9967:9964], addr_2491_6);

wire[27:0] addr_2492_6;

Selector_2 s2492_6(wires_623_5[0], addr_623_5, addr_positional[9971:9968], addr_2492_6);

wire[27:0] addr_2493_6;

Selector_2 s2493_6(wires_623_5[1], addr_623_5, addr_positional[9975:9972], addr_2493_6);

wire[27:0] addr_2494_6;

Selector_2 s2494_6(wires_623_5[2], addr_623_5, addr_positional[9979:9976], addr_2494_6);

wire[27:0] addr_2495_6;

Selector_2 s2495_6(wires_623_5[3], addr_623_5, addr_positional[9983:9980], addr_2495_6);

wire[27:0] addr_2496_6;

Selector_2 s2496_6(wires_624_5[0], addr_624_5, addr_positional[9987:9984], addr_2496_6);

wire[27:0] addr_2497_6;

Selector_2 s2497_6(wires_624_5[1], addr_624_5, addr_positional[9991:9988], addr_2497_6);

wire[27:0] addr_2498_6;

Selector_2 s2498_6(wires_624_5[2], addr_624_5, addr_positional[9995:9992], addr_2498_6);

wire[27:0] addr_2499_6;

Selector_2 s2499_6(wires_624_5[3], addr_624_5, addr_positional[9999:9996], addr_2499_6);

wire[27:0] addr_2500_6;

Selector_2 s2500_6(wires_625_5[0], addr_625_5, addr_positional[10003:10000], addr_2500_6);

wire[27:0] addr_2501_6;

Selector_2 s2501_6(wires_625_5[1], addr_625_5, addr_positional[10007:10004], addr_2501_6);

wire[27:0] addr_2502_6;

Selector_2 s2502_6(wires_625_5[2], addr_625_5, addr_positional[10011:10008], addr_2502_6);

wire[27:0] addr_2503_6;

Selector_2 s2503_6(wires_625_5[3], addr_625_5, addr_positional[10015:10012], addr_2503_6);

wire[27:0] addr_2504_6;

Selector_2 s2504_6(wires_626_5[0], addr_626_5, addr_positional[10019:10016], addr_2504_6);

wire[27:0] addr_2505_6;

Selector_2 s2505_6(wires_626_5[1], addr_626_5, addr_positional[10023:10020], addr_2505_6);

wire[27:0] addr_2506_6;

Selector_2 s2506_6(wires_626_5[2], addr_626_5, addr_positional[10027:10024], addr_2506_6);

wire[27:0] addr_2507_6;

Selector_2 s2507_6(wires_626_5[3], addr_626_5, addr_positional[10031:10028], addr_2507_6);

wire[27:0] addr_2508_6;

Selector_2 s2508_6(wires_627_5[0], addr_627_5, addr_positional[10035:10032], addr_2508_6);

wire[27:0] addr_2509_6;

Selector_2 s2509_6(wires_627_5[1], addr_627_5, addr_positional[10039:10036], addr_2509_6);

wire[27:0] addr_2510_6;

Selector_2 s2510_6(wires_627_5[2], addr_627_5, addr_positional[10043:10040], addr_2510_6);

wire[27:0] addr_2511_6;

Selector_2 s2511_6(wires_627_5[3], addr_627_5, addr_positional[10047:10044], addr_2511_6);

wire[27:0] addr_2512_6;

Selector_2 s2512_6(wires_628_5[0], addr_628_5, addr_positional[10051:10048], addr_2512_6);

wire[27:0] addr_2513_6;

Selector_2 s2513_6(wires_628_5[1], addr_628_5, addr_positional[10055:10052], addr_2513_6);

wire[27:0] addr_2514_6;

Selector_2 s2514_6(wires_628_5[2], addr_628_5, addr_positional[10059:10056], addr_2514_6);

wire[27:0] addr_2515_6;

Selector_2 s2515_6(wires_628_5[3], addr_628_5, addr_positional[10063:10060], addr_2515_6);

wire[27:0] addr_2516_6;

Selector_2 s2516_6(wires_629_5[0], addr_629_5, addr_positional[10067:10064], addr_2516_6);

wire[27:0] addr_2517_6;

Selector_2 s2517_6(wires_629_5[1], addr_629_5, addr_positional[10071:10068], addr_2517_6);

wire[27:0] addr_2518_6;

Selector_2 s2518_6(wires_629_5[2], addr_629_5, addr_positional[10075:10072], addr_2518_6);

wire[27:0] addr_2519_6;

Selector_2 s2519_6(wires_629_5[3], addr_629_5, addr_positional[10079:10076], addr_2519_6);

wire[27:0] addr_2520_6;

Selector_2 s2520_6(wires_630_5[0], addr_630_5, addr_positional[10083:10080], addr_2520_6);

wire[27:0] addr_2521_6;

Selector_2 s2521_6(wires_630_5[1], addr_630_5, addr_positional[10087:10084], addr_2521_6);

wire[27:0] addr_2522_6;

Selector_2 s2522_6(wires_630_5[2], addr_630_5, addr_positional[10091:10088], addr_2522_6);

wire[27:0] addr_2523_6;

Selector_2 s2523_6(wires_630_5[3], addr_630_5, addr_positional[10095:10092], addr_2523_6);

wire[27:0] addr_2524_6;

Selector_2 s2524_6(wires_631_5[0], addr_631_5, addr_positional[10099:10096], addr_2524_6);

wire[27:0] addr_2525_6;

Selector_2 s2525_6(wires_631_5[1], addr_631_5, addr_positional[10103:10100], addr_2525_6);

wire[27:0] addr_2526_6;

Selector_2 s2526_6(wires_631_5[2], addr_631_5, addr_positional[10107:10104], addr_2526_6);

wire[27:0] addr_2527_6;

Selector_2 s2527_6(wires_631_5[3], addr_631_5, addr_positional[10111:10108], addr_2527_6);

wire[27:0] addr_2528_6;

Selector_2 s2528_6(wires_632_5[0], addr_632_5, addr_positional[10115:10112], addr_2528_6);

wire[27:0] addr_2529_6;

Selector_2 s2529_6(wires_632_5[1], addr_632_5, addr_positional[10119:10116], addr_2529_6);

wire[27:0] addr_2530_6;

Selector_2 s2530_6(wires_632_5[2], addr_632_5, addr_positional[10123:10120], addr_2530_6);

wire[27:0] addr_2531_6;

Selector_2 s2531_6(wires_632_5[3], addr_632_5, addr_positional[10127:10124], addr_2531_6);

wire[27:0] addr_2532_6;

Selector_2 s2532_6(wires_633_5[0], addr_633_5, addr_positional[10131:10128], addr_2532_6);

wire[27:0] addr_2533_6;

Selector_2 s2533_6(wires_633_5[1], addr_633_5, addr_positional[10135:10132], addr_2533_6);

wire[27:0] addr_2534_6;

Selector_2 s2534_6(wires_633_5[2], addr_633_5, addr_positional[10139:10136], addr_2534_6);

wire[27:0] addr_2535_6;

Selector_2 s2535_6(wires_633_5[3], addr_633_5, addr_positional[10143:10140], addr_2535_6);

wire[27:0] addr_2536_6;

Selector_2 s2536_6(wires_634_5[0], addr_634_5, addr_positional[10147:10144], addr_2536_6);

wire[27:0] addr_2537_6;

Selector_2 s2537_6(wires_634_5[1], addr_634_5, addr_positional[10151:10148], addr_2537_6);

wire[27:0] addr_2538_6;

Selector_2 s2538_6(wires_634_5[2], addr_634_5, addr_positional[10155:10152], addr_2538_6);

wire[27:0] addr_2539_6;

Selector_2 s2539_6(wires_634_5[3], addr_634_5, addr_positional[10159:10156], addr_2539_6);

wire[27:0] addr_2540_6;

Selector_2 s2540_6(wires_635_5[0], addr_635_5, addr_positional[10163:10160], addr_2540_6);

wire[27:0] addr_2541_6;

Selector_2 s2541_6(wires_635_5[1], addr_635_5, addr_positional[10167:10164], addr_2541_6);

wire[27:0] addr_2542_6;

Selector_2 s2542_6(wires_635_5[2], addr_635_5, addr_positional[10171:10168], addr_2542_6);

wire[27:0] addr_2543_6;

Selector_2 s2543_6(wires_635_5[3], addr_635_5, addr_positional[10175:10172], addr_2543_6);

wire[27:0] addr_2544_6;

Selector_2 s2544_6(wires_636_5[0], addr_636_5, addr_positional[10179:10176], addr_2544_6);

wire[27:0] addr_2545_6;

Selector_2 s2545_6(wires_636_5[1], addr_636_5, addr_positional[10183:10180], addr_2545_6);

wire[27:0] addr_2546_6;

Selector_2 s2546_6(wires_636_5[2], addr_636_5, addr_positional[10187:10184], addr_2546_6);

wire[27:0] addr_2547_6;

Selector_2 s2547_6(wires_636_5[3], addr_636_5, addr_positional[10191:10188], addr_2547_6);

wire[27:0] addr_2548_6;

Selector_2 s2548_6(wires_637_5[0], addr_637_5, addr_positional[10195:10192], addr_2548_6);

wire[27:0] addr_2549_6;

Selector_2 s2549_6(wires_637_5[1], addr_637_5, addr_positional[10199:10196], addr_2549_6);

wire[27:0] addr_2550_6;

Selector_2 s2550_6(wires_637_5[2], addr_637_5, addr_positional[10203:10200], addr_2550_6);

wire[27:0] addr_2551_6;

Selector_2 s2551_6(wires_637_5[3], addr_637_5, addr_positional[10207:10204], addr_2551_6);

wire[27:0] addr_2552_6;

Selector_2 s2552_6(wires_638_5[0], addr_638_5, addr_positional[10211:10208], addr_2552_6);

wire[27:0] addr_2553_6;

Selector_2 s2553_6(wires_638_5[1], addr_638_5, addr_positional[10215:10212], addr_2553_6);

wire[27:0] addr_2554_6;

Selector_2 s2554_6(wires_638_5[2], addr_638_5, addr_positional[10219:10216], addr_2554_6);

wire[27:0] addr_2555_6;

Selector_2 s2555_6(wires_638_5[3], addr_638_5, addr_positional[10223:10220], addr_2555_6);

wire[27:0] addr_2556_6;

Selector_2 s2556_6(wires_639_5[0], addr_639_5, addr_positional[10227:10224], addr_2556_6);

wire[27:0] addr_2557_6;

Selector_2 s2557_6(wires_639_5[1], addr_639_5, addr_positional[10231:10228], addr_2557_6);

wire[27:0] addr_2558_6;

Selector_2 s2558_6(wires_639_5[2], addr_639_5, addr_positional[10235:10232], addr_2558_6);

wire[27:0] addr_2559_6;

Selector_2 s2559_6(wires_639_5[3], addr_639_5, addr_positional[10239:10236], addr_2559_6);

wire[27:0] addr_2560_6;

Selector_2 s2560_6(wires_640_5[0], addr_640_5, addr_positional[10243:10240], addr_2560_6);

wire[27:0] addr_2561_6;

Selector_2 s2561_6(wires_640_5[1], addr_640_5, addr_positional[10247:10244], addr_2561_6);

wire[27:0] addr_2562_6;

Selector_2 s2562_6(wires_640_5[2], addr_640_5, addr_positional[10251:10248], addr_2562_6);

wire[27:0] addr_2563_6;

Selector_2 s2563_6(wires_640_5[3], addr_640_5, addr_positional[10255:10252], addr_2563_6);

wire[27:0] addr_2564_6;

Selector_2 s2564_6(wires_641_5[0], addr_641_5, addr_positional[10259:10256], addr_2564_6);

wire[27:0] addr_2565_6;

Selector_2 s2565_6(wires_641_5[1], addr_641_5, addr_positional[10263:10260], addr_2565_6);

wire[27:0] addr_2566_6;

Selector_2 s2566_6(wires_641_5[2], addr_641_5, addr_positional[10267:10264], addr_2566_6);

wire[27:0] addr_2567_6;

Selector_2 s2567_6(wires_641_5[3], addr_641_5, addr_positional[10271:10268], addr_2567_6);

wire[27:0] addr_2568_6;

Selector_2 s2568_6(wires_642_5[0], addr_642_5, addr_positional[10275:10272], addr_2568_6);

wire[27:0] addr_2569_6;

Selector_2 s2569_6(wires_642_5[1], addr_642_5, addr_positional[10279:10276], addr_2569_6);

wire[27:0] addr_2570_6;

Selector_2 s2570_6(wires_642_5[2], addr_642_5, addr_positional[10283:10280], addr_2570_6);

wire[27:0] addr_2571_6;

Selector_2 s2571_6(wires_642_5[3], addr_642_5, addr_positional[10287:10284], addr_2571_6);

wire[27:0] addr_2572_6;

Selector_2 s2572_6(wires_643_5[0], addr_643_5, addr_positional[10291:10288], addr_2572_6);

wire[27:0] addr_2573_6;

Selector_2 s2573_6(wires_643_5[1], addr_643_5, addr_positional[10295:10292], addr_2573_6);

wire[27:0] addr_2574_6;

Selector_2 s2574_6(wires_643_5[2], addr_643_5, addr_positional[10299:10296], addr_2574_6);

wire[27:0] addr_2575_6;

Selector_2 s2575_6(wires_643_5[3], addr_643_5, addr_positional[10303:10300], addr_2575_6);

wire[27:0] addr_2576_6;

Selector_2 s2576_6(wires_644_5[0], addr_644_5, addr_positional[10307:10304], addr_2576_6);

wire[27:0] addr_2577_6;

Selector_2 s2577_6(wires_644_5[1], addr_644_5, addr_positional[10311:10308], addr_2577_6);

wire[27:0] addr_2578_6;

Selector_2 s2578_6(wires_644_5[2], addr_644_5, addr_positional[10315:10312], addr_2578_6);

wire[27:0] addr_2579_6;

Selector_2 s2579_6(wires_644_5[3], addr_644_5, addr_positional[10319:10316], addr_2579_6);

wire[27:0] addr_2580_6;

Selector_2 s2580_6(wires_645_5[0], addr_645_5, addr_positional[10323:10320], addr_2580_6);

wire[27:0] addr_2581_6;

Selector_2 s2581_6(wires_645_5[1], addr_645_5, addr_positional[10327:10324], addr_2581_6);

wire[27:0] addr_2582_6;

Selector_2 s2582_6(wires_645_5[2], addr_645_5, addr_positional[10331:10328], addr_2582_6);

wire[27:0] addr_2583_6;

Selector_2 s2583_6(wires_645_5[3], addr_645_5, addr_positional[10335:10332], addr_2583_6);

wire[27:0] addr_2584_6;

Selector_2 s2584_6(wires_646_5[0], addr_646_5, addr_positional[10339:10336], addr_2584_6);

wire[27:0] addr_2585_6;

Selector_2 s2585_6(wires_646_5[1], addr_646_5, addr_positional[10343:10340], addr_2585_6);

wire[27:0] addr_2586_6;

Selector_2 s2586_6(wires_646_5[2], addr_646_5, addr_positional[10347:10344], addr_2586_6);

wire[27:0] addr_2587_6;

Selector_2 s2587_6(wires_646_5[3], addr_646_5, addr_positional[10351:10348], addr_2587_6);

wire[27:0] addr_2588_6;

Selector_2 s2588_6(wires_647_5[0], addr_647_5, addr_positional[10355:10352], addr_2588_6);

wire[27:0] addr_2589_6;

Selector_2 s2589_6(wires_647_5[1], addr_647_5, addr_positional[10359:10356], addr_2589_6);

wire[27:0] addr_2590_6;

Selector_2 s2590_6(wires_647_5[2], addr_647_5, addr_positional[10363:10360], addr_2590_6);

wire[27:0] addr_2591_6;

Selector_2 s2591_6(wires_647_5[3], addr_647_5, addr_positional[10367:10364], addr_2591_6);

wire[27:0] addr_2592_6;

Selector_2 s2592_6(wires_648_5[0], addr_648_5, addr_positional[10371:10368], addr_2592_6);

wire[27:0] addr_2593_6;

Selector_2 s2593_6(wires_648_5[1], addr_648_5, addr_positional[10375:10372], addr_2593_6);

wire[27:0] addr_2594_6;

Selector_2 s2594_6(wires_648_5[2], addr_648_5, addr_positional[10379:10376], addr_2594_6);

wire[27:0] addr_2595_6;

Selector_2 s2595_6(wires_648_5[3], addr_648_5, addr_positional[10383:10380], addr_2595_6);

wire[27:0] addr_2596_6;

Selector_2 s2596_6(wires_649_5[0], addr_649_5, addr_positional[10387:10384], addr_2596_6);

wire[27:0] addr_2597_6;

Selector_2 s2597_6(wires_649_5[1], addr_649_5, addr_positional[10391:10388], addr_2597_6);

wire[27:0] addr_2598_6;

Selector_2 s2598_6(wires_649_5[2], addr_649_5, addr_positional[10395:10392], addr_2598_6);

wire[27:0] addr_2599_6;

Selector_2 s2599_6(wires_649_5[3], addr_649_5, addr_positional[10399:10396], addr_2599_6);

wire[27:0] addr_2600_6;

Selector_2 s2600_6(wires_650_5[0], addr_650_5, addr_positional[10403:10400], addr_2600_6);

wire[27:0] addr_2601_6;

Selector_2 s2601_6(wires_650_5[1], addr_650_5, addr_positional[10407:10404], addr_2601_6);

wire[27:0] addr_2602_6;

Selector_2 s2602_6(wires_650_5[2], addr_650_5, addr_positional[10411:10408], addr_2602_6);

wire[27:0] addr_2603_6;

Selector_2 s2603_6(wires_650_5[3], addr_650_5, addr_positional[10415:10412], addr_2603_6);

wire[27:0] addr_2604_6;

Selector_2 s2604_6(wires_651_5[0], addr_651_5, addr_positional[10419:10416], addr_2604_6);

wire[27:0] addr_2605_6;

Selector_2 s2605_6(wires_651_5[1], addr_651_5, addr_positional[10423:10420], addr_2605_6);

wire[27:0] addr_2606_6;

Selector_2 s2606_6(wires_651_5[2], addr_651_5, addr_positional[10427:10424], addr_2606_6);

wire[27:0] addr_2607_6;

Selector_2 s2607_6(wires_651_5[3], addr_651_5, addr_positional[10431:10428], addr_2607_6);

wire[27:0] addr_2608_6;

Selector_2 s2608_6(wires_652_5[0], addr_652_5, addr_positional[10435:10432], addr_2608_6);

wire[27:0] addr_2609_6;

Selector_2 s2609_6(wires_652_5[1], addr_652_5, addr_positional[10439:10436], addr_2609_6);

wire[27:0] addr_2610_6;

Selector_2 s2610_6(wires_652_5[2], addr_652_5, addr_positional[10443:10440], addr_2610_6);

wire[27:0] addr_2611_6;

Selector_2 s2611_6(wires_652_5[3], addr_652_5, addr_positional[10447:10444], addr_2611_6);

wire[27:0] addr_2612_6;

Selector_2 s2612_6(wires_653_5[0], addr_653_5, addr_positional[10451:10448], addr_2612_6);

wire[27:0] addr_2613_6;

Selector_2 s2613_6(wires_653_5[1], addr_653_5, addr_positional[10455:10452], addr_2613_6);

wire[27:0] addr_2614_6;

Selector_2 s2614_6(wires_653_5[2], addr_653_5, addr_positional[10459:10456], addr_2614_6);

wire[27:0] addr_2615_6;

Selector_2 s2615_6(wires_653_5[3], addr_653_5, addr_positional[10463:10460], addr_2615_6);

wire[27:0] addr_2616_6;

Selector_2 s2616_6(wires_654_5[0], addr_654_5, addr_positional[10467:10464], addr_2616_6);

wire[27:0] addr_2617_6;

Selector_2 s2617_6(wires_654_5[1], addr_654_5, addr_positional[10471:10468], addr_2617_6);

wire[27:0] addr_2618_6;

Selector_2 s2618_6(wires_654_5[2], addr_654_5, addr_positional[10475:10472], addr_2618_6);

wire[27:0] addr_2619_6;

Selector_2 s2619_6(wires_654_5[3], addr_654_5, addr_positional[10479:10476], addr_2619_6);

wire[27:0] addr_2620_6;

Selector_2 s2620_6(wires_655_5[0], addr_655_5, addr_positional[10483:10480], addr_2620_6);

wire[27:0] addr_2621_6;

Selector_2 s2621_6(wires_655_5[1], addr_655_5, addr_positional[10487:10484], addr_2621_6);

wire[27:0] addr_2622_6;

Selector_2 s2622_6(wires_655_5[2], addr_655_5, addr_positional[10491:10488], addr_2622_6);

wire[27:0] addr_2623_6;

Selector_2 s2623_6(wires_655_5[3], addr_655_5, addr_positional[10495:10492], addr_2623_6);

wire[27:0] addr_2624_6;

Selector_2 s2624_6(wires_656_5[0], addr_656_5, addr_positional[10499:10496], addr_2624_6);

wire[27:0] addr_2625_6;

Selector_2 s2625_6(wires_656_5[1], addr_656_5, addr_positional[10503:10500], addr_2625_6);

wire[27:0] addr_2626_6;

Selector_2 s2626_6(wires_656_5[2], addr_656_5, addr_positional[10507:10504], addr_2626_6);

wire[27:0] addr_2627_6;

Selector_2 s2627_6(wires_656_5[3], addr_656_5, addr_positional[10511:10508], addr_2627_6);

wire[27:0] addr_2628_6;

Selector_2 s2628_6(wires_657_5[0], addr_657_5, addr_positional[10515:10512], addr_2628_6);

wire[27:0] addr_2629_6;

Selector_2 s2629_6(wires_657_5[1], addr_657_5, addr_positional[10519:10516], addr_2629_6);

wire[27:0] addr_2630_6;

Selector_2 s2630_6(wires_657_5[2], addr_657_5, addr_positional[10523:10520], addr_2630_6);

wire[27:0] addr_2631_6;

Selector_2 s2631_6(wires_657_5[3], addr_657_5, addr_positional[10527:10524], addr_2631_6);

wire[27:0] addr_2632_6;

Selector_2 s2632_6(wires_658_5[0], addr_658_5, addr_positional[10531:10528], addr_2632_6);

wire[27:0] addr_2633_6;

Selector_2 s2633_6(wires_658_5[1], addr_658_5, addr_positional[10535:10532], addr_2633_6);

wire[27:0] addr_2634_6;

Selector_2 s2634_6(wires_658_5[2], addr_658_5, addr_positional[10539:10536], addr_2634_6);

wire[27:0] addr_2635_6;

Selector_2 s2635_6(wires_658_5[3], addr_658_5, addr_positional[10543:10540], addr_2635_6);

wire[27:0] addr_2636_6;

Selector_2 s2636_6(wires_659_5[0], addr_659_5, addr_positional[10547:10544], addr_2636_6);

wire[27:0] addr_2637_6;

Selector_2 s2637_6(wires_659_5[1], addr_659_5, addr_positional[10551:10548], addr_2637_6);

wire[27:0] addr_2638_6;

Selector_2 s2638_6(wires_659_5[2], addr_659_5, addr_positional[10555:10552], addr_2638_6);

wire[27:0] addr_2639_6;

Selector_2 s2639_6(wires_659_5[3], addr_659_5, addr_positional[10559:10556], addr_2639_6);

wire[27:0] addr_2640_6;

Selector_2 s2640_6(wires_660_5[0], addr_660_5, addr_positional[10563:10560], addr_2640_6);

wire[27:0] addr_2641_6;

Selector_2 s2641_6(wires_660_5[1], addr_660_5, addr_positional[10567:10564], addr_2641_6);

wire[27:0] addr_2642_6;

Selector_2 s2642_6(wires_660_5[2], addr_660_5, addr_positional[10571:10568], addr_2642_6);

wire[27:0] addr_2643_6;

Selector_2 s2643_6(wires_660_5[3], addr_660_5, addr_positional[10575:10572], addr_2643_6);

wire[27:0] addr_2644_6;

Selector_2 s2644_6(wires_661_5[0], addr_661_5, addr_positional[10579:10576], addr_2644_6);

wire[27:0] addr_2645_6;

Selector_2 s2645_6(wires_661_5[1], addr_661_5, addr_positional[10583:10580], addr_2645_6);

wire[27:0] addr_2646_6;

Selector_2 s2646_6(wires_661_5[2], addr_661_5, addr_positional[10587:10584], addr_2646_6);

wire[27:0] addr_2647_6;

Selector_2 s2647_6(wires_661_5[3], addr_661_5, addr_positional[10591:10588], addr_2647_6);

wire[27:0] addr_2648_6;

Selector_2 s2648_6(wires_662_5[0], addr_662_5, addr_positional[10595:10592], addr_2648_6);

wire[27:0] addr_2649_6;

Selector_2 s2649_6(wires_662_5[1], addr_662_5, addr_positional[10599:10596], addr_2649_6);

wire[27:0] addr_2650_6;

Selector_2 s2650_6(wires_662_5[2], addr_662_5, addr_positional[10603:10600], addr_2650_6);

wire[27:0] addr_2651_6;

Selector_2 s2651_6(wires_662_5[3], addr_662_5, addr_positional[10607:10604], addr_2651_6);

wire[27:0] addr_2652_6;

Selector_2 s2652_6(wires_663_5[0], addr_663_5, addr_positional[10611:10608], addr_2652_6);

wire[27:0] addr_2653_6;

Selector_2 s2653_6(wires_663_5[1], addr_663_5, addr_positional[10615:10612], addr_2653_6);

wire[27:0] addr_2654_6;

Selector_2 s2654_6(wires_663_5[2], addr_663_5, addr_positional[10619:10616], addr_2654_6);

wire[27:0] addr_2655_6;

Selector_2 s2655_6(wires_663_5[3], addr_663_5, addr_positional[10623:10620], addr_2655_6);

wire[27:0] addr_2656_6;

Selector_2 s2656_6(wires_664_5[0], addr_664_5, addr_positional[10627:10624], addr_2656_6);

wire[27:0] addr_2657_6;

Selector_2 s2657_6(wires_664_5[1], addr_664_5, addr_positional[10631:10628], addr_2657_6);

wire[27:0] addr_2658_6;

Selector_2 s2658_6(wires_664_5[2], addr_664_5, addr_positional[10635:10632], addr_2658_6);

wire[27:0] addr_2659_6;

Selector_2 s2659_6(wires_664_5[3], addr_664_5, addr_positional[10639:10636], addr_2659_6);

wire[27:0] addr_2660_6;

Selector_2 s2660_6(wires_665_5[0], addr_665_5, addr_positional[10643:10640], addr_2660_6);

wire[27:0] addr_2661_6;

Selector_2 s2661_6(wires_665_5[1], addr_665_5, addr_positional[10647:10644], addr_2661_6);

wire[27:0] addr_2662_6;

Selector_2 s2662_6(wires_665_5[2], addr_665_5, addr_positional[10651:10648], addr_2662_6);

wire[27:0] addr_2663_6;

Selector_2 s2663_6(wires_665_5[3], addr_665_5, addr_positional[10655:10652], addr_2663_6);

wire[27:0] addr_2664_6;

Selector_2 s2664_6(wires_666_5[0], addr_666_5, addr_positional[10659:10656], addr_2664_6);

wire[27:0] addr_2665_6;

Selector_2 s2665_6(wires_666_5[1], addr_666_5, addr_positional[10663:10660], addr_2665_6);

wire[27:0] addr_2666_6;

Selector_2 s2666_6(wires_666_5[2], addr_666_5, addr_positional[10667:10664], addr_2666_6);

wire[27:0] addr_2667_6;

Selector_2 s2667_6(wires_666_5[3], addr_666_5, addr_positional[10671:10668], addr_2667_6);

wire[27:0] addr_2668_6;

Selector_2 s2668_6(wires_667_5[0], addr_667_5, addr_positional[10675:10672], addr_2668_6);

wire[27:0] addr_2669_6;

Selector_2 s2669_6(wires_667_5[1], addr_667_5, addr_positional[10679:10676], addr_2669_6);

wire[27:0] addr_2670_6;

Selector_2 s2670_6(wires_667_5[2], addr_667_5, addr_positional[10683:10680], addr_2670_6);

wire[27:0] addr_2671_6;

Selector_2 s2671_6(wires_667_5[3], addr_667_5, addr_positional[10687:10684], addr_2671_6);

wire[27:0] addr_2672_6;

Selector_2 s2672_6(wires_668_5[0], addr_668_5, addr_positional[10691:10688], addr_2672_6);

wire[27:0] addr_2673_6;

Selector_2 s2673_6(wires_668_5[1], addr_668_5, addr_positional[10695:10692], addr_2673_6);

wire[27:0] addr_2674_6;

Selector_2 s2674_6(wires_668_5[2], addr_668_5, addr_positional[10699:10696], addr_2674_6);

wire[27:0] addr_2675_6;

Selector_2 s2675_6(wires_668_5[3], addr_668_5, addr_positional[10703:10700], addr_2675_6);

wire[27:0] addr_2676_6;

Selector_2 s2676_6(wires_669_5[0], addr_669_5, addr_positional[10707:10704], addr_2676_6);

wire[27:0] addr_2677_6;

Selector_2 s2677_6(wires_669_5[1], addr_669_5, addr_positional[10711:10708], addr_2677_6);

wire[27:0] addr_2678_6;

Selector_2 s2678_6(wires_669_5[2], addr_669_5, addr_positional[10715:10712], addr_2678_6);

wire[27:0] addr_2679_6;

Selector_2 s2679_6(wires_669_5[3], addr_669_5, addr_positional[10719:10716], addr_2679_6);

wire[27:0] addr_2680_6;

Selector_2 s2680_6(wires_670_5[0], addr_670_5, addr_positional[10723:10720], addr_2680_6);

wire[27:0] addr_2681_6;

Selector_2 s2681_6(wires_670_5[1], addr_670_5, addr_positional[10727:10724], addr_2681_6);

wire[27:0] addr_2682_6;

Selector_2 s2682_6(wires_670_5[2], addr_670_5, addr_positional[10731:10728], addr_2682_6);

wire[27:0] addr_2683_6;

Selector_2 s2683_6(wires_670_5[3], addr_670_5, addr_positional[10735:10732], addr_2683_6);

wire[27:0] addr_2684_6;

Selector_2 s2684_6(wires_671_5[0], addr_671_5, addr_positional[10739:10736], addr_2684_6);

wire[27:0] addr_2685_6;

Selector_2 s2685_6(wires_671_5[1], addr_671_5, addr_positional[10743:10740], addr_2685_6);

wire[27:0] addr_2686_6;

Selector_2 s2686_6(wires_671_5[2], addr_671_5, addr_positional[10747:10744], addr_2686_6);

wire[27:0] addr_2687_6;

Selector_2 s2687_6(wires_671_5[3], addr_671_5, addr_positional[10751:10748], addr_2687_6);

wire[27:0] addr_2688_6;

Selector_2 s2688_6(wires_672_5[0], addr_672_5, addr_positional[10755:10752], addr_2688_6);

wire[27:0] addr_2689_6;

Selector_2 s2689_6(wires_672_5[1], addr_672_5, addr_positional[10759:10756], addr_2689_6);

wire[27:0] addr_2690_6;

Selector_2 s2690_6(wires_672_5[2], addr_672_5, addr_positional[10763:10760], addr_2690_6);

wire[27:0] addr_2691_6;

Selector_2 s2691_6(wires_672_5[3], addr_672_5, addr_positional[10767:10764], addr_2691_6);

wire[27:0] addr_2692_6;

Selector_2 s2692_6(wires_673_5[0], addr_673_5, addr_positional[10771:10768], addr_2692_6);

wire[27:0] addr_2693_6;

Selector_2 s2693_6(wires_673_5[1], addr_673_5, addr_positional[10775:10772], addr_2693_6);

wire[27:0] addr_2694_6;

Selector_2 s2694_6(wires_673_5[2], addr_673_5, addr_positional[10779:10776], addr_2694_6);

wire[27:0] addr_2695_6;

Selector_2 s2695_6(wires_673_5[3], addr_673_5, addr_positional[10783:10780], addr_2695_6);

wire[27:0] addr_2696_6;

Selector_2 s2696_6(wires_674_5[0], addr_674_5, addr_positional[10787:10784], addr_2696_6);

wire[27:0] addr_2697_6;

Selector_2 s2697_6(wires_674_5[1], addr_674_5, addr_positional[10791:10788], addr_2697_6);

wire[27:0] addr_2698_6;

Selector_2 s2698_6(wires_674_5[2], addr_674_5, addr_positional[10795:10792], addr_2698_6);

wire[27:0] addr_2699_6;

Selector_2 s2699_6(wires_674_5[3], addr_674_5, addr_positional[10799:10796], addr_2699_6);

wire[27:0] addr_2700_6;

Selector_2 s2700_6(wires_675_5[0], addr_675_5, addr_positional[10803:10800], addr_2700_6);

wire[27:0] addr_2701_6;

Selector_2 s2701_6(wires_675_5[1], addr_675_5, addr_positional[10807:10804], addr_2701_6);

wire[27:0] addr_2702_6;

Selector_2 s2702_6(wires_675_5[2], addr_675_5, addr_positional[10811:10808], addr_2702_6);

wire[27:0] addr_2703_6;

Selector_2 s2703_6(wires_675_5[3], addr_675_5, addr_positional[10815:10812], addr_2703_6);

wire[27:0] addr_2704_6;

Selector_2 s2704_6(wires_676_5[0], addr_676_5, addr_positional[10819:10816], addr_2704_6);

wire[27:0] addr_2705_6;

Selector_2 s2705_6(wires_676_5[1], addr_676_5, addr_positional[10823:10820], addr_2705_6);

wire[27:0] addr_2706_6;

Selector_2 s2706_6(wires_676_5[2], addr_676_5, addr_positional[10827:10824], addr_2706_6);

wire[27:0] addr_2707_6;

Selector_2 s2707_6(wires_676_5[3], addr_676_5, addr_positional[10831:10828], addr_2707_6);

wire[27:0] addr_2708_6;

Selector_2 s2708_6(wires_677_5[0], addr_677_5, addr_positional[10835:10832], addr_2708_6);

wire[27:0] addr_2709_6;

Selector_2 s2709_6(wires_677_5[1], addr_677_5, addr_positional[10839:10836], addr_2709_6);

wire[27:0] addr_2710_6;

Selector_2 s2710_6(wires_677_5[2], addr_677_5, addr_positional[10843:10840], addr_2710_6);

wire[27:0] addr_2711_6;

Selector_2 s2711_6(wires_677_5[3], addr_677_5, addr_positional[10847:10844], addr_2711_6);

wire[27:0] addr_2712_6;

Selector_2 s2712_6(wires_678_5[0], addr_678_5, addr_positional[10851:10848], addr_2712_6);

wire[27:0] addr_2713_6;

Selector_2 s2713_6(wires_678_5[1], addr_678_5, addr_positional[10855:10852], addr_2713_6);

wire[27:0] addr_2714_6;

Selector_2 s2714_6(wires_678_5[2], addr_678_5, addr_positional[10859:10856], addr_2714_6);

wire[27:0] addr_2715_6;

Selector_2 s2715_6(wires_678_5[3], addr_678_5, addr_positional[10863:10860], addr_2715_6);

wire[27:0] addr_2716_6;

Selector_2 s2716_6(wires_679_5[0], addr_679_5, addr_positional[10867:10864], addr_2716_6);

wire[27:0] addr_2717_6;

Selector_2 s2717_6(wires_679_5[1], addr_679_5, addr_positional[10871:10868], addr_2717_6);

wire[27:0] addr_2718_6;

Selector_2 s2718_6(wires_679_5[2], addr_679_5, addr_positional[10875:10872], addr_2718_6);

wire[27:0] addr_2719_6;

Selector_2 s2719_6(wires_679_5[3], addr_679_5, addr_positional[10879:10876], addr_2719_6);

wire[27:0] addr_2720_6;

Selector_2 s2720_6(wires_680_5[0], addr_680_5, addr_positional[10883:10880], addr_2720_6);

wire[27:0] addr_2721_6;

Selector_2 s2721_6(wires_680_5[1], addr_680_5, addr_positional[10887:10884], addr_2721_6);

wire[27:0] addr_2722_6;

Selector_2 s2722_6(wires_680_5[2], addr_680_5, addr_positional[10891:10888], addr_2722_6);

wire[27:0] addr_2723_6;

Selector_2 s2723_6(wires_680_5[3], addr_680_5, addr_positional[10895:10892], addr_2723_6);

wire[27:0] addr_2724_6;

Selector_2 s2724_6(wires_681_5[0], addr_681_5, addr_positional[10899:10896], addr_2724_6);

wire[27:0] addr_2725_6;

Selector_2 s2725_6(wires_681_5[1], addr_681_5, addr_positional[10903:10900], addr_2725_6);

wire[27:0] addr_2726_6;

Selector_2 s2726_6(wires_681_5[2], addr_681_5, addr_positional[10907:10904], addr_2726_6);

wire[27:0] addr_2727_6;

Selector_2 s2727_6(wires_681_5[3], addr_681_5, addr_positional[10911:10908], addr_2727_6);

wire[27:0] addr_2728_6;

Selector_2 s2728_6(wires_682_5[0], addr_682_5, addr_positional[10915:10912], addr_2728_6);

wire[27:0] addr_2729_6;

Selector_2 s2729_6(wires_682_5[1], addr_682_5, addr_positional[10919:10916], addr_2729_6);

wire[27:0] addr_2730_6;

Selector_2 s2730_6(wires_682_5[2], addr_682_5, addr_positional[10923:10920], addr_2730_6);

wire[27:0] addr_2731_6;

Selector_2 s2731_6(wires_682_5[3], addr_682_5, addr_positional[10927:10924], addr_2731_6);

wire[27:0] addr_2732_6;

Selector_2 s2732_6(wires_683_5[0], addr_683_5, addr_positional[10931:10928], addr_2732_6);

wire[27:0] addr_2733_6;

Selector_2 s2733_6(wires_683_5[1], addr_683_5, addr_positional[10935:10932], addr_2733_6);

wire[27:0] addr_2734_6;

Selector_2 s2734_6(wires_683_5[2], addr_683_5, addr_positional[10939:10936], addr_2734_6);

wire[27:0] addr_2735_6;

Selector_2 s2735_6(wires_683_5[3], addr_683_5, addr_positional[10943:10940], addr_2735_6);

wire[27:0] addr_2736_6;

Selector_2 s2736_6(wires_684_5[0], addr_684_5, addr_positional[10947:10944], addr_2736_6);

wire[27:0] addr_2737_6;

Selector_2 s2737_6(wires_684_5[1], addr_684_5, addr_positional[10951:10948], addr_2737_6);

wire[27:0] addr_2738_6;

Selector_2 s2738_6(wires_684_5[2], addr_684_5, addr_positional[10955:10952], addr_2738_6);

wire[27:0] addr_2739_6;

Selector_2 s2739_6(wires_684_5[3], addr_684_5, addr_positional[10959:10956], addr_2739_6);

wire[27:0] addr_2740_6;

Selector_2 s2740_6(wires_685_5[0], addr_685_5, addr_positional[10963:10960], addr_2740_6);

wire[27:0] addr_2741_6;

Selector_2 s2741_6(wires_685_5[1], addr_685_5, addr_positional[10967:10964], addr_2741_6);

wire[27:0] addr_2742_6;

Selector_2 s2742_6(wires_685_5[2], addr_685_5, addr_positional[10971:10968], addr_2742_6);

wire[27:0] addr_2743_6;

Selector_2 s2743_6(wires_685_5[3], addr_685_5, addr_positional[10975:10972], addr_2743_6);

wire[27:0] addr_2744_6;

Selector_2 s2744_6(wires_686_5[0], addr_686_5, addr_positional[10979:10976], addr_2744_6);

wire[27:0] addr_2745_6;

Selector_2 s2745_6(wires_686_5[1], addr_686_5, addr_positional[10983:10980], addr_2745_6);

wire[27:0] addr_2746_6;

Selector_2 s2746_6(wires_686_5[2], addr_686_5, addr_positional[10987:10984], addr_2746_6);

wire[27:0] addr_2747_6;

Selector_2 s2747_6(wires_686_5[3], addr_686_5, addr_positional[10991:10988], addr_2747_6);

wire[27:0] addr_2748_6;

Selector_2 s2748_6(wires_687_5[0], addr_687_5, addr_positional[10995:10992], addr_2748_6);

wire[27:0] addr_2749_6;

Selector_2 s2749_6(wires_687_5[1], addr_687_5, addr_positional[10999:10996], addr_2749_6);

wire[27:0] addr_2750_6;

Selector_2 s2750_6(wires_687_5[2], addr_687_5, addr_positional[11003:11000], addr_2750_6);

wire[27:0] addr_2751_6;

Selector_2 s2751_6(wires_687_5[3], addr_687_5, addr_positional[11007:11004], addr_2751_6);

wire[27:0] addr_2752_6;

Selector_2 s2752_6(wires_688_5[0], addr_688_5, addr_positional[11011:11008], addr_2752_6);

wire[27:0] addr_2753_6;

Selector_2 s2753_6(wires_688_5[1], addr_688_5, addr_positional[11015:11012], addr_2753_6);

wire[27:0] addr_2754_6;

Selector_2 s2754_6(wires_688_5[2], addr_688_5, addr_positional[11019:11016], addr_2754_6);

wire[27:0] addr_2755_6;

Selector_2 s2755_6(wires_688_5[3], addr_688_5, addr_positional[11023:11020], addr_2755_6);

wire[27:0] addr_2756_6;

Selector_2 s2756_6(wires_689_5[0], addr_689_5, addr_positional[11027:11024], addr_2756_6);

wire[27:0] addr_2757_6;

Selector_2 s2757_6(wires_689_5[1], addr_689_5, addr_positional[11031:11028], addr_2757_6);

wire[27:0] addr_2758_6;

Selector_2 s2758_6(wires_689_5[2], addr_689_5, addr_positional[11035:11032], addr_2758_6);

wire[27:0] addr_2759_6;

Selector_2 s2759_6(wires_689_5[3], addr_689_5, addr_positional[11039:11036], addr_2759_6);

wire[27:0] addr_2760_6;

Selector_2 s2760_6(wires_690_5[0], addr_690_5, addr_positional[11043:11040], addr_2760_6);

wire[27:0] addr_2761_6;

Selector_2 s2761_6(wires_690_5[1], addr_690_5, addr_positional[11047:11044], addr_2761_6);

wire[27:0] addr_2762_6;

Selector_2 s2762_6(wires_690_5[2], addr_690_5, addr_positional[11051:11048], addr_2762_6);

wire[27:0] addr_2763_6;

Selector_2 s2763_6(wires_690_5[3], addr_690_5, addr_positional[11055:11052], addr_2763_6);

wire[27:0] addr_2764_6;

Selector_2 s2764_6(wires_691_5[0], addr_691_5, addr_positional[11059:11056], addr_2764_6);

wire[27:0] addr_2765_6;

Selector_2 s2765_6(wires_691_5[1], addr_691_5, addr_positional[11063:11060], addr_2765_6);

wire[27:0] addr_2766_6;

Selector_2 s2766_6(wires_691_5[2], addr_691_5, addr_positional[11067:11064], addr_2766_6);

wire[27:0] addr_2767_6;

Selector_2 s2767_6(wires_691_5[3], addr_691_5, addr_positional[11071:11068], addr_2767_6);

wire[27:0] addr_2768_6;

Selector_2 s2768_6(wires_692_5[0], addr_692_5, addr_positional[11075:11072], addr_2768_6);

wire[27:0] addr_2769_6;

Selector_2 s2769_6(wires_692_5[1], addr_692_5, addr_positional[11079:11076], addr_2769_6);

wire[27:0] addr_2770_6;

Selector_2 s2770_6(wires_692_5[2], addr_692_5, addr_positional[11083:11080], addr_2770_6);

wire[27:0] addr_2771_6;

Selector_2 s2771_6(wires_692_5[3], addr_692_5, addr_positional[11087:11084], addr_2771_6);

wire[27:0] addr_2772_6;

Selector_2 s2772_6(wires_693_5[0], addr_693_5, addr_positional[11091:11088], addr_2772_6);

wire[27:0] addr_2773_6;

Selector_2 s2773_6(wires_693_5[1], addr_693_5, addr_positional[11095:11092], addr_2773_6);

wire[27:0] addr_2774_6;

Selector_2 s2774_6(wires_693_5[2], addr_693_5, addr_positional[11099:11096], addr_2774_6);

wire[27:0] addr_2775_6;

Selector_2 s2775_6(wires_693_5[3], addr_693_5, addr_positional[11103:11100], addr_2775_6);

wire[27:0] addr_2776_6;

Selector_2 s2776_6(wires_694_5[0], addr_694_5, addr_positional[11107:11104], addr_2776_6);

wire[27:0] addr_2777_6;

Selector_2 s2777_6(wires_694_5[1], addr_694_5, addr_positional[11111:11108], addr_2777_6);

wire[27:0] addr_2778_6;

Selector_2 s2778_6(wires_694_5[2], addr_694_5, addr_positional[11115:11112], addr_2778_6);

wire[27:0] addr_2779_6;

Selector_2 s2779_6(wires_694_5[3], addr_694_5, addr_positional[11119:11116], addr_2779_6);

wire[27:0] addr_2780_6;

Selector_2 s2780_6(wires_695_5[0], addr_695_5, addr_positional[11123:11120], addr_2780_6);

wire[27:0] addr_2781_6;

Selector_2 s2781_6(wires_695_5[1], addr_695_5, addr_positional[11127:11124], addr_2781_6);

wire[27:0] addr_2782_6;

Selector_2 s2782_6(wires_695_5[2], addr_695_5, addr_positional[11131:11128], addr_2782_6);

wire[27:0] addr_2783_6;

Selector_2 s2783_6(wires_695_5[3], addr_695_5, addr_positional[11135:11132], addr_2783_6);

wire[27:0] addr_2784_6;

Selector_2 s2784_6(wires_696_5[0], addr_696_5, addr_positional[11139:11136], addr_2784_6);

wire[27:0] addr_2785_6;

Selector_2 s2785_6(wires_696_5[1], addr_696_5, addr_positional[11143:11140], addr_2785_6);

wire[27:0] addr_2786_6;

Selector_2 s2786_6(wires_696_5[2], addr_696_5, addr_positional[11147:11144], addr_2786_6);

wire[27:0] addr_2787_6;

Selector_2 s2787_6(wires_696_5[3], addr_696_5, addr_positional[11151:11148], addr_2787_6);

wire[27:0] addr_2788_6;

Selector_2 s2788_6(wires_697_5[0], addr_697_5, addr_positional[11155:11152], addr_2788_6);

wire[27:0] addr_2789_6;

Selector_2 s2789_6(wires_697_5[1], addr_697_5, addr_positional[11159:11156], addr_2789_6);

wire[27:0] addr_2790_6;

Selector_2 s2790_6(wires_697_5[2], addr_697_5, addr_positional[11163:11160], addr_2790_6);

wire[27:0] addr_2791_6;

Selector_2 s2791_6(wires_697_5[3], addr_697_5, addr_positional[11167:11164], addr_2791_6);

wire[27:0] addr_2792_6;

Selector_2 s2792_6(wires_698_5[0], addr_698_5, addr_positional[11171:11168], addr_2792_6);

wire[27:0] addr_2793_6;

Selector_2 s2793_6(wires_698_5[1], addr_698_5, addr_positional[11175:11172], addr_2793_6);

wire[27:0] addr_2794_6;

Selector_2 s2794_6(wires_698_5[2], addr_698_5, addr_positional[11179:11176], addr_2794_6);

wire[27:0] addr_2795_6;

Selector_2 s2795_6(wires_698_5[3], addr_698_5, addr_positional[11183:11180], addr_2795_6);

wire[27:0] addr_2796_6;

Selector_2 s2796_6(wires_699_5[0], addr_699_5, addr_positional[11187:11184], addr_2796_6);

wire[27:0] addr_2797_6;

Selector_2 s2797_6(wires_699_5[1], addr_699_5, addr_positional[11191:11188], addr_2797_6);

wire[27:0] addr_2798_6;

Selector_2 s2798_6(wires_699_5[2], addr_699_5, addr_positional[11195:11192], addr_2798_6);

wire[27:0] addr_2799_6;

Selector_2 s2799_6(wires_699_5[3], addr_699_5, addr_positional[11199:11196], addr_2799_6);

wire[27:0] addr_2800_6;

Selector_2 s2800_6(wires_700_5[0], addr_700_5, addr_positional[11203:11200], addr_2800_6);

wire[27:0] addr_2801_6;

Selector_2 s2801_6(wires_700_5[1], addr_700_5, addr_positional[11207:11204], addr_2801_6);

wire[27:0] addr_2802_6;

Selector_2 s2802_6(wires_700_5[2], addr_700_5, addr_positional[11211:11208], addr_2802_6);

wire[27:0] addr_2803_6;

Selector_2 s2803_6(wires_700_5[3], addr_700_5, addr_positional[11215:11212], addr_2803_6);

wire[27:0] addr_2804_6;

Selector_2 s2804_6(wires_701_5[0], addr_701_5, addr_positional[11219:11216], addr_2804_6);

wire[27:0] addr_2805_6;

Selector_2 s2805_6(wires_701_5[1], addr_701_5, addr_positional[11223:11220], addr_2805_6);

wire[27:0] addr_2806_6;

Selector_2 s2806_6(wires_701_5[2], addr_701_5, addr_positional[11227:11224], addr_2806_6);

wire[27:0] addr_2807_6;

Selector_2 s2807_6(wires_701_5[3], addr_701_5, addr_positional[11231:11228], addr_2807_6);

wire[27:0] addr_2808_6;

Selector_2 s2808_6(wires_702_5[0], addr_702_5, addr_positional[11235:11232], addr_2808_6);

wire[27:0] addr_2809_6;

Selector_2 s2809_6(wires_702_5[1], addr_702_5, addr_positional[11239:11236], addr_2809_6);

wire[27:0] addr_2810_6;

Selector_2 s2810_6(wires_702_5[2], addr_702_5, addr_positional[11243:11240], addr_2810_6);

wire[27:0] addr_2811_6;

Selector_2 s2811_6(wires_702_5[3], addr_702_5, addr_positional[11247:11244], addr_2811_6);

wire[27:0] addr_2812_6;

Selector_2 s2812_6(wires_703_5[0], addr_703_5, addr_positional[11251:11248], addr_2812_6);

wire[27:0] addr_2813_6;

Selector_2 s2813_6(wires_703_5[1], addr_703_5, addr_positional[11255:11252], addr_2813_6);

wire[27:0] addr_2814_6;

Selector_2 s2814_6(wires_703_5[2], addr_703_5, addr_positional[11259:11256], addr_2814_6);

wire[27:0] addr_2815_6;

Selector_2 s2815_6(wires_703_5[3], addr_703_5, addr_positional[11263:11260], addr_2815_6);

wire[27:0] addr_2816_6;

Selector_2 s2816_6(wires_704_5[0], addr_704_5, addr_positional[11267:11264], addr_2816_6);

wire[27:0] addr_2817_6;

Selector_2 s2817_6(wires_704_5[1], addr_704_5, addr_positional[11271:11268], addr_2817_6);

wire[27:0] addr_2818_6;

Selector_2 s2818_6(wires_704_5[2], addr_704_5, addr_positional[11275:11272], addr_2818_6);

wire[27:0] addr_2819_6;

Selector_2 s2819_6(wires_704_5[3], addr_704_5, addr_positional[11279:11276], addr_2819_6);

wire[27:0] addr_2820_6;

Selector_2 s2820_6(wires_705_5[0], addr_705_5, addr_positional[11283:11280], addr_2820_6);

wire[27:0] addr_2821_6;

Selector_2 s2821_6(wires_705_5[1], addr_705_5, addr_positional[11287:11284], addr_2821_6);

wire[27:0] addr_2822_6;

Selector_2 s2822_6(wires_705_5[2], addr_705_5, addr_positional[11291:11288], addr_2822_6);

wire[27:0] addr_2823_6;

Selector_2 s2823_6(wires_705_5[3], addr_705_5, addr_positional[11295:11292], addr_2823_6);

wire[27:0] addr_2824_6;

Selector_2 s2824_6(wires_706_5[0], addr_706_5, addr_positional[11299:11296], addr_2824_6);

wire[27:0] addr_2825_6;

Selector_2 s2825_6(wires_706_5[1], addr_706_5, addr_positional[11303:11300], addr_2825_6);

wire[27:0] addr_2826_6;

Selector_2 s2826_6(wires_706_5[2], addr_706_5, addr_positional[11307:11304], addr_2826_6);

wire[27:0] addr_2827_6;

Selector_2 s2827_6(wires_706_5[3], addr_706_5, addr_positional[11311:11308], addr_2827_6);

wire[27:0] addr_2828_6;

Selector_2 s2828_6(wires_707_5[0], addr_707_5, addr_positional[11315:11312], addr_2828_6);

wire[27:0] addr_2829_6;

Selector_2 s2829_6(wires_707_5[1], addr_707_5, addr_positional[11319:11316], addr_2829_6);

wire[27:0] addr_2830_6;

Selector_2 s2830_6(wires_707_5[2], addr_707_5, addr_positional[11323:11320], addr_2830_6);

wire[27:0] addr_2831_6;

Selector_2 s2831_6(wires_707_5[3], addr_707_5, addr_positional[11327:11324], addr_2831_6);

wire[27:0] addr_2832_6;

Selector_2 s2832_6(wires_708_5[0], addr_708_5, addr_positional[11331:11328], addr_2832_6);

wire[27:0] addr_2833_6;

Selector_2 s2833_6(wires_708_5[1], addr_708_5, addr_positional[11335:11332], addr_2833_6);

wire[27:0] addr_2834_6;

Selector_2 s2834_6(wires_708_5[2], addr_708_5, addr_positional[11339:11336], addr_2834_6);

wire[27:0] addr_2835_6;

Selector_2 s2835_6(wires_708_5[3], addr_708_5, addr_positional[11343:11340], addr_2835_6);

wire[27:0] addr_2836_6;

Selector_2 s2836_6(wires_709_5[0], addr_709_5, addr_positional[11347:11344], addr_2836_6);

wire[27:0] addr_2837_6;

Selector_2 s2837_6(wires_709_5[1], addr_709_5, addr_positional[11351:11348], addr_2837_6);

wire[27:0] addr_2838_6;

Selector_2 s2838_6(wires_709_5[2], addr_709_5, addr_positional[11355:11352], addr_2838_6);

wire[27:0] addr_2839_6;

Selector_2 s2839_6(wires_709_5[3], addr_709_5, addr_positional[11359:11356], addr_2839_6);

wire[27:0] addr_2840_6;

Selector_2 s2840_6(wires_710_5[0], addr_710_5, addr_positional[11363:11360], addr_2840_6);

wire[27:0] addr_2841_6;

Selector_2 s2841_6(wires_710_5[1], addr_710_5, addr_positional[11367:11364], addr_2841_6);

wire[27:0] addr_2842_6;

Selector_2 s2842_6(wires_710_5[2], addr_710_5, addr_positional[11371:11368], addr_2842_6);

wire[27:0] addr_2843_6;

Selector_2 s2843_6(wires_710_5[3], addr_710_5, addr_positional[11375:11372], addr_2843_6);

wire[27:0] addr_2844_6;

Selector_2 s2844_6(wires_711_5[0], addr_711_5, addr_positional[11379:11376], addr_2844_6);

wire[27:0] addr_2845_6;

Selector_2 s2845_6(wires_711_5[1], addr_711_5, addr_positional[11383:11380], addr_2845_6);

wire[27:0] addr_2846_6;

Selector_2 s2846_6(wires_711_5[2], addr_711_5, addr_positional[11387:11384], addr_2846_6);

wire[27:0] addr_2847_6;

Selector_2 s2847_6(wires_711_5[3], addr_711_5, addr_positional[11391:11388], addr_2847_6);

wire[27:0] addr_2848_6;

Selector_2 s2848_6(wires_712_5[0], addr_712_5, addr_positional[11395:11392], addr_2848_6);

wire[27:0] addr_2849_6;

Selector_2 s2849_6(wires_712_5[1], addr_712_5, addr_positional[11399:11396], addr_2849_6);

wire[27:0] addr_2850_6;

Selector_2 s2850_6(wires_712_5[2], addr_712_5, addr_positional[11403:11400], addr_2850_6);

wire[27:0] addr_2851_6;

Selector_2 s2851_6(wires_712_5[3], addr_712_5, addr_positional[11407:11404], addr_2851_6);

wire[27:0] addr_2852_6;

Selector_2 s2852_6(wires_713_5[0], addr_713_5, addr_positional[11411:11408], addr_2852_6);

wire[27:0] addr_2853_6;

Selector_2 s2853_6(wires_713_5[1], addr_713_5, addr_positional[11415:11412], addr_2853_6);

wire[27:0] addr_2854_6;

Selector_2 s2854_6(wires_713_5[2], addr_713_5, addr_positional[11419:11416], addr_2854_6);

wire[27:0] addr_2855_6;

Selector_2 s2855_6(wires_713_5[3], addr_713_5, addr_positional[11423:11420], addr_2855_6);

wire[27:0] addr_2856_6;

Selector_2 s2856_6(wires_714_5[0], addr_714_5, addr_positional[11427:11424], addr_2856_6);

wire[27:0] addr_2857_6;

Selector_2 s2857_6(wires_714_5[1], addr_714_5, addr_positional[11431:11428], addr_2857_6);

wire[27:0] addr_2858_6;

Selector_2 s2858_6(wires_714_5[2], addr_714_5, addr_positional[11435:11432], addr_2858_6);

wire[27:0] addr_2859_6;

Selector_2 s2859_6(wires_714_5[3], addr_714_5, addr_positional[11439:11436], addr_2859_6);

wire[27:0] addr_2860_6;

Selector_2 s2860_6(wires_715_5[0], addr_715_5, addr_positional[11443:11440], addr_2860_6);

wire[27:0] addr_2861_6;

Selector_2 s2861_6(wires_715_5[1], addr_715_5, addr_positional[11447:11444], addr_2861_6);

wire[27:0] addr_2862_6;

Selector_2 s2862_6(wires_715_5[2], addr_715_5, addr_positional[11451:11448], addr_2862_6);

wire[27:0] addr_2863_6;

Selector_2 s2863_6(wires_715_5[3], addr_715_5, addr_positional[11455:11452], addr_2863_6);

wire[27:0] addr_2864_6;

Selector_2 s2864_6(wires_716_5[0], addr_716_5, addr_positional[11459:11456], addr_2864_6);

wire[27:0] addr_2865_6;

Selector_2 s2865_6(wires_716_5[1], addr_716_5, addr_positional[11463:11460], addr_2865_6);

wire[27:0] addr_2866_6;

Selector_2 s2866_6(wires_716_5[2], addr_716_5, addr_positional[11467:11464], addr_2866_6);

wire[27:0] addr_2867_6;

Selector_2 s2867_6(wires_716_5[3], addr_716_5, addr_positional[11471:11468], addr_2867_6);

wire[27:0] addr_2868_6;

Selector_2 s2868_6(wires_717_5[0], addr_717_5, addr_positional[11475:11472], addr_2868_6);

wire[27:0] addr_2869_6;

Selector_2 s2869_6(wires_717_5[1], addr_717_5, addr_positional[11479:11476], addr_2869_6);

wire[27:0] addr_2870_6;

Selector_2 s2870_6(wires_717_5[2], addr_717_5, addr_positional[11483:11480], addr_2870_6);

wire[27:0] addr_2871_6;

Selector_2 s2871_6(wires_717_5[3], addr_717_5, addr_positional[11487:11484], addr_2871_6);

wire[27:0] addr_2872_6;

Selector_2 s2872_6(wires_718_5[0], addr_718_5, addr_positional[11491:11488], addr_2872_6);

wire[27:0] addr_2873_6;

Selector_2 s2873_6(wires_718_5[1], addr_718_5, addr_positional[11495:11492], addr_2873_6);

wire[27:0] addr_2874_6;

Selector_2 s2874_6(wires_718_5[2], addr_718_5, addr_positional[11499:11496], addr_2874_6);

wire[27:0] addr_2875_6;

Selector_2 s2875_6(wires_718_5[3], addr_718_5, addr_positional[11503:11500], addr_2875_6);

wire[27:0] addr_2876_6;

Selector_2 s2876_6(wires_719_5[0], addr_719_5, addr_positional[11507:11504], addr_2876_6);

wire[27:0] addr_2877_6;

Selector_2 s2877_6(wires_719_5[1], addr_719_5, addr_positional[11511:11508], addr_2877_6);

wire[27:0] addr_2878_6;

Selector_2 s2878_6(wires_719_5[2], addr_719_5, addr_positional[11515:11512], addr_2878_6);

wire[27:0] addr_2879_6;

Selector_2 s2879_6(wires_719_5[3], addr_719_5, addr_positional[11519:11516], addr_2879_6);

wire[27:0] addr_2880_6;

Selector_2 s2880_6(wires_720_5[0], addr_720_5, addr_positional[11523:11520], addr_2880_6);

wire[27:0] addr_2881_6;

Selector_2 s2881_6(wires_720_5[1], addr_720_5, addr_positional[11527:11524], addr_2881_6);

wire[27:0] addr_2882_6;

Selector_2 s2882_6(wires_720_5[2], addr_720_5, addr_positional[11531:11528], addr_2882_6);

wire[27:0] addr_2883_6;

Selector_2 s2883_6(wires_720_5[3], addr_720_5, addr_positional[11535:11532], addr_2883_6);

wire[27:0] addr_2884_6;

Selector_2 s2884_6(wires_721_5[0], addr_721_5, addr_positional[11539:11536], addr_2884_6);

wire[27:0] addr_2885_6;

Selector_2 s2885_6(wires_721_5[1], addr_721_5, addr_positional[11543:11540], addr_2885_6);

wire[27:0] addr_2886_6;

Selector_2 s2886_6(wires_721_5[2], addr_721_5, addr_positional[11547:11544], addr_2886_6);

wire[27:0] addr_2887_6;

Selector_2 s2887_6(wires_721_5[3], addr_721_5, addr_positional[11551:11548], addr_2887_6);

wire[27:0] addr_2888_6;

Selector_2 s2888_6(wires_722_5[0], addr_722_5, addr_positional[11555:11552], addr_2888_6);

wire[27:0] addr_2889_6;

Selector_2 s2889_6(wires_722_5[1], addr_722_5, addr_positional[11559:11556], addr_2889_6);

wire[27:0] addr_2890_6;

Selector_2 s2890_6(wires_722_5[2], addr_722_5, addr_positional[11563:11560], addr_2890_6);

wire[27:0] addr_2891_6;

Selector_2 s2891_6(wires_722_5[3], addr_722_5, addr_positional[11567:11564], addr_2891_6);

wire[27:0] addr_2892_6;

Selector_2 s2892_6(wires_723_5[0], addr_723_5, addr_positional[11571:11568], addr_2892_6);

wire[27:0] addr_2893_6;

Selector_2 s2893_6(wires_723_5[1], addr_723_5, addr_positional[11575:11572], addr_2893_6);

wire[27:0] addr_2894_6;

Selector_2 s2894_6(wires_723_5[2], addr_723_5, addr_positional[11579:11576], addr_2894_6);

wire[27:0] addr_2895_6;

Selector_2 s2895_6(wires_723_5[3], addr_723_5, addr_positional[11583:11580], addr_2895_6);

wire[27:0] addr_2896_6;

Selector_2 s2896_6(wires_724_5[0], addr_724_5, addr_positional[11587:11584], addr_2896_6);

wire[27:0] addr_2897_6;

Selector_2 s2897_6(wires_724_5[1], addr_724_5, addr_positional[11591:11588], addr_2897_6);

wire[27:0] addr_2898_6;

Selector_2 s2898_6(wires_724_5[2], addr_724_5, addr_positional[11595:11592], addr_2898_6);

wire[27:0] addr_2899_6;

Selector_2 s2899_6(wires_724_5[3], addr_724_5, addr_positional[11599:11596], addr_2899_6);

wire[27:0] addr_2900_6;

Selector_2 s2900_6(wires_725_5[0], addr_725_5, addr_positional[11603:11600], addr_2900_6);

wire[27:0] addr_2901_6;

Selector_2 s2901_6(wires_725_5[1], addr_725_5, addr_positional[11607:11604], addr_2901_6);

wire[27:0] addr_2902_6;

Selector_2 s2902_6(wires_725_5[2], addr_725_5, addr_positional[11611:11608], addr_2902_6);

wire[27:0] addr_2903_6;

Selector_2 s2903_6(wires_725_5[3], addr_725_5, addr_positional[11615:11612], addr_2903_6);

wire[27:0] addr_2904_6;

Selector_2 s2904_6(wires_726_5[0], addr_726_5, addr_positional[11619:11616], addr_2904_6);

wire[27:0] addr_2905_6;

Selector_2 s2905_6(wires_726_5[1], addr_726_5, addr_positional[11623:11620], addr_2905_6);

wire[27:0] addr_2906_6;

Selector_2 s2906_6(wires_726_5[2], addr_726_5, addr_positional[11627:11624], addr_2906_6);

wire[27:0] addr_2907_6;

Selector_2 s2907_6(wires_726_5[3], addr_726_5, addr_positional[11631:11628], addr_2907_6);

wire[27:0] addr_2908_6;

Selector_2 s2908_6(wires_727_5[0], addr_727_5, addr_positional[11635:11632], addr_2908_6);

wire[27:0] addr_2909_6;

Selector_2 s2909_6(wires_727_5[1], addr_727_5, addr_positional[11639:11636], addr_2909_6);

wire[27:0] addr_2910_6;

Selector_2 s2910_6(wires_727_5[2], addr_727_5, addr_positional[11643:11640], addr_2910_6);

wire[27:0] addr_2911_6;

Selector_2 s2911_6(wires_727_5[3], addr_727_5, addr_positional[11647:11644], addr_2911_6);

wire[27:0] addr_2912_6;

Selector_2 s2912_6(wires_728_5[0], addr_728_5, addr_positional[11651:11648], addr_2912_6);

wire[27:0] addr_2913_6;

Selector_2 s2913_6(wires_728_5[1], addr_728_5, addr_positional[11655:11652], addr_2913_6);

wire[27:0] addr_2914_6;

Selector_2 s2914_6(wires_728_5[2], addr_728_5, addr_positional[11659:11656], addr_2914_6);

wire[27:0] addr_2915_6;

Selector_2 s2915_6(wires_728_5[3], addr_728_5, addr_positional[11663:11660], addr_2915_6);

wire[27:0] addr_2916_6;

Selector_2 s2916_6(wires_729_5[0], addr_729_5, addr_positional[11667:11664], addr_2916_6);

wire[27:0] addr_2917_6;

Selector_2 s2917_6(wires_729_5[1], addr_729_5, addr_positional[11671:11668], addr_2917_6);

wire[27:0] addr_2918_6;

Selector_2 s2918_6(wires_729_5[2], addr_729_5, addr_positional[11675:11672], addr_2918_6);

wire[27:0] addr_2919_6;

Selector_2 s2919_6(wires_729_5[3], addr_729_5, addr_positional[11679:11676], addr_2919_6);

wire[27:0] addr_2920_6;

Selector_2 s2920_6(wires_730_5[0], addr_730_5, addr_positional[11683:11680], addr_2920_6);

wire[27:0] addr_2921_6;

Selector_2 s2921_6(wires_730_5[1], addr_730_5, addr_positional[11687:11684], addr_2921_6);

wire[27:0] addr_2922_6;

Selector_2 s2922_6(wires_730_5[2], addr_730_5, addr_positional[11691:11688], addr_2922_6);

wire[27:0] addr_2923_6;

Selector_2 s2923_6(wires_730_5[3], addr_730_5, addr_positional[11695:11692], addr_2923_6);

wire[27:0] addr_2924_6;

Selector_2 s2924_6(wires_731_5[0], addr_731_5, addr_positional[11699:11696], addr_2924_6);

wire[27:0] addr_2925_6;

Selector_2 s2925_6(wires_731_5[1], addr_731_5, addr_positional[11703:11700], addr_2925_6);

wire[27:0] addr_2926_6;

Selector_2 s2926_6(wires_731_5[2], addr_731_5, addr_positional[11707:11704], addr_2926_6);

wire[27:0] addr_2927_6;

Selector_2 s2927_6(wires_731_5[3], addr_731_5, addr_positional[11711:11708], addr_2927_6);

wire[27:0] addr_2928_6;

Selector_2 s2928_6(wires_732_5[0], addr_732_5, addr_positional[11715:11712], addr_2928_6);

wire[27:0] addr_2929_6;

Selector_2 s2929_6(wires_732_5[1], addr_732_5, addr_positional[11719:11716], addr_2929_6);

wire[27:0] addr_2930_6;

Selector_2 s2930_6(wires_732_5[2], addr_732_5, addr_positional[11723:11720], addr_2930_6);

wire[27:0] addr_2931_6;

Selector_2 s2931_6(wires_732_5[3], addr_732_5, addr_positional[11727:11724], addr_2931_6);

wire[27:0] addr_2932_6;

Selector_2 s2932_6(wires_733_5[0], addr_733_5, addr_positional[11731:11728], addr_2932_6);

wire[27:0] addr_2933_6;

Selector_2 s2933_6(wires_733_5[1], addr_733_5, addr_positional[11735:11732], addr_2933_6);

wire[27:0] addr_2934_6;

Selector_2 s2934_6(wires_733_5[2], addr_733_5, addr_positional[11739:11736], addr_2934_6);

wire[27:0] addr_2935_6;

Selector_2 s2935_6(wires_733_5[3], addr_733_5, addr_positional[11743:11740], addr_2935_6);

wire[27:0] addr_2936_6;

Selector_2 s2936_6(wires_734_5[0], addr_734_5, addr_positional[11747:11744], addr_2936_6);

wire[27:0] addr_2937_6;

Selector_2 s2937_6(wires_734_5[1], addr_734_5, addr_positional[11751:11748], addr_2937_6);

wire[27:0] addr_2938_6;

Selector_2 s2938_6(wires_734_5[2], addr_734_5, addr_positional[11755:11752], addr_2938_6);

wire[27:0] addr_2939_6;

Selector_2 s2939_6(wires_734_5[3], addr_734_5, addr_positional[11759:11756], addr_2939_6);

wire[27:0] addr_2940_6;

Selector_2 s2940_6(wires_735_5[0], addr_735_5, addr_positional[11763:11760], addr_2940_6);

wire[27:0] addr_2941_6;

Selector_2 s2941_6(wires_735_5[1], addr_735_5, addr_positional[11767:11764], addr_2941_6);

wire[27:0] addr_2942_6;

Selector_2 s2942_6(wires_735_5[2], addr_735_5, addr_positional[11771:11768], addr_2942_6);

wire[27:0] addr_2943_6;

Selector_2 s2943_6(wires_735_5[3], addr_735_5, addr_positional[11775:11772], addr_2943_6);

wire[27:0] addr_2944_6;

Selector_2 s2944_6(wires_736_5[0], addr_736_5, addr_positional[11779:11776], addr_2944_6);

wire[27:0] addr_2945_6;

Selector_2 s2945_6(wires_736_5[1], addr_736_5, addr_positional[11783:11780], addr_2945_6);

wire[27:0] addr_2946_6;

Selector_2 s2946_6(wires_736_5[2], addr_736_5, addr_positional[11787:11784], addr_2946_6);

wire[27:0] addr_2947_6;

Selector_2 s2947_6(wires_736_5[3], addr_736_5, addr_positional[11791:11788], addr_2947_6);

wire[27:0] addr_2948_6;

Selector_2 s2948_6(wires_737_5[0], addr_737_5, addr_positional[11795:11792], addr_2948_6);

wire[27:0] addr_2949_6;

Selector_2 s2949_6(wires_737_5[1], addr_737_5, addr_positional[11799:11796], addr_2949_6);

wire[27:0] addr_2950_6;

Selector_2 s2950_6(wires_737_5[2], addr_737_5, addr_positional[11803:11800], addr_2950_6);

wire[27:0] addr_2951_6;

Selector_2 s2951_6(wires_737_5[3], addr_737_5, addr_positional[11807:11804], addr_2951_6);

wire[27:0] addr_2952_6;

Selector_2 s2952_6(wires_738_5[0], addr_738_5, addr_positional[11811:11808], addr_2952_6);

wire[27:0] addr_2953_6;

Selector_2 s2953_6(wires_738_5[1], addr_738_5, addr_positional[11815:11812], addr_2953_6);

wire[27:0] addr_2954_6;

Selector_2 s2954_6(wires_738_5[2], addr_738_5, addr_positional[11819:11816], addr_2954_6);

wire[27:0] addr_2955_6;

Selector_2 s2955_6(wires_738_5[3], addr_738_5, addr_positional[11823:11820], addr_2955_6);

wire[27:0] addr_2956_6;

Selector_2 s2956_6(wires_739_5[0], addr_739_5, addr_positional[11827:11824], addr_2956_6);

wire[27:0] addr_2957_6;

Selector_2 s2957_6(wires_739_5[1], addr_739_5, addr_positional[11831:11828], addr_2957_6);

wire[27:0] addr_2958_6;

Selector_2 s2958_6(wires_739_5[2], addr_739_5, addr_positional[11835:11832], addr_2958_6);

wire[27:0] addr_2959_6;

Selector_2 s2959_6(wires_739_5[3], addr_739_5, addr_positional[11839:11836], addr_2959_6);

wire[27:0] addr_2960_6;

Selector_2 s2960_6(wires_740_5[0], addr_740_5, addr_positional[11843:11840], addr_2960_6);

wire[27:0] addr_2961_6;

Selector_2 s2961_6(wires_740_5[1], addr_740_5, addr_positional[11847:11844], addr_2961_6);

wire[27:0] addr_2962_6;

Selector_2 s2962_6(wires_740_5[2], addr_740_5, addr_positional[11851:11848], addr_2962_6);

wire[27:0] addr_2963_6;

Selector_2 s2963_6(wires_740_5[3], addr_740_5, addr_positional[11855:11852], addr_2963_6);

wire[27:0] addr_2964_6;

Selector_2 s2964_6(wires_741_5[0], addr_741_5, addr_positional[11859:11856], addr_2964_6);

wire[27:0] addr_2965_6;

Selector_2 s2965_6(wires_741_5[1], addr_741_5, addr_positional[11863:11860], addr_2965_6);

wire[27:0] addr_2966_6;

Selector_2 s2966_6(wires_741_5[2], addr_741_5, addr_positional[11867:11864], addr_2966_6);

wire[27:0] addr_2967_6;

Selector_2 s2967_6(wires_741_5[3], addr_741_5, addr_positional[11871:11868], addr_2967_6);

wire[27:0] addr_2968_6;

Selector_2 s2968_6(wires_742_5[0], addr_742_5, addr_positional[11875:11872], addr_2968_6);

wire[27:0] addr_2969_6;

Selector_2 s2969_6(wires_742_5[1], addr_742_5, addr_positional[11879:11876], addr_2969_6);

wire[27:0] addr_2970_6;

Selector_2 s2970_6(wires_742_5[2], addr_742_5, addr_positional[11883:11880], addr_2970_6);

wire[27:0] addr_2971_6;

Selector_2 s2971_6(wires_742_5[3], addr_742_5, addr_positional[11887:11884], addr_2971_6);

wire[27:0] addr_2972_6;

Selector_2 s2972_6(wires_743_5[0], addr_743_5, addr_positional[11891:11888], addr_2972_6);

wire[27:0] addr_2973_6;

Selector_2 s2973_6(wires_743_5[1], addr_743_5, addr_positional[11895:11892], addr_2973_6);

wire[27:0] addr_2974_6;

Selector_2 s2974_6(wires_743_5[2], addr_743_5, addr_positional[11899:11896], addr_2974_6);

wire[27:0] addr_2975_6;

Selector_2 s2975_6(wires_743_5[3], addr_743_5, addr_positional[11903:11900], addr_2975_6);

wire[27:0] addr_2976_6;

Selector_2 s2976_6(wires_744_5[0], addr_744_5, addr_positional[11907:11904], addr_2976_6);

wire[27:0] addr_2977_6;

Selector_2 s2977_6(wires_744_5[1], addr_744_5, addr_positional[11911:11908], addr_2977_6);

wire[27:0] addr_2978_6;

Selector_2 s2978_6(wires_744_5[2], addr_744_5, addr_positional[11915:11912], addr_2978_6);

wire[27:0] addr_2979_6;

Selector_2 s2979_6(wires_744_5[3], addr_744_5, addr_positional[11919:11916], addr_2979_6);

wire[27:0] addr_2980_6;

Selector_2 s2980_6(wires_745_5[0], addr_745_5, addr_positional[11923:11920], addr_2980_6);

wire[27:0] addr_2981_6;

Selector_2 s2981_6(wires_745_5[1], addr_745_5, addr_positional[11927:11924], addr_2981_6);

wire[27:0] addr_2982_6;

Selector_2 s2982_6(wires_745_5[2], addr_745_5, addr_positional[11931:11928], addr_2982_6);

wire[27:0] addr_2983_6;

Selector_2 s2983_6(wires_745_5[3], addr_745_5, addr_positional[11935:11932], addr_2983_6);

wire[27:0] addr_2984_6;

Selector_2 s2984_6(wires_746_5[0], addr_746_5, addr_positional[11939:11936], addr_2984_6);

wire[27:0] addr_2985_6;

Selector_2 s2985_6(wires_746_5[1], addr_746_5, addr_positional[11943:11940], addr_2985_6);

wire[27:0] addr_2986_6;

Selector_2 s2986_6(wires_746_5[2], addr_746_5, addr_positional[11947:11944], addr_2986_6);

wire[27:0] addr_2987_6;

Selector_2 s2987_6(wires_746_5[3], addr_746_5, addr_positional[11951:11948], addr_2987_6);

wire[27:0] addr_2988_6;

Selector_2 s2988_6(wires_747_5[0], addr_747_5, addr_positional[11955:11952], addr_2988_6);

wire[27:0] addr_2989_6;

Selector_2 s2989_6(wires_747_5[1], addr_747_5, addr_positional[11959:11956], addr_2989_6);

wire[27:0] addr_2990_6;

Selector_2 s2990_6(wires_747_5[2], addr_747_5, addr_positional[11963:11960], addr_2990_6);

wire[27:0] addr_2991_6;

Selector_2 s2991_6(wires_747_5[3], addr_747_5, addr_positional[11967:11964], addr_2991_6);

wire[27:0] addr_2992_6;

Selector_2 s2992_6(wires_748_5[0], addr_748_5, addr_positional[11971:11968], addr_2992_6);

wire[27:0] addr_2993_6;

Selector_2 s2993_6(wires_748_5[1], addr_748_5, addr_positional[11975:11972], addr_2993_6);

wire[27:0] addr_2994_6;

Selector_2 s2994_6(wires_748_5[2], addr_748_5, addr_positional[11979:11976], addr_2994_6);

wire[27:0] addr_2995_6;

Selector_2 s2995_6(wires_748_5[3], addr_748_5, addr_positional[11983:11980], addr_2995_6);

wire[27:0] addr_2996_6;

Selector_2 s2996_6(wires_749_5[0], addr_749_5, addr_positional[11987:11984], addr_2996_6);

wire[27:0] addr_2997_6;

Selector_2 s2997_6(wires_749_5[1], addr_749_5, addr_positional[11991:11988], addr_2997_6);

wire[27:0] addr_2998_6;

Selector_2 s2998_6(wires_749_5[2], addr_749_5, addr_positional[11995:11992], addr_2998_6);

wire[27:0] addr_2999_6;

Selector_2 s2999_6(wires_749_5[3], addr_749_5, addr_positional[11999:11996], addr_2999_6);

wire[27:0] addr_3000_6;

Selector_2 s3000_6(wires_750_5[0], addr_750_5, addr_positional[12003:12000], addr_3000_6);

wire[27:0] addr_3001_6;

Selector_2 s3001_6(wires_750_5[1], addr_750_5, addr_positional[12007:12004], addr_3001_6);

wire[27:0] addr_3002_6;

Selector_2 s3002_6(wires_750_5[2], addr_750_5, addr_positional[12011:12008], addr_3002_6);

wire[27:0] addr_3003_6;

Selector_2 s3003_6(wires_750_5[3], addr_750_5, addr_positional[12015:12012], addr_3003_6);

wire[27:0] addr_3004_6;

Selector_2 s3004_6(wires_751_5[0], addr_751_5, addr_positional[12019:12016], addr_3004_6);

wire[27:0] addr_3005_6;

Selector_2 s3005_6(wires_751_5[1], addr_751_5, addr_positional[12023:12020], addr_3005_6);

wire[27:0] addr_3006_6;

Selector_2 s3006_6(wires_751_5[2], addr_751_5, addr_positional[12027:12024], addr_3006_6);

wire[27:0] addr_3007_6;

Selector_2 s3007_6(wires_751_5[3], addr_751_5, addr_positional[12031:12028], addr_3007_6);

wire[27:0] addr_3008_6;

Selector_2 s3008_6(wires_752_5[0], addr_752_5, addr_positional[12035:12032], addr_3008_6);

wire[27:0] addr_3009_6;

Selector_2 s3009_6(wires_752_5[1], addr_752_5, addr_positional[12039:12036], addr_3009_6);

wire[27:0] addr_3010_6;

Selector_2 s3010_6(wires_752_5[2], addr_752_5, addr_positional[12043:12040], addr_3010_6);

wire[27:0] addr_3011_6;

Selector_2 s3011_6(wires_752_5[3], addr_752_5, addr_positional[12047:12044], addr_3011_6);

wire[27:0] addr_3012_6;

Selector_2 s3012_6(wires_753_5[0], addr_753_5, addr_positional[12051:12048], addr_3012_6);

wire[27:0] addr_3013_6;

Selector_2 s3013_6(wires_753_5[1], addr_753_5, addr_positional[12055:12052], addr_3013_6);

wire[27:0] addr_3014_6;

Selector_2 s3014_6(wires_753_5[2], addr_753_5, addr_positional[12059:12056], addr_3014_6);

wire[27:0] addr_3015_6;

Selector_2 s3015_6(wires_753_5[3], addr_753_5, addr_positional[12063:12060], addr_3015_6);

wire[27:0] addr_3016_6;

Selector_2 s3016_6(wires_754_5[0], addr_754_5, addr_positional[12067:12064], addr_3016_6);

wire[27:0] addr_3017_6;

Selector_2 s3017_6(wires_754_5[1], addr_754_5, addr_positional[12071:12068], addr_3017_6);

wire[27:0] addr_3018_6;

Selector_2 s3018_6(wires_754_5[2], addr_754_5, addr_positional[12075:12072], addr_3018_6);

wire[27:0] addr_3019_6;

Selector_2 s3019_6(wires_754_5[3], addr_754_5, addr_positional[12079:12076], addr_3019_6);

wire[27:0] addr_3020_6;

Selector_2 s3020_6(wires_755_5[0], addr_755_5, addr_positional[12083:12080], addr_3020_6);

wire[27:0] addr_3021_6;

Selector_2 s3021_6(wires_755_5[1], addr_755_5, addr_positional[12087:12084], addr_3021_6);

wire[27:0] addr_3022_6;

Selector_2 s3022_6(wires_755_5[2], addr_755_5, addr_positional[12091:12088], addr_3022_6);

wire[27:0] addr_3023_6;

Selector_2 s3023_6(wires_755_5[3], addr_755_5, addr_positional[12095:12092], addr_3023_6);

wire[27:0] addr_3024_6;

Selector_2 s3024_6(wires_756_5[0], addr_756_5, addr_positional[12099:12096], addr_3024_6);

wire[27:0] addr_3025_6;

Selector_2 s3025_6(wires_756_5[1], addr_756_5, addr_positional[12103:12100], addr_3025_6);

wire[27:0] addr_3026_6;

Selector_2 s3026_6(wires_756_5[2], addr_756_5, addr_positional[12107:12104], addr_3026_6);

wire[27:0] addr_3027_6;

Selector_2 s3027_6(wires_756_5[3], addr_756_5, addr_positional[12111:12108], addr_3027_6);

wire[27:0] addr_3028_6;

Selector_2 s3028_6(wires_757_5[0], addr_757_5, addr_positional[12115:12112], addr_3028_6);

wire[27:0] addr_3029_6;

Selector_2 s3029_6(wires_757_5[1], addr_757_5, addr_positional[12119:12116], addr_3029_6);

wire[27:0] addr_3030_6;

Selector_2 s3030_6(wires_757_5[2], addr_757_5, addr_positional[12123:12120], addr_3030_6);

wire[27:0] addr_3031_6;

Selector_2 s3031_6(wires_757_5[3], addr_757_5, addr_positional[12127:12124], addr_3031_6);

wire[27:0] addr_3032_6;

Selector_2 s3032_6(wires_758_5[0], addr_758_5, addr_positional[12131:12128], addr_3032_6);

wire[27:0] addr_3033_6;

Selector_2 s3033_6(wires_758_5[1], addr_758_5, addr_positional[12135:12132], addr_3033_6);

wire[27:0] addr_3034_6;

Selector_2 s3034_6(wires_758_5[2], addr_758_5, addr_positional[12139:12136], addr_3034_6);

wire[27:0] addr_3035_6;

Selector_2 s3035_6(wires_758_5[3], addr_758_5, addr_positional[12143:12140], addr_3035_6);

wire[27:0] addr_3036_6;

Selector_2 s3036_6(wires_759_5[0], addr_759_5, addr_positional[12147:12144], addr_3036_6);

wire[27:0] addr_3037_6;

Selector_2 s3037_6(wires_759_5[1], addr_759_5, addr_positional[12151:12148], addr_3037_6);

wire[27:0] addr_3038_6;

Selector_2 s3038_6(wires_759_5[2], addr_759_5, addr_positional[12155:12152], addr_3038_6);

wire[27:0] addr_3039_6;

Selector_2 s3039_6(wires_759_5[3], addr_759_5, addr_positional[12159:12156], addr_3039_6);

wire[27:0] addr_3040_6;

Selector_2 s3040_6(wires_760_5[0], addr_760_5, addr_positional[12163:12160], addr_3040_6);

wire[27:0] addr_3041_6;

Selector_2 s3041_6(wires_760_5[1], addr_760_5, addr_positional[12167:12164], addr_3041_6);

wire[27:0] addr_3042_6;

Selector_2 s3042_6(wires_760_5[2], addr_760_5, addr_positional[12171:12168], addr_3042_6);

wire[27:0] addr_3043_6;

Selector_2 s3043_6(wires_760_5[3], addr_760_5, addr_positional[12175:12172], addr_3043_6);

wire[27:0] addr_3044_6;

Selector_2 s3044_6(wires_761_5[0], addr_761_5, addr_positional[12179:12176], addr_3044_6);

wire[27:0] addr_3045_6;

Selector_2 s3045_6(wires_761_5[1], addr_761_5, addr_positional[12183:12180], addr_3045_6);

wire[27:0] addr_3046_6;

Selector_2 s3046_6(wires_761_5[2], addr_761_5, addr_positional[12187:12184], addr_3046_6);

wire[27:0] addr_3047_6;

Selector_2 s3047_6(wires_761_5[3], addr_761_5, addr_positional[12191:12188], addr_3047_6);

wire[27:0] addr_3048_6;

Selector_2 s3048_6(wires_762_5[0], addr_762_5, addr_positional[12195:12192], addr_3048_6);

wire[27:0] addr_3049_6;

Selector_2 s3049_6(wires_762_5[1], addr_762_5, addr_positional[12199:12196], addr_3049_6);

wire[27:0] addr_3050_6;

Selector_2 s3050_6(wires_762_5[2], addr_762_5, addr_positional[12203:12200], addr_3050_6);

wire[27:0] addr_3051_6;

Selector_2 s3051_6(wires_762_5[3], addr_762_5, addr_positional[12207:12204], addr_3051_6);

wire[27:0] addr_3052_6;

Selector_2 s3052_6(wires_763_5[0], addr_763_5, addr_positional[12211:12208], addr_3052_6);

wire[27:0] addr_3053_6;

Selector_2 s3053_6(wires_763_5[1], addr_763_5, addr_positional[12215:12212], addr_3053_6);

wire[27:0] addr_3054_6;

Selector_2 s3054_6(wires_763_5[2], addr_763_5, addr_positional[12219:12216], addr_3054_6);

wire[27:0] addr_3055_6;

Selector_2 s3055_6(wires_763_5[3], addr_763_5, addr_positional[12223:12220], addr_3055_6);

wire[27:0] addr_3056_6;

Selector_2 s3056_6(wires_764_5[0], addr_764_5, addr_positional[12227:12224], addr_3056_6);

wire[27:0] addr_3057_6;

Selector_2 s3057_6(wires_764_5[1], addr_764_5, addr_positional[12231:12228], addr_3057_6);

wire[27:0] addr_3058_6;

Selector_2 s3058_6(wires_764_5[2], addr_764_5, addr_positional[12235:12232], addr_3058_6);

wire[27:0] addr_3059_6;

Selector_2 s3059_6(wires_764_5[3], addr_764_5, addr_positional[12239:12236], addr_3059_6);

wire[27:0] addr_3060_6;

Selector_2 s3060_6(wires_765_5[0], addr_765_5, addr_positional[12243:12240], addr_3060_6);

wire[27:0] addr_3061_6;

Selector_2 s3061_6(wires_765_5[1], addr_765_5, addr_positional[12247:12244], addr_3061_6);

wire[27:0] addr_3062_6;

Selector_2 s3062_6(wires_765_5[2], addr_765_5, addr_positional[12251:12248], addr_3062_6);

wire[27:0] addr_3063_6;

Selector_2 s3063_6(wires_765_5[3], addr_765_5, addr_positional[12255:12252], addr_3063_6);

wire[27:0] addr_3064_6;

Selector_2 s3064_6(wires_766_5[0], addr_766_5, addr_positional[12259:12256], addr_3064_6);

wire[27:0] addr_3065_6;

Selector_2 s3065_6(wires_766_5[1], addr_766_5, addr_positional[12263:12260], addr_3065_6);

wire[27:0] addr_3066_6;

Selector_2 s3066_6(wires_766_5[2], addr_766_5, addr_positional[12267:12264], addr_3066_6);

wire[27:0] addr_3067_6;

Selector_2 s3067_6(wires_766_5[3], addr_766_5, addr_positional[12271:12268], addr_3067_6);

wire[27:0] addr_3068_6;

Selector_2 s3068_6(wires_767_5[0], addr_767_5, addr_positional[12275:12272], addr_3068_6);

wire[27:0] addr_3069_6;

Selector_2 s3069_6(wires_767_5[1], addr_767_5, addr_positional[12279:12276], addr_3069_6);

wire[27:0] addr_3070_6;

Selector_2 s3070_6(wires_767_5[2], addr_767_5, addr_positional[12283:12280], addr_3070_6);

wire[27:0] addr_3071_6;

Selector_2 s3071_6(wires_767_5[3], addr_767_5, addr_positional[12287:12284], addr_3071_6);

wire[27:0] addr_3072_6;

Selector_2 s3072_6(wires_768_5[0], addr_768_5, addr_positional[12291:12288], addr_3072_6);

wire[27:0] addr_3073_6;

Selector_2 s3073_6(wires_768_5[1], addr_768_5, addr_positional[12295:12292], addr_3073_6);

wire[27:0] addr_3074_6;

Selector_2 s3074_6(wires_768_5[2], addr_768_5, addr_positional[12299:12296], addr_3074_6);

wire[27:0] addr_3075_6;

Selector_2 s3075_6(wires_768_5[3], addr_768_5, addr_positional[12303:12300], addr_3075_6);

wire[27:0] addr_3076_6;

Selector_2 s3076_6(wires_769_5[0], addr_769_5, addr_positional[12307:12304], addr_3076_6);

wire[27:0] addr_3077_6;

Selector_2 s3077_6(wires_769_5[1], addr_769_5, addr_positional[12311:12308], addr_3077_6);

wire[27:0] addr_3078_6;

Selector_2 s3078_6(wires_769_5[2], addr_769_5, addr_positional[12315:12312], addr_3078_6);

wire[27:0] addr_3079_6;

Selector_2 s3079_6(wires_769_5[3], addr_769_5, addr_positional[12319:12316], addr_3079_6);

wire[27:0] addr_3080_6;

Selector_2 s3080_6(wires_770_5[0], addr_770_5, addr_positional[12323:12320], addr_3080_6);

wire[27:0] addr_3081_6;

Selector_2 s3081_6(wires_770_5[1], addr_770_5, addr_positional[12327:12324], addr_3081_6);

wire[27:0] addr_3082_6;

Selector_2 s3082_6(wires_770_5[2], addr_770_5, addr_positional[12331:12328], addr_3082_6);

wire[27:0] addr_3083_6;

Selector_2 s3083_6(wires_770_5[3], addr_770_5, addr_positional[12335:12332], addr_3083_6);

wire[27:0] addr_3084_6;

Selector_2 s3084_6(wires_771_5[0], addr_771_5, addr_positional[12339:12336], addr_3084_6);

wire[27:0] addr_3085_6;

Selector_2 s3085_6(wires_771_5[1], addr_771_5, addr_positional[12343:12340], addr_3085_6);

wire[27:0] addr_3086_6;

Selector_2 s3086_6(wires_771_5[2], addr_771_5, addr_positional[12347:12344], addr_3086_6);

wire[27:0] addr_3087_6;

Selector_2 s3087_6(wires_771_5[3], addr_771_5, addr_positional[12351:12348], addr_3087_6);

wire[27:0] addr_3088_6;

Selector_2 s3088_6(wires_772_5[0], addr_772_5, addr_positional[12355:12352], addr_3088_6);

wire[27:0] addr_3089_6;

Selector_2 s3089_6(wires_772_5[1], addr_772_5, addr_positional[12359:12356], addr_3089_6);

wire[27:0] addr_3090_6;

Selector_2 s3090_6(wires_772_5[2], addr_772_5, addr_positional[12363:12360], addr_3090_6);

wire[27:0] addr_3091_6;

Selector_2 s3091_6(wires_772_5[3], addr_772_5, addr_positional[12367:12364], addr_3091_6);

wire[27:0] addr_3092_6;

Selector_2 s3092_6(wires_773_5[0], addr_773_5, addr_positional[12371:12368], addr_3092_6);

wire[27:0] addr_3093_6;

Selector_2 s3093_6(wires_773_5[1], addr_773_5, addr_positional[12375:12372], addr_3093_6);

wire[27:0] addr_3094_6;

Selector_2 s3094_6(wires_773_5[2], addr_773_5, addr_positional[12379:12376], addr_3094_6);

wire[27:0] addr_3095_6;

Selector_2 s3095_6(wires_773_5[3], addr_773_5, addr_positional[12383:12380], addr_3095_6);

wire[27:0] addr_3096_6;

Selector_2 s3096_6(wires_774_5[0], addr_774_5, addr_positional[12387:12384], addr_3096_6);

wire[27:0] addr_3097_6;

Selector_2 s3097_6(wires_774_5[1], addr_774_5, addr_positional[12391:12388], addr_3097_6);

wire[27:0] addr_3098_6;

Selector_2 s3098_6(wires_774_5[2], addr_774_5, addr_positional[12395:12392], addr_3098_6);

wire[27:0] addr_3099_6;

Selector_2 s3099_6(wires_774_5[3], addr_774_5, addr_positional[12399:12396], addr_3099_6);

wire[27:0] addr_3100_6;

Selector_2 s3100_6(wires_775_5[0], addr_775_5, addr_positional[12403:12400], addr_3100_6);

wire[27:0] addr_3101_6;

Selector_2 s3101_6(wires_775_5[1], addr_775_5, addr_positional[12407:12404], addr_3101_6);

wire[27:0] addr_3102_6;

Selector_2 s3102_6(wires_775_5[2], addr_775_5, addr_positional[12411:12408], addr_3102_6);

wire[27:0] addr_3103_6;

Selector_2 s3103_6(wires_775_5[3], addr_775_5, addr_positional[12415:12412], addr_3103_6);

wire[27:0] addr_3104_6;

Selector_2 s3104_6(wires_776_5[0], addr_776_5, addr_positional[12419:12416], addr_3104_6);

wire[27:0] addr_3105_6;

Selector_2 s3105_6(wires_776_5[1], addr_776_5, addr_positional[12423:12420], addr_3105_6);

wire[27:0] addr_3106_6;

Selector_2 s3106_6(wires_776_5[2], addr_776_5, addr_positional[12427:12424], addr_3106_6);

wire[27:0] addr_3107_6;

Selector_2 s3107_6(wires_776_5[3], addr_776_5, addr_positional[12431:12428], addr_3107_6);

wire[27:0] addr_3108_6;

Selector_2 s3108_6(wires_777_5[0], addr_777_5, addr_positional[12435:12432], addr_3108_6);

wire[27:0] addr_3109_6;

Selector_2 s3109_6(wires_777_5[1], addr_777_5, addr_positional[12439:12436], addr_3109_6);

wire[27:0] addr_3110_6;

Selector_2 s3110_6(wires_777_5[2], addr_777_5, addr_positional[12443:12440], addr_3110_6);

wire[27:0] addr_3111_6;

Selector_2 s3111_6(wires_777_5[3], addr_777_5, addr_positional[12447:12444], addr_3111_6);

wire[27:0] addr_3112_6;

Selector_2 s3112_6(wires_778_5[0], addr_778_5, addr_positional[12451:12448], addr_3112_6);

wire[27:0] addr_3113_6;

Selector_2 s3113_6(wires_778_5[1], addr_778_5, addr_positional[12455:12452], addr_3113_6);

wire[27:0] addr_3114_6;

Selector_2 s3114_6(wires_778_5[2], addr_778_5, addr_positional[12459:12456], addr_3114_6);

wire[27:0] addr_3115_6;

Selector_2 s3115_6(wires_778_5[3], addr_778_5, addr_positional[12463:12460], addr_3115_6);

wire[27:0] addr_3116_6;

Selector_2 s3116_6(wires_779_5[0], addr_779_5, addr_positional[12467:12464], addr_3116_6);

wire[27:0] addr_3117_6;

Selector_2 s3117_6(wires_779_5[1], addr_779_5, addr_positional[12471:12468], addr_3117_6);

wire[27:0] addr_3118_6;

Selector_2 s3118_6(wires_779_5[2], addr_779_5, addr_positional[12475:12472], addr_3118_6);

wire[27:0] addr_3119_6;

Selector_2 s3119_6(wires_779_5[3], addr_779_5, addr_positional[12479:12476], addr_3119_6);

wire[27:0] addr_3120_6;

Selector_2 s3120_6(wires_780_5[0], addr_780_5, addr_positional[12483:12480], addr_3120_6);

wire[27:0] addr_3121_6;

Selector_2 s3121_6(wires_780_5[1], addr_780_5, addr_positional[12487:12484], addr_3121_6);

wire[27:0] addr_3122_6;

Selector_2 s3122_6(wires_780_5[2], addr_780_5, addr_positional[12491:12488], addr_3122_6);

wire[27:0] addr_3123_6;

Selector_2 s3123_6(wires_780_5[3], addr_780_5, addr_positional[12495:12492], addr_3123_6);

wire[27:0] addr_3124_6;

Selector_2 s3124_6(wires_781_5[0], addr_781_5, addr_positional[12499:12496], addr_3124_6);

wire[27:0] addr_3125_6;

Selector_2 s3125_6(wires_781_5[1], addr_781_5, addr_positional[12503:12500], addr_3125_6);

wire[27:0] addr_3126_6;

Selector_2 s3126_6(wires_781_5[2], addr_781_5, addr_positional[12507:12504], addr_3126_6);

wire[27:0] addr_3127_6;

Selector_2 s3127_6(wires_781_5[3], addr_781_5, addr_positional[12511:12508], addr_3127_6);

wire[27:0] addr_3128_6;

Selector_2 s3128_6(wires_782_5[0], addr_782_5, addr_positional[12515:12512], addr_3128_6);

wire[27:0] addr_3129_6;

Selector_2 s3129_6(wires_782_5[1], addr_782_5, addr_positional[12519:12516], addr_3129_6);

wire[27:0] addr_3130_6;

Selector_2 s3130_6(wires_782_5[2], addr_782_5, addr_positional[12523:12520], addr_3130_6);

wire[27:0] addr_3131_6;

Selector_2 s3131_6(wires_782_5[3], addr_782_5, addr_positional[12527:12524], addr_3131_6);

wire[27:0] addr_3132_6;

Selector_2 s3132_6(wires_783_5[0], addr_783_5, addr_positional[12531:12528], addr_3132_6);

wire[27:0] addr_3133_6;

Selector_2 s3133_6(wires_783_5[1], addr_783_5, addr_positional[12535:12532], addr_3133_6);

wire[27:0] addr_3134_6;

Selector_2 s3134_6(wires_783_5[2], addr_783_5, addr_positional[12539:12536], addr_3134_6);

wire[27:0] addr_3135_6;

Selector_2 s3135_6(wires_783_5[3], addr_783_5, addr_positional[12543:12540], addr_3135_6);

wire[27:0] addr_3136_6;

Selector_2 s3136_6(wires_784_5[0], addr_784_5, addr_positional[12547:12544], addr_3136_6);

wire[27:0] addr_3137_6;

Selector_2 s3137_6(wires_784_5[1], addr_784_5, addr_positional[12551:12548], addr_3137_6);

wire[27:0] addr_3138_6;

Selector_2 s3138_6(wires_784_5[2], addr_784_5, addr_positional[12555:12552], addr_3138_6);

wire[27:0] addr_3139_6;

Selector_2 s3139_6(wires_784_5[3], addr_784_5, addr_positional[12559:12556], addr_3139_6);

wire[27:0] addr_3140_6;

Selector_2 s3140_6(wires_785_5[0], addr_785_5, addr_positional[12563:12560], addr_3140_6);

wire[27:0] addr_3141_6;

Selector_2 s3141_6(wires_785_5[1], addr_785_5, addr_positional[12567:12564], addr_3141_6);

wire[27:0] addr_3142_6;

Selector_2 s3142_6(wires_785_5[2], addr_785_5, addr_positional[12571:12568], addr_3142_6);

wire[27:0] addr_3143_6;

Selector_2 s3143_6(wires_785_5[3], addr_785_5, addr_positional[12575:12572], addr_3143_6);

wire[27:0] addr_3144_6;

Selector_2 s3144_6(wires_786_5[0], addr_786_5, addr_positional[12579:12576], addr_3144_6);

wire[27:0] addr_3145_6;

Selector_2 s3145_6(wires_786_5[1], addr_786_5, addr_positional[12583:12580], addr_3145_6);

wire[27:0] addr_3146_6;

Selector_2 s3146_6(wires_786_5[2], addr_786_5, addr_positional[12587:12584], addr_3146_6);

wire[27:0] addr_3147_6;

Selector_2 s3147_6(wires_786_5[3], addr_786_5, addr_positional[12591:12588], addr_3147_6);

wire[27:0] addr_3148_6;

Selector_2 s3148_6(wires_787_5[0], addr_787_5, addr_positional[12595:12592], addr_3148_6);

wire[27:0] addr_3149_6;

Selector_2 s3149_6(wires_787_5[1], addr_787_5, addr_positional[12599:12596], addr_3149_6);

wire[27:0] addr_3150_6;

Selector_2 s3150_6(wires_787_5[2], addr_787_5, addr_positional[12603:12600], addr_3150_6);

wire[27:0] addr_3151_6;

Selector_2 s3151_6(wires_787_5[3], addr_787_5, addr_positional[12607:12604], addr_3151_6);

wire[27:0] addr_3152_6;

Selector_2 s3152_6(wires_788_5[0], addr_788_5, addr_positional[12611:12608], addr_3152_6);

wire[27:0] addr_3153_6;

Selector_2 s3153_6(wires_788_5[1], addr_788_5, addr_positional[12615:12612], addr_3153_6);

wire[27:0] addr_3154_6;

Selector_2 s3154_6(wires_788_5[2], addr_788_5, addr_positional[12619:12616], addr_3154_6);

wire[27:0] addr_3155_6;

Selector_2 s3155_6(wires_788_5[3], addr_788_5, addr_positional[12623:12620], addr_3155_6);

wire[27:0] addr_3156_6;

Selector_2 s3156_6(wires_789_5[0], addr_789_5, addr_positional[12627:12624], addr_3156_6);

wire[27:0] addr_3157_6;

Selector_2 s3157_6(wires_789_5[1], addr_789_5, addr_positional[12631:12628], addr_3157_6);

wire[27:0] addr_3158_6;

Selector_2 s3158_6(wires_789_5[2], addr_789_5, addr_positional[12635:12632], addr_3158_6);

wire[27:0] addr_3159_6;

Selector_2 s3159_6(wires_789_5[3], addr_789_5, addr_positional[12639:12636], addr_3159_6);

wire[27:0] addr_3160_6;

Selector_2 s3160_6(wires_790_5[0], addr_790_5, addr_positional[12643:12640], addr_3160_6);

wire[27:0] addr_3161_6;

Selector_2 s3161_6(wires_790_5[1], addr_790_5, addr_positional[12647:12644], addr_3161_6);

wire[27:0] addr_3162_6;

Selector_2 s3162_6(wires_790_5[2], addr_790_5, addr_positional[12651:12648], addr_3162_6);

wire[27:0] addr_3163_6;

Selector_2 s3163_6(wires_790_5[3], addr_790_5, addr_positional[12655:12652], addr_3163_6);

wire[27:0] addr_3164_6;

Selector_2 s3164_6(wires_791_5[0], addr_791_5, addr_positional[12659:12656], addr_3164_6);

wire[27:0] addr_3165_6;

Selector_2 s3165_6(wires_791_5[1], addr_791_5, addr_positional[12663:12660], addr_3165_6);

wire[27:0] addr_3166_6;

Selector_2 s3166_6(wires_791_5[2], addr_791_5, addr_positional[12667:12664], addr_3166_6);

wire[27:0] addr_3167_6;

Selector_2 s3167_6(wires_791_5[3], addr_791_5, addr_positional[12671:12668], addr_3167_6);

wire[27:0] addr_3168_6;

Selector_2 s3168_6(wires_792_5[0], addr_792_5, addr_positional[12675:12672], addr_3168_6);

wire[27:0] addr_3169_6;

Selector_2 s3169_6(wires_792_5[1], addr_792_5, addr_positional[12679:12676], addr_3169_6);

wire[27:0] addr_3170_6;

Selector_2 s3170_6(wires_792_5[2], addr_792_5, addr_positional[12683:12680], addr_3170_6);

wire[27:0] addr_3171_6;

Selector_2 s3171_6(wires_792_5[3], addr_792_5, addr_positional[12687:12684], addr_3171_6);

wire[27:0] addr_3172_6;

Selector_2 s3172_6(wires_793_5[0], addr_793_5, addr_positional[12691:12688], addr_3172_6);

wire[27:0] addr_3173_6;

Selector_2 s3173_6(wires_793_5[1], addr_793_5, addr_positional[12695:12692], addr_3173_6);

wire[27:0] addr_3174_6;

Selector_2 s3174_6(wires_793_5[2], addr_793_5, addr_positional[12699:12696], addr_3174_6);

wire[27:0] addr_3175_6;

Selector_2 s3175_6(wires_793_5[3], addr_793_5, addr_positional[12703:12700], addr_3175_6);

wire[27:0] addr_3176_6;

Selector_2 s3176_6(wires_794_5[0], addr_794_5, addr_positional[12707:12704], addr_3176_6);

wire[27:0] addr_3177_6;

Selector_2 s3177_6(wires_794_5[1], addr_794_5, addr_positional[12711:12708], addr_3177_6);

wire[27:0] addr_3178_6;

Selector_2 s3178_6(wires_794_5[2], addr_794_5, addr_positional[12715:12712], addr_3178_6);

wire[27:0] addr_3179_6;

Selector_2 s3179_6(wires_794_5[3], addr_794_5, addr_positional[12719:12716], addr_3179_6);

wire[27:0] addr_3180_6;

Selector_2 s3180_6(wires_795_5[0], addr_795_5, addr_positional[12723:12720], addr_3180_6);

wire[27:0] addr_3181_6;

Selector_2 s3181_6(wires_795_5[1], addr_795_5, addr_positional[12727:12724], addr_3181_6);

wire[27:0] addr_3182_6;

Selector_2 s3182_6(wires_795_5[2], addr_795_5, addr_positional[12731:12728], addr_3182_6);

wire[27:0] addr_3183_6;

Selector_2 s3183_6(wires_795_5[3], addr_795_5, addr_positional[12735:12732], addr_3183_6);

wire[27:0] addr_3184_6;

Selector_2 s3184_6(wires_796_5[0], addr_796_5, addr_positional[12739:12736], addr_3184_6);

wire[27:0] addr_3185_6;

Selector_2 s3185_6(wires_796_5[1], addr_796_5, addr_positional[12743:12740], addr_3185_6);

wire[27:0] addr_3186_6;

Selector_2 s3186_6(wires_796_5[2], addr_796_5, addr_positional[12747:12744], addr_3186_6);

wire[27:0] addr_3187_6;

Selector_2 s3187_6(wires_796_5[3], addr_796_5, addr_positional[12751:12748], addr_3187_6);

wire[27:0] addr_3188_6;

Selector_2 s3188_6(wires_797_5[0], addr_797_5, addr_positional[12755:12752], addr_3188_6);

wire[27:0] addr_3189_6;

Selector_2 s3189_6(wires_797_5[1], addr_797_5, addr_positional[12759:12756], addr_3189_6);

wire[27:0] addr_3190_6;

Selector_2 s3190_6(wires_797_5[2], addr_797_5, addr_positional[12763:12760], addr_3190_6);

wire[27:0] addr_3191_6;

Selector_2 s3191_6(wires_797_5[3], addr_797_5, addr_positional[12767:12764], addr_3191_6);

wire[27:0] addr_3192_6;

Selector_2 s3192_6(wires_798_5[0], addr_798_5, addr_positional[12771:12768], addr_3192_6);

wire[27:0] addr_3193_6;

Selector_2 s3193_6(wires_798_5[1], addr_798_5, addr_positional[12775:12772], addr_3193_6);

wire[27:0] addr_3194_6;

Selector_2 s3194_6(wires_798_5[2], addr_798_5, addr_positional[12779:12776], addr_3194_6);

wire[27:0] addr_3195_6;

Selector_2 s3195_6(wires_798_5[3], addr_798_5, addr_positional[12783:12780], addr_3195_6);

wire[27:0] addr_3196_6;

Selector_2 s3196_6(wires_799_5[0], addr_799_5, addr_positional[12787:12784], addr_3196_6);

wire[27:0] addr_3197_6;

Selector_2 s3197_6(wires_799_5[1], addr_799_5, addr_positional[12791:12788], addr_3197_6);

wire[27:0] addr_3198_6;

Selector_2 s3198_6(wires_799_5[2], addr_799_5, addr_positional[12795:12792], addr_3198_6);

wire[27:0] addr_3199_6;

Selector_2 s3199_6(wires_799_5[3], addr_799_5, addr_positional[12799:12796], addr_3199_6);

wire[27:0] addr_3200_6;

Selector_2 s3200_6(wires_800_5[0], addr_800_5, addr_positional[12803:12800], addr_3200_6);

wire[27:0] addr_3201_6;

Selector_2 s3201_6(wires_800_5[1], addr_800_5, addr_positional[12807:12804], addr_3201_6);

wire[27:0] addr_3202_6;

Selector_2 s3202_6(wires_800_5[2], addr_800_5, addr_positional[12811:12808], addr_3202_6);

wire[27:0] addr_3203_6;

Selector_2 s3203_6(wires_800_5[3], addr_800_5, addr_positional[12815:12812], addr_3203_6);

wire[27:0] addr_3204_6;

Selector_2 s3204_6(wires_801_5[0], addr_801_5, addr_positional[12819:12816], addr_3204_6);

wire[27:0] addr_3205_6;

Selector_2 s3205_6(wires_801_5[1], addr_801_5, addr_positional[12823:12820], addr_3205_6);

wire[27:0] addr_3206_6;

Selector_2 s3206_6(wires_801_5[2], addr_801_5, addr_positional[12827:12824], addr_3206_6);

wire[27:0] addr_3207_6;

Selector_2 s3207_6(wires_801_5[3], addr_801_5, addr_positional[12831:12828], addr_3207_6);

wire[27:0] addr_3208_6;

Selector_2 s3208_6(wires_802_5[0], addr_802_5, addr_positional[12835:12832], addr_3208_6);

wire[27:0] addr_3209_6;

Selector_2 s3209_6(wires_802_5[1], addr_802_5, addr_positional[12839:12836], addr_3209_6);

wire[27:0] addr_3210_6;

Selector_2 s3210_6(wires_802_5[2], addr_802_5, addr_positional[12843:12840], addr_3210_6);

wire[27:0] addr_3211_6;

Selector_2 s3211_6(wires_802_5[3], addr_802_5, addr_positional[12847:12844], addr_3211_6);

wire[27:0] addr_3212_6;

Selector_2 s3212_6(wires_803_5[0], addr_803_5, addr_positional[12851:12848], addr_3212_6);

wire[27:0] addr_3213_6;

Selector_2 s3213_6(wires_803_5[1], addr_803_5, addr_positional[12855:12852], addr_3213_6);

wire[27:0] addr_3214_6;

Selector_2 s3214_6(wires_803_5[2], addr_803_5, addr_positional[12859:12856], addr_3214_6);

wire[27:0] addr_3215_6;

Selector_2 s3215_6(wires_803_5[3], addr_803_5, addr_positional[12863:12860], addr_3215_6);

wire[27:0] addr_3216_6;

Selector_2 s3216_6(wires_804_5[0], addr_804_5, addr_positional[12867:12864], addr_3216_6);

wire[27:0] addr_3217_6;

Selector_2 s3217_6(wires_804_5[1], addr_804_5, addr_positional[12871:12868], addr_3217_6);

wire[27:0] addr_3218_6;

Selector_2 s3218_6(wires_804_5[2], addr_804_5, addr_positional[12875:12872], addr_3218_6);

wire[27:0] addr_3219_6;

Selector_2 s3219_6(wires_804_5[3], addr_804_5, addr_positional[12879:12876], addr_3219_6);

wire[27:0] addr_3220_6;

Selector_2 s3220_6(wires_805_5[0], addr_805_5, addr_positional[12883:12880], addr_3220_6);

wire[27:0] addr_3221_6;

Selector_2 s3221_6(wires_805_5[1], addr_805_5, addr_positional[12887:12884], addr_3221_6);

wire[27:0] addr_3222_6;

Selector_2 s3222_6(wires_805_5[2], addr_805_5, addr_positional[12891:12888], addr_3222_6);

wire[27:0] addr_3223_6;

Selector_2 s3223_6(wires_805_5[3], addr_805_5, addr_positional[12895:12892], addr_3223_6);

wire[27:0] addr_3224_6;

Selector_2 s3224_6(wires_806_5[0], addr_806_5, addr_positional[12899:12896], addr_3224_6);

wire[27:0] addr_3225_6;

Selector_2 s3225_6(wires_806_5[1], addr_806_5, addr_positional[12903:12900], addr_3225_6);

wire[27:0] addr_3226_6;

Selector_2 s3226_6(wires_806_5[2], addr_806_5, addr_positional[12907:12904], addr_3226_6);

wire[27:0] addr_3227_6;

Selector_2 s3227_6(wires_806_5[3], addr_806_5, addr_positional[12911:12908], addr_3227_6);

wire[27:0] addr_3228_6;

Selector_2 s3228_6(wires_807_5[0], addr_807_5, addr_positional[12915:12912], addr_3228_6);

wire[27:0] addr_3229_6;

Selector_2 s3229_6(wires_807_5[1], addr_807_5, addr_positional[12919:12916], addr_3229_6);

wire[27:0] addr_3230_6;

Selector_2 s3230_6(wires_807_5[2], addr_807_5, addr_positional[12923:12920], addr_3230_6);

wire[27:0] addr_3231_6;

Selector_2 s3231_6(wires_807_5[3], addr_807_5, addr_positional[12927:12924], addr_3231_6);

wire[27:0] addr_3232_6;

Selector_2 s3232_6(wires_808_5[0], addr_808_5, addr_positional[12931:12928], addr_3232_6);

wire[27:0] addr_3233_6;

Selector_2 s3233_6(wires_808_5[1], addr_808_5, addr_positional[12935:12932], addr_3233_6);

wire[27:0] addr_3234_6;

Selector_2 s3234_6(wires_808_5[2], addr_808_5, addr_positional[12939:12936], addr_3234_6);

wire[27:0] addr_3235_6;

Selector_2 s3235_6(wires_808_5[3], addr_808_5, addr_positional[12943:12940], addr_3235_6);

wire[27:0] addr_3236_6;

Selector_2 s3236_6(wires_809_5[0], addr_809_5, addr_positional[12947:12944], addr_3236_6);

wire[27:0] addr_3237_6;

Selector_2 s3237_6(wires_809_5[1], addr_809_5, addr_positional[12951:12948], addr_3237_6);

wire[27:0] addr_3238_6;

Selector_2 s3238_6(wires_809_5[2], addr_809_5, addr_positional[12955:12952], addr_3238_6);

wire[27:0] addr_3239_6;

Selector_2 s3239_6(wires_809_5[3], addr_809_5, addr_positional[12959:12956], addr_3239_6);

wire[27:0] addr_3240_6;

Selector_2 s3240_6(wires_810_5[0], addr_810_5, addr_positional[12963:12960], addr_3240_6);

wire[27:0] addr_3241_6;

Selector_2 s3241_6(wires_810_5[1], addr_810_5, addr_positional[12967:12964], addr_3241_6);

wire[27:0] addr_3242_6;

Selector_2 s3242_6(wires_810_5[2], addr_810_5, addr_positional[12971:12968], addr_3242_6);

wire[27:0] addr_3243_6;

Selector_2 s3243_6(wires_810_5[3], addr_810_5, addr_positional[12975:12972], addr_3243_6);

wire[27:0] addr_3244_6;

Selector_2 s3244_6(wires_811_5[0], addr_811_5, addr_positional[12979:12976], addr_3244_6);

wire[27:0] addr_3245_6;

Selector_2 s3245_6(wires_811_5[1], addr_811_5, addr_positional[12983:12980], addr_3245_6);

wire[27:0] addr_3246_6;

Selector_2 s3246_6(wires_811_5[2], addr_811_5, addr_positional[12987:12984], addr_3246_6);

wire[27:0] addr_3247_6;

Selector_2 s3247_6(wires_811_5[3], addr_811_5, addr_positional[12991:12988], addr_3247_6);

wire[27:0] addr_3248_6;

Selector_2 s3248_6(wires_812_5[0], addr_812_5, addr_positional[12995:12992], addr_3248_6);

wire[27:0] addr_3249_6;

Selector_2 s3249_6(wires_812_5[1], addr_812_5, addr_positional[12999:12996], addr_3249_6);

wire[27:0] addr_3250_6;

Selector_2 s3250_6(wires_812_5[2], addr_812_5, addr_positional[13003:13000], addr_3250_6);

wire[27:0] addr_3251_6;

Selector_2 s3251_6(wires_812_5[3], addr_812_5, addr_positional[13007:13004], addr_3251_6);

wire[27:0] addr_3252_6;

Selector_2 s3252_6(wires_813_5[0], addr_813_5, addr_positional[13011:13008], addr_3252_6);

wire[27:0] addr_3253_6;

Selector_2 s3253_6(wires_813_5[1], addr_813_5, addr_positional[13015:13012], addr_3253_6);

wire[27:0] addr_3254_6;

Selector_2 s3254_6(wires_813_5[2], addr_813_5, addr_positional[13019:13016], addr_3254_6);

wire[27:0] addr_3255_6;

Selector_2 s3255_6(wires_813_5[3], addr_813_5, addr_positional[13023:13020], addr_3255_6);

wire[27:0] addr_3256_6;

Selector_2 s3256_6(wires_814_5[0], addr_814_5, addr_positional[13027:13024], addr_3256_6);

wire[27:0] addr_3257_6;

Selector_2 s3257_6(wires_814_5[1], addr_814_5, addr_positional[13031:13028], addr_3257_6);

wire[27:0] addr_3258_6;

Selector_2 s3258_6(wires_814_5[2], addr_814_5, addr_positional[13035:13032], addr_3258_6);

wire[27:0] addr_3259_6;

Selector_2 s3259_6(wires_814_5[3], addr_814_5, addr_positional[13039:13036], addr_3259_6);

wire[27:0] addr_3260_6;

Selector_2 s3260_6(wires_815_5[0], addr_815_5, addr_positional[13043:13040], addr_3260_6);

wire[27:0] addr_3261_6;

Selector_2 s3261_6(wires_815_5[1], addr_815_5, addr_positional[13047:13044], addr_3261_6);

wire[27:0] addr_3262_6;

Selector_2 s3262_6(wires_815_5[2], addr_815_5, addr_positional[13051:13048], addr_3262_6);

wire[27:0] addr_3263_6;

Selector_2 s3263_6(wires_815_5[3], addr_815_5, addr_positional[13055:13052], addr_3263_6);

wire[27:0] addr_3264_6;

Selector_2 s3264_6(wires_816_5[0], addr_816_5, addr_positional[13059:13056], addr_3264_6);

wire[27:0] addr_3265_6;

Selector_2 s3265_6(wires_816_5[1], addr_816_5, addr_positional[13063:13060], addr_3265_6);

wire[27:0] addr_3266_6;

Selector_2 s3266_6(wires_816_5[2], addr_816_5, addr_positional[13067:13064], addr_3266_6);

wire[27:0] addr_3267_6;

Selector_2 s3267_6(wires_816_5[3], addr_816_5, addr_positional[13071:13068], addr_3267_6);

wire[27:0] addr_3268_6;

Selector_2 s3268_6(wires_817_5[0], addr_817_5, addr_positional[13075:13072], addr_3268_6);

wire[27:0] addr_3269_6;

Selector_2 s3269_6(wires_817_5[1], addr_817_5, addr_positional[13079:13076], addr_3269_6);

wire[27:0] addr_3270_6;

Selector_2 s3270_6(wires_817_5[2], addr_817_5, addr_positional[13083:13080], addr_3270_6);

wire[27:0] addr_3271_6;

Selector_2 s3271_6(wires_817_5[3], addr_817_5, addr_positional[13087:13084], addr_3271_6);

wire[27:0] addr_3272_6;

Selector_2 s3272_6(wires_818_5[0], addr_818_5, addr_positional[13091:13088], addr_3272_6);

wire[27:0] addr_3273_6;

Selector_2 s3273_6(wires_818_5[1], addr_818_5, addr_positional[13095:13092], addr_3273_6);

wire[27:0] addr_3274_6;

Selector_2 s3274_6(wires_818_5[2], addr_818_5, addr_positional[13099:13096], addr_3274_6);

wire[27:0] addr_3275_6;

Selector_2 s3275_6(wires_818_5[3], addr_818_5, addr_positional[13103:13100], addr_3275_6);

wire[27:0] addr_3276_6;

Selector_2 s3276_6(wires_819_5[0], addr_819_5, addr_positional[13107:13104], addr_3276_6);

wire[27:0] addr_3277_6;

Selector_2 s3277_6(wires_819_5[1], addr_819_5, addr_positional[13111:13108], addr_3277_6);

wire[27:0] addr_3278_6;

Selector_2 s3278_6(wires_819_5[2], addr_819_5, addr_positional[13115:13112], addr_3278_6);

wire[27:0] addr_3279_6;

Selector_2 s3279_6(wires_819_5[3], addr_819_5, addr_positional[13119:13116], addr_3279_6);

wire[27:0] addr_3280_6;

Selector_2 s3280_6(wires_820_5[0], addr_820_5, addr_positional[13123:13120], addr_3280_6);

wire[27:0] addr_3281_6;

Selector_2 s3281_6(wires_820_5[1], addr_820_5, addr_positional[13127:13124], addr_3281_6);

wire[27:0] addr_3282_6;

Selector_2 s3282_6(wires_820_5[2], addr_820_5, addr_positional[13131:13128], addr_3282_6);

wire[27:0] addr_3283_6;

Selector_2 s3283_6(wires_820_5[3], addr_820_5, addr_positional[13135:13132], addr_3283_6);

wire[27:0] addr_3284_6;

Selector_2 s3284_6(wires_821_5[0], addr_821_5, addr_positional[13139:13136], addr_3284_6);

wire[27:0] addr_3285_6;

Selector_2 s3285_6(wires_821_5[1], addr_821_5, addr_positional[13143:13140], addr_3285_6);

wire[27:0] addr_3286_6;

Selector_2 s3286_6(wires_821_5[2], addr_821_5, addr_positional[13147:13144], addr_3286_6);

wire[27:0] addr_3287_6;

Selector_2 s3287_6(wires_821_5[3], addr_821_5, addr_positional[13151:13148], addr_3287_6);

wire[27:0] addr_3288_6;

Selector_2 s3288_6(wires_822_5[0], addr_822_5, addr_positional[13155:13152], addr_3288_6);

wire[27:0] addr_3289_6;

Selector_2 s3289_6(wires_822_5[1], addr_822_5, addr_positional[13159:13156], addr_3289_6);

wire[27:0] addr_3290_6;

Selector_2 s3290_6(wires_822_5[2], addr_822_5, addr_positional[13163:13160], addr_3290_6);

wire[27:0] addr_3291_6;

Selector_2 s3291_6(wires_822_5[3], addr_822_5, addr_positional[13167:13164], addr_3291_6);

wire[27:0] addr_3292_6;

Selector_2 s3292_6(wires_823_5[0], addr_823_5, addr_positional[13171:13168], addr_3292_6);

wire[27:0] addr_3293_6;

Selector_2 s3293_6(wires_823_5[1], addr_823_5, addr_positional[13175:13172], addr_3293_6);

wire[27:0] addr_3294_6;

Selector_2 s3294_6(wires_823_5[2], addr_823_5, addr_positional[13179:13176], addr_3294_6);

wire[27:0] addr_3295_6;

Selector_2 s3295_6(wires_823_5[3], addr_823_5, addr_positional[13183:13180], addr_3295_6);

wire[27:0] addr_3296_6;

Selector_2 s3296_6(wires_824_5[0], addr_824_5, addr_positional[13187:13184], addr_3296_6);

wire[27:0] addr_3297_6;

Selector_2 s3297_6(wires_824_5[1], addr_824_5, addr_positional[13191:13188], addr_3297_6);

wire[27:0] addr_3298_6;

Selector_2 s3298_6(wires_824_5[2], addr_824_5, addr_positional[13195:13192], addr_3298_6);

wire[27:0] addr_3299_6;

Selector_2 s3299_6(wires_824_5[3], addr_824_5, addr_positional[13199:13196], addr_3299_6);

wire[27:0] addr_3300_6;

Selector_2 s3300_6(wires_825_5[0], addr_825_5, addr_positional[13203:13200], addr_3300_6);

wire[27:0] addr_3301_6;

Selector_2 s3301_6(wires_825_5[1], addr_825_5, addr_positional[13207:13204], addr_3301_6);

wire[27:0] addr_3302_6;

Selector_2 s3302_6(wires_825_5[2], addr_825_5, addr_positional[13211:13208], addr_3302_6);

wire[27:0] addr_3303_6;

Selector_2 s3303_6(wires_825_5[3], addr_825_5, addr_positional[13215:13212], addr_3303_6);

wire[27:0] addr_3304_6;

Selector_2 s3304_6(wires_826_5[0], addr_826_5, addr_positional[13219:13216], addr_3304_6);

wire[27:0] addr_3305_6;

Selector_2 s3305_6(wires_826_5[1], addr_826_5, addr_positional[13223:13220], addr_3305_6);

wire[27:0] addr_3306_6;

Selector_2 s3306_6(wires_826_5[2], addr_826_5, addr_positional[13227:13224], addr_3306_6);

wire[27:0] addr_3307_6;

Selector_2 s3307_6(wires_826_5[3], addr_826_5, addr_positional[13231:13228], addr_3307_6);

wire[27:0] addr_3308_6;

Selector_2 s3308_6(wires_827_5[0], addr_827_5, addr_positional[13235:13232], addr_3308_6);

wire[27:0] addr_3309_6;

Selector_2 s3309_6(wires_827_5[1], addr_827_5, addr_positional[13239:13236], addr_3309_6);

wire[27:0] addr_3310_6;

Selector_2 s3310_6(wires_827_5[2], addr_827_5, addr_positional[13243:13240], addr_3310_6);

wire[27:0] addr_3311_6;

Selector_2 s3311_6(wires_827_5[3], addr_827_5, addr_positional[13247:13244], addr_3311_6);

wire[27:0] addr_3312_6;

Selector_2 s3312_6(wires_828_5[0], addr_828_5, addr_positional[13251:13248], addr_3312_6);

wire[27:0] addr_3313_6;

Selector_2 s3313_6(wires_828_5[1], addr_828_5, addr_positional[13255:13252], addr_3313_6);

wire[27:0] addr_3314_6;

Selector_2 s3314_6(wires_828_5[2], addr_828_5, addr_positional[13259:13256], addr_3314_6);

wire[27:0] addr_3315_6;

Selector_2 s3315_6(wires_828_5[3], addr_828_5, addr_positional[13263:13260], addr_3315_6);

wire[27:0] addr_3316_6;

Selector_2 s3316_6(wires_829_5[0], addr_829_5, addr_positional[13267:13264], addr_3316_6);

wire[27:0] addr_3317_6;

Selector_2 s3317_6(wires_829_5[1], addr_829_5, addr_positional[13271:13268], addr_3317_6);

wire[27:0] addr_3318_6;

Selector_2 s3318_6(wires_829_5[2], addr_829_5, addr_positional[13275:13272], addr_3318_6);

wire[27:0] addr_3319_6;

Selector_2 s3319_6(wires_829_5[3], addr_829_5, addr_positional[13279:13276], addr_3319_6);

wire[27:0] addr_3320_6;

Selector_2 s3320_6(wires_830_5[0], addr_830_5, addr_positional[13283:13280], addr_3320_6);

wire[27:0] addr_3321_6;

Selector_2 s3321_6(wires_830_5[1], addr_830_5, addr_positional[13287:13284], addr_3321_6);

wire[27:0] addr_3322_6;

Selector_2 s3322_6(wires_830_5[2], addr_830_5, addr_positional[13291:13288], addr_3322_6);

wire[27:0] addr_3323_6;

Selector_2 s3323_6(wires_830_5[3], addr_830_5, addr_positional[13295:13292], addr_3323_6);

wire[27:0] addr_3324_6;

Selector_2 s3324_6(wires_831_5[0], addr_831_5, addr_positional[13299:13296], addr_3324_6);

wire[27:0] addr_3325_6;

Selector_2 s3325_6(wires_831_5[1], addr_831_5, addr_positional[13303:13300], addr_3325_6);

wire[27:0] addr_3326_6;

Selector_2 s3326_6(wires_831_5[2], addr_831_5, addr_positional[13307:13304], addr_3326_6);

wire[27:0] addr_3327_6;

Selector_2 s3327_6(wires_831_5[3], addr_831_5, addr_positional[13311:13308], addr_3327_6);

wire[27:0] addr_3328_6;

Selector_2 s3328_6(wires_832_5[0], addr_832_5, addr_positional[13315:13312], addr_3328_6);

wire[27:0] addr_3329_6;

Selector_2 s3329_6(wires_832_5[1], addr_832_5, addr_positional[13319:13316], addr_3329_6);

wire[27:0] addr_3330_6;

Selector_2 s3330_6(wires_832_5[2], addr_832_5, addr_positional[13323:13320], addr_3330_6);

wire[27:0] addr_3331_6;

Selector_2 s3331_6(wires_832_5[3], addr_832_5, addr_positional[13327:13324], addr_3331_6);

wire[27:0] addr_3332_6;

Selector_2 s3332_6(wires_833_5[0], addr_833_5, addr_positional[13331:13328], addr_3332_6);

wire[27:0] addr_3333_6;

Selector_2 s3333_6(wires_833_5[1], addr_833_5, addr_positional[13335:13332], addr_3333_6);

wire[27:0] addr_3334_6;

Selector_2 s3334_6(wires_833_5[2], addr_833_5, addr_positional[13339:13336], addr_3334_6);

wire[27:0] addr_3335_6;

Selector_2 s3335_6(wires_833_5[3], addr_833_5, addr_positional[13343:13340], addr_3335_6);

wire[27:0] addr_3336_6;

Selector_2 s3336_6(wires_834_5[0], addr_834_5, addr_positional[13347:13344], addr_3336_6);

wire[27:0] addr_3337_6;

Selector_2 s3337_6(wires_834_5[1], addr_834_5, addr_positional[13351:13348], addr_3337_6);

wire[27:0] addr_3338_6;

Selector_2 s3338_6(wires_834_5[2], addr_834_5, addr_positional[13355:13352], addr_3338_6);

wire[27:0] addr_3339_6;

Selector_2 s3339_6(wires_834_5[3], addr_834_5, addr_positional[13359:13356], addr_3339_6);

wire[27:0] addr_3340_6;

Selector_2 s3340_6(wires_835_5[0], addr_835_5, addr_positional[13363:13360], addr_3340_6);

wire[27:0] addr_3341_6;

Selector_2 s3341_6(wires_835_5[1], addr_835_5, addr_positional[13367:13364], addr_3341_6);

wire[27:0] addr_3342_6;

Selector_2 s3342_6(wires_835_5[2], addr_835_5, addr_positional[13371:13368], addr_3342_6);

wire[27:0] addr_3343_6;

Selector_2 s3343_6(wires_835_5[3], addr_835_5, addr_positional[13375:13372], addr_3343_6);

wire[27:0] addr_3344_6;

Selector_2 s3344_6(wires_836_5[0], addr_836_5, addr_positional[13379:13376], addr_3344_6);

wire[27:0] addr_3345_6;

Selector_2 s3345_6(wires_836_5[1], addr_836_5, addr_positional[13383:13380], addr_3345_6);

wire[27:0] addr_3346_6;

Selector_2 s3346_6(wires_836_5[2], addr_836_5, addr_positional[13387:13384], addr_3346_6);

wire[27:0] addr_3347_6;

Selector_2 s3347_6(wires_836_5[3], addr_836_5, addr_positional[13391:13388], addr_3347_6);

wire[27:0] addr_3348_6;

Selector_2 s3348_6(wires_837_5[0], addr_837_5, addr_positional[13395:13392], addr_3348_6);

wire[27:0] addr_3349_6;

Selector_2 s3349_6(wires_837_5[1], addr_837_5, addr_positional[13399:13396], addr_3349_6);

wire[27:0] addr_3350_6;

Selector_2 s3350_6(wires_837_5[2], addr_837_5, addr_positional[13403:13400], addr_3350_6);

wire[27:0] addr_3351_6;

Selector_2 s3351_6(wires_837_5[3], addr_837_5, addr_positional[13407:13404], addr_3351_6);

wire[27:0] addr_3352_6;

Selector_2 s3352_6(wires_838_5[0], addr_838_5, addr_positional[13411:13408], addr_3352_6);

wire[27:0] addr_3353_6;

Selector_2 s3353_6(wires_838_5[1], addr_838_5, addr_positional[13415:13412], addr_3353_6);

wire[27:0] addr_3354_6;

Selector_2 s3354_6(wires_838_5[2], addr_838_5, addr_positional[13419:13416], addr_3354_6);

wire[27:0] addr_3355_6;

Selector_2 s3355_6(wires_838_5[3], addr_838_5, addr_positional[13423:13420], addr_3355_6);

wire[27:0] addr_3356_6;

Selector_2 s3356_6(wires_839_5[0], addr_839_5, addr_positional[13427:13424], addr_3356_6);

wire[27:0] addr_3357_6;

Selector_2 s3357_6(wires_839_5[1], addr_839_5, addr_positional[13431:13428], addr_3357_6);

wire[27:0] addr_3358_6;

Selector_2 s3358_6(wires_839_5[2], addr_839_5, addr_positional[13435:13432], addr_3358_6);

wire[27:0] addr_3359_6;

Selector_2 s3359_6(wires_839_5[3], addr_839_5, addr_positional[13439:13436], addr_3359_6);

wire[27:0] addr_3360_6;

Selector_2 s3360_6(wires_840_5[0], addr_840_5, addr_positional[13443:13440], addr_3360_6);

wire[27:0] addr_3361_6;

Selector_2 s3361_6(wires_840_5[1], addr_840_5, addr_positional[13447:13444], addr_3361_6);

wire[27:0] addr_3362_6;

Selector_2 s3362_6(wires_840_5[2], addr_840_5, addr_positional[13451:13448], addr_3362_6);

wire[27:0] addr_3363_6;

Selector_2 s3363_6(wires_840_5[3], addr_840_5, addr_positional[13455:13452], addr_3363_6);

wire[27:0] addr_3364_6;

Selector_2 s3364_6(wires_841_5[0], addr_841_5, addr_positional[13459:13456], addr_3364_6);

wire[27:0] addr_3365_6;

Selector_2 s3365_6(wires_841_5[1], addr_841_5, addr_positional[13463:13460], addr_3365_6);

wire[27:0] addr_3366_6;

Selector_2 s3366_6(wires_841_5[2], addr_841_5, addr_positional[13467:13464], addr_3366_6);

wire[27:0] addr_3367_6;

Selector_2 s3367_6(wires_841_5[3], addr_841_5, addr_positional[13471:13468], addr_3367_6);

wire[27:0] addr_3368_6;

Selector_2 s3368_6(wires_842_5[0], addr_842_5, addr_positional[13475:13472], addr_3368_6);

wire[27:0] addr_3369_6;

Selector_2 s3369_6(wires_842_5[1], addr_842_5, addr_positional[13479:13476], addr_3369_6);

wire[27:0] addr_3370_6;

Selector_2 s3370_6(wires_842_5[2], addr_842_5, addr_positional[13483:13480], addr_3370_6);

wire[27:0] addr_3371_6;

Selector_2 s3371_6(wires_842_5[3], addr_842_5, addr_positional[13487:13484], addr_3371_6);

wire[27:0] addr_3372_6;

Selector_2 s3372_6(wires_843_5[0], addr_843_5, addr_positional[13491:13488], addr_3372_6);

wire[27:0] addr_3373_6;

Selector_2 s3373_6(wires_843_5[1], addr_843_5, addr_positional[13495:13492], addr_3373_6);

wire[27:0] addr_3374_6;

Selector_2 s3374_6(wires_843_5[2], addr_843_5, addr_positional[13499:13496], addr_3374_6);

wire[27:0] addr_3375_6;

Selector_2 s3375_6(wires_843_5[3], addr_843_5, addr_positional[13503:13500], addr_3375_6);

wire[27:0] addr_3376_6;

Selector_2 s3376_6(wires_844_5[0], addr_844_5, addr_positional[13507:13504], addr_3376_6);

wire[27:0] addr_3377_6;

Selector_2 s3377_6(wires_844_5[1], addr_844_5, addr_positional[13511:13508], addr_3377_6);

wire[27:0] addr_3378_6;

Selector_2 s3378_6(wires_844_5[2], addr_844_5, addr_positional[13515:13512], addr_3378_6);

wire[27:0] addr_3379_6;

Selector_2 s3379_6(wires_844_5[3], addr_844_5, addr_positional[13519:13516], addr_3379_6);

wire[27:0] addr_3380_6;

Selector_2 s3380_6(wires_845_5[0], addr_845_5, addr_positional[13523:13520], addr_3380_6);

wire[27:0] addr_3381_6;

Selector_2 s3381_6(wires_845_5[1], addr_845_5, addr_positional[13527:13524], addr_3381_6);

wire[27:0] addr_3382_6;

Selector_2 s3382_6(wires_845_5[2], addr_845_5, addr_positional[13531:13528], addr_3382_6);

wire[27:0] addr_3383_6;

Selector_2 s3383_6(wires_845_5[3], addr_845_5, addr_positional[13535:13532], addr_3383_6);

wire[27:0] addr_3384_6;

Selector_2 s3384_6(wires_846_5[0], addr_846_5, addr_positional[13539:13536], addr_3384_6);

wire[27:0] addr_3385_6;

Selector_2 s3385_6(wires_846_5[1], addr_846_5, addr_positional[13543:13540], addr_3385_6);

wire[27:0] addr_3386_6;

Selector_2 s3386_6(wires_846_5[2], addr_846_5, addr_positional[13547:13544], addr_3386_6);

wire[27:0] addr_3387_6;

Selector_2 s3387_6(wires_846_5[3], addr_846_5, addr_positional[13551:13548], addr_3387_6);

wire[27:0] addr_3388_6;

Selector_2 s3388_6(wires_847_5[0], addr_847_5, addr_positional[13555:13552], addr_3388_6);

wire[27:0] addr_3389_6;

Selector_2 s3389_6(wires_847_5[1], addr_847_5, addr_positional[13559:13556], addr_3389_6);

wire[27:0] addr_3390_6;

Selector_2 s3390_6(wires_847_5[2], addr_847_5, addr_positional[13563:13560], addr_3390_6);

wire[27:0] addr_3391_6;

Selector_2 s3391_6(wires_847_5[3], addr_847_5, addr_positional[13567:13564], addr_3391_6);

wire[27:0] addr_3392_6;

Selector_2 s3392_6(wires_848_5[0], addr_848_5, addr_positional[13571:13568], addr_3392_6);

wire[27:0] addr_3393_6;

Selector_2 s3393_6(wires_848_5[1], addr_848_5, addr_positional[13575:13572], addr_3393_6);

wire[27:0] addr_3394_6;

Selector_2 s3394_6(wires_848_5[2], addr_848_5, addr_positional[13579:13576], addr_3394_6);

wire[27:0] addr_3395_6;

Selector_2 s3395_6(wires_848_5[3], addr_848_5, addr_positional[13583:13580], addr_3395_6);

wire[27:0] addr_3396_6;

Selector_2 s3396_6(wires_849_5[0], addr_849_5, addr_positional[13587:13584], addr_3396_6);

wire[27:0] addr_3397_6;

Selector_2 s3397_6(wires_849_5[1], addr_849_5, addr_positional[13591:13588], addr_3397_6);

wire[27:0] addr_3398_6;

Selector_2 s3398_6(wires_849_5[2], addr_849_5, addr_positional[13595:13592], addr_3398_6);

wire[27:0] addr_3399_6;

Selector_2 s3399_6(wires_849_5[3], addr_849_5, addr_positional[13599:13596], addr_3399_6);

wire[27:0] addr_3400_6;

Selector_2 s3400_6(wires_850_5[0], addr_850_5, addr_positional[13603:13600], addr_3400_6);

wire[27:0] addr_3401_6;

Selector_2 s3401_6(wires_850_5[1], addr_850_5, addr_positional[13607:13604], addr_3401_6);

wire[27:0] addr_3402_6;

Selector_2 s3402_6(wires_850_5[2], addr_850_5, addr_positional[13611:13608], addr_3402_6);

wire[27:0] addr_3403_6;

Selector_2 s3403_6(wires_850_5[3], addr_850_5, addr_positional[13615:13612], addr_3403_6);

wire[27:0] addr_3404_6;

Selector_2 s3404_6(wires_851_5[0], addr_851_5, addr_positional[13619:13616], addr_3404_6);

wire[27:0] addr_3405_6;

Selector_2 s3405_6(wires_851_5[1], addr_851_5, addr_positional[13623:13620], addr_3405_6);

wire[27:0] addr_3406_6;

Selector_2 s3406_6(wires_851_5[2], addr_851_5, addr_positional[13627:13624], addr_3406_6);

wire[27:0] addr_3407_6;

Selector_2 s3407_6(wires_851_5[3], addr_851_5, addr_positional[13631:13628], addr_3407_6);

wire[27:0] addr_3408_6;

Selector_2 s3408_6(wires_852_5[0], addr_852_5, addr_positional[13635:13632], addr_3408_6);

wire[27:0] addr_3409_6;

Selector_2 s3409_6(wires_852_5[1], addr_852_5, addr_positional[13639:13636], addr_3409_6);

wire[27:0] addr_3410_6;

Selector_2 s3410_6(wires_852_5[2], addr_852_5, addr_positional[13643:13640], addr_3410_6);

wire[27:0] addr_3411_6;

Selector_2 s3411_6(wires_852_5[3], addr_852_5, addr_positional[13647:13644], addr_3411_6);

wire[27:0] addr_3412_6;

Selector_2 s3412_6(wires_853_5[0], addr_853_5, addr_positional[13651:13648], addr_3412_6);

wire[27:0] addr_3413_6;

Selector_2 s3413_6(wires_853_5[1], addr_853_5, addr_positional[13655:13652], addr_3413_6);

wire[27:0] addr_3414_6;

Selector_2 s3414_6(wires_853_5[2], addr_853_5, addr_positional[13659:13656], addr_3414_6);

wire[27:0] addr_3415_6;

Selector_2 s3415_6(wires_853_5[3], addr_853_5, addr_positional[13663:13660], addr_3415_6);

wire[27:0] addr_3416_6;

Selector_2 s3416_6(wires_854_5[0], addr_854_5, addr_positional[13667:13664], addr_3416_6);

wire[27:0] addr_3417_6;

Selector_2 s3417_6(wires_854_5[1], addr_854_5, addr_positional[13671:13668], addr_3417_6);

wire[27:0] addr_3418_6;

Selector_2 s3418_6(wires_854_5[2], addr_854_5, addr_positional[13675:13672], addr_3418_6);

wire[27:0] addr_3419_6;

Selector_2 s3419_6(wires_854_5[3], addr_854_5, addr_positional[13679:13676], addr_3419_6);

wire[27:0] addr_3420_6;

Selector_2 s3420_6(wires_855_5[0], addr_855_5, addr_positional[13683:13680], addr_3420_6);

wire[27:0] addr_3421_6;

Selector_2 s3421_6(wires_855_5[1], addr_855_5, addr_positional[13687:13684], addr_3421_6);

wire[27:0] addr_3422_6;

Selector_2 s3422_6(wires_855_5[2], addr_855_5, addr_positional[13691:13688], addr_3422_6);

wire[27:0] addr_3423_6;

Selector_2 s3423_6(wires_855_5[3], addr_855_5, addr_positional[13695:13692], addr_3423_6);

wire[27:0] addr_3424_6;

Selector_2 s3424_6(wires_856_5[0], addr_856_5, addr_positional[13699:13696], addr_3424_6);

wire[27:0] addr_3425_6;

Selector_2 s3425_6(wires_856_5[1], addr_856_5, addr_positional[13703:13700], addr_3425_6);

wire[27:0] addr_3426_6;

Selector_2 s3426_6(wires_856_5[2], addr_856_5, addr_positional[13707:13704], addr_3426_6);

wire[27:0] addr_3427_6;

Selector_2 s3427_6(wires_856_5[3], addr_856_5, addr_positional[13711:13708], addr_3427_6);

wire[27:0] addr_3428_6;

Selector_2 s3428_6(wires_857_5[0], addr_857_5, addr_positional[13715:13712], addr_3428_6);

wire[27:0] addr_3429_6;

Selector_2 s3429_6(wires_857_5[1], addr_857_5, addr_positional[13719:13716], addr_3429_6);

wire[27:0] addr_3430_6;

Selector_2 s3430_6(wires_857_5[2], addr_857_5, addr_positional[13723:13720], addr_3430_6);

wire[27:0] addr_3431_6;

Selector_2 s3431_6(wires_857_5[3], addr_857_5, addr_positional[13727:13724], addr_3431_6);

wire[27:0] addr_3432_6;

Selector_2 s3432_6(wires_858_5[0], addr_858_5, addr_positional[13731:13728], addr_3432_6);

wire[27:0] addr_3433_6;

Selector_2 s3433_6(wires_858_5[1], addr_858_5, addr_positional[13735:13732], addr_3433_6);

wire[27:0] addr_3434_6;

Selector_2 s3434_6(wires_858_5[2], addr_858_5, addr_positional[13739:13736], addr_3434_6);

wire[27:0] addr_3435_6;

Selector_2 s3435_6(wires_858_5[3], addr_858_5, addr_positional[13743:13740], addr_3435_6);

wire[27:0] addr_3436_6;

Selector_2 s3436_6(wires_859_5[0], addr_859_5, addr_positional[13747:13744], addr_3436_6);

wire[27:0] addr_3437_6;

Selector_2 s3437_6(wires_859_5[1], addr_859_5, addr_positional[13751:13748], addr_3437_6);

wire[27:0] addr_3438_6;

Selector_2 s3438_6(wires_859_5[2], addr_859_5, addr_positional[13755:13752], addr_3438_6);

wire[27:0] addr_3439_6;

Selector_2 s3439_6(wires_859_5[3], addr_859_5, addr_positional[13759:13756], addr_3439_6);

wire[27:0] addr_3440_6;

Selector_2 s3440_6(wires_860_5[0], addr_860_5, addr_positional[13763:13760], addr_3440_6);

wire[27:0] addr_3441_6;

Selector_2 s3441_6(wires_860_5[1], addr_860_5, addr_positional[13767:13764], addr_3441_6);

wire[27:0] addr_3442_6;

Selector_2 s3442_6(wires_860_5[2], addr_860_5, addr_positional[13771:13768], addr_3442_6);

wire[27:0] addr_3443_6;

Selector_2 s3443_6(wires_860_5[3], addr_860_5, addr_positional[13775:13772], addr_3443_6);

wire[27:0] addr_3444_6;

Selector_2 s3444_6(wires_861_5[0], addr_861_5, addr_positional[13779:13776], addr_3444_6);

wire[27:0] addr_3445_6;

Selector_2 s3445_6(wires_861_5[1], addr_861_5, addr_positional[13783:13780], addr_3445_6);

wire[27:0] addr_3446_6;

Selector_2 s3446_6(wires_861_5[2], addr_861_5, addr_positional[13787:13784], addr_3446_6);

wire[27:0] addr_3447_6;

Selector_2 s3447_6(wires_861_5[3], addr_861_5, addr_positional[13791:13788], addr_3447_6);

wire[27:0] addr_3448_6;

Selector_2 s3448_6(wires_862_5[0], addr_862_5, addr_positional[13795:13792], addr_3448_6);

wire[27:0] addr_3449_6;

Selector_2 s3449_6(wires_862_5[1], addr_862_5, addr_positional[13799:13796], addr_3449_6);

wire[27:0] addr_3450_6;

Selector_2 s3450_6(wires_862_5[2], addr_862_5, addr_positional[13803:13800], addr_3450_6);

wire[27:0] addr_3451_6;

Selector_2 s3451_6(wires_862_5[3], addr_862_5, addr_positional[13807:13804], addr_3451_6);

wire[27:0] addr_3452_6;

Selector_2 s3452_6(wires_863_5[0], addr_863_5, addr_positional[13811:13808], addr_3452_6);

wire[27:0] addr_3453_6;

Selector_2 s3453_6(wires_863_5[1], addr_863_5, addr_positional[13815:13812], addr_3453_6);

wire[27:0] addr_3454_6;

Selector_2 s3454_6(wires_863_5[2], addr_863_5, addr_positional[13819:13816], addr_3454_6);

wire[27:0] addr_3455_6;

Selector_2 s3455_6(wires_863_5[3], addr_863_5, addr_positional[13823:13820], addr_3455_6);

wire[27:0] addr_3456_6;

Selector_2 s3456_6(wires_864_5[0], addr_864_5, addr_positional[13827:13824], addr_3456_6);

wire[27:0] addr_3457_6;

Selector_2 s3457_6(wires_864_5[1], addr_864_5, addr_positional[13831:13828], addr_3457_6);

wire[27:0] addr_3458_6;

Selector_2 s3458_6(wires_864_5[2], addr_864_5, addr_positional[13835:13832], addr_3458_6);

wire[27:0] addr_3459_6;

Selector_2 s3459_6(wires_864_5[3], addr_864_5, addr_positional[13839:13836], addr_3459_6);

wire[27:0] addr_3460_6;

Selector_2 s3460_6(wires_865_5[0], addr_865_5, addr_positional[13843:13840], addr_3460_6);

wire[27:0] addr_3461_6;

Selector_2 s3461_6(wires_865_5[1], addr_865_5, addr_positional[13847:13844], addr_3461_6);

wire[27:0] addr_3462_6;

Selector_2 s3462_6(wires_865_5[2], addr_865_5, addr_positional[13851:13848], addr_3462_6);

wire[27:0] addr_3463_6;

Selector_2 s3463_6(wires_865_5[3], addr_865_5, addr_positional[13855:13852], addr_3463_6);

wire[27:0] addr_3464_6;

Selector_2 s3464_6(wires_866_5[0], addr_866_5, addr_positional[13859:13856], addr_3464_6);

wire[27:0] addr_3465_6;

Selector_2 s3465_6(wires_866_5[1], addr_866_5, addr_positional[13863:13860], addr_3465_6);

wire[27:0] addr_3466_6;

Selector_2 s3466_6(wires_866_5[2], addr_866_5, addr_positional[13867:13864], addr_3466_6);

wire[27:0] addr_3467_6;

Selector_2 s3467_6(wires_866_5[3], addr_866_5, addr_positional[13871:13868], addr_3467_6);

wire[27:0] addr_3468_6;

Selector_2 s3468_6(wires_867_5[0], addr_867_5, addr_positional[13875:13872], addr_3468_6);

wire[27:0] addr_3469_6;

Selector_2 s3469_6(wires_867_5[1], addr_867_5, addr_positional[13879:13876], addr_3469_6);

wire[27:0] addr_3470_6;

Selector_2 s3470_6(wires_867_5[2], addr_867_5, addr_positional[13883:13880], addr_3470_6);

wire[27:0] addr_3471_6;

Selector_2 s3471_6(wires_867_5[3], addr_867_5, addr_positional[13887:13884], addr_3471_6);

wire[27:0] addr_3472_6;

Selector_2 s3472_6(wires_868_5[0], addr_868_5, addr_positional[13891:13888], addr_3472_6);

wire[27:0] addr_3473_6;

Selector_2 s3473_6(wires_868_5[1], addr_868_5, addr_positional[13895:13892], addr_3473_6);

wire[27:0] addr_3474_6;

Selector_2 s3474_6(wires_868_5[2], addr_868_5, addr_positional[13899:13896], addr_3474_6);

wire[27:0] addr_3475_6;

Selector_2 s3475_6(wires_868_5[3], addr_868_5, addr_positional[13903:13900], addr_3475_6);

wire[27:0] addr_3476_6;

Selector_2 s3476_6(wires_869_5[0], addr_869_5, addr_positional[13907:13904], addr_3476_6);

wire[27:0] addr_3477_6;

Selector_2 s3477_6(wires_869_5[1], addr_869_5, addr_positional[13911:13908], addr_3477_6);

wire[27:0] addr_3478_6;

Selector_2 s3478_6(wires_869_5[2], addr_869_5, addr_positional[13915:13912], addr_3478_6);

wire[27:0] addr_3479_6;

Selector_2 s3479_6(wires_869_5[3], addr_869_5, addr_positional[13919:13916], addr_3479_6);

wire[27:0] addr_3480_6;

Selector_2 s3480_6(wires_870_5[0], addr_870_5, addr_positional[13923:13920], addr_3480_6);

wire[27:0] addr_3481_6;

Selector_2 s3481_6(wires_870_5[1], addr_870_5, addr_positional[13927:13924], addr_3481_6);

wire[27:0] addr_3482_6;

Selector_2 s3482_6(wires_870_5[2], addr_870_5, addr_positional[13931:13928], addr_3482_6);

wire[27:0] addr_3483_6;

Selector_2 s3483_6(wires_870_5[3], addr_870_5, addr_positional[13935:13932], addr_3483_6);

wire[27:0] addr_3484_6;

Selector_2 s3484_6(wires_871_5[0], addr_871_5, addr_positional[13939:13936], addr_3484_6);

wire[27:0] addr_3485_6;

Selector_2 s3485_6(wires_871_5[1], addr_871_5, addr_positional[13943:13940], addr_3485_6);

wire[27:0] addr_3486_6;

Selector_2 s3486_6(wires_871_5[2], addr_871_5, addr_positional[13947:13944], addr_3486_6);

wire[27:0] addr_3487_6;

Selector_2 s3487_6(wires_871_5[3], addr_871_5, addr_positional[13951:13948], addr_3487_6);

wire[27:0] addr_3488_6;

Selector_2 s3488_6(wires_872_5[0], addr_872_5, addr_positional[13955:13952], addr_3488_6);

wire[27:0] addr_3489_6;

Selector_2 s3489_6(wires_872_5[1], addr_872_5, addr_positional[13959:13956], addr_3489_6);

wire[27:0] addr_3490_6;

Selector_2 s3490_6(wires_872_5[2], addr_872_5, addr_positional[13963:13960], addr_3490_6);

wire[27:0] addr_3491_6;

Selector_2 s3491_6(wires_872_5[3], addr_872_5, addr_positional[13967:13964], addr_3491_6);

wire[27:0] addr_3492_6;

Selector_2 s3492_6(wires_873_5[0], addr_873_5, addr_positional[13971:13968], addr_3492_6);

wire[27:0] addr_3493_6;

Selector_2 s3493_6(wires_873_5[1], addr_873_5, addr_positional[13975:13972], addr_3493_6);

wire[27:0] addr_3494_6;

Selector_2 s3494_6(wires_873_5[2], addr_873_5, addr_positional[13979:13976], addr_3494_6);

wire[27:0] addr_3495_6;

Selector_2 s3495_6(wires_873_5[3], addr_873_5, addr_positional[13983:13980], addr_3495_6);

wire[27:0] addr_3496_6;

Selector_2 s3496_6(wires_874_5[0], addr_874_5, addr_positional[13987:13984], addr_3496_6);

wire[27:0] addr_3497_6;

Selector_2 s3497_6(wires_874_5[1], addr_874_5, addr_positional[13991:13988], addr_3497_6);

wire[27:0] addr_3498_6;

Selector_2 s3498_6(wires_874_5[2], addr_874_5, addr_positional[13995:13992], addr_3498_6);

wire[27:0] addr_3499_6;

Selector_2 s3499_6(wires_874_5[3], addr_874_5, addr_positional[13999:13996], addr_3499_6);

wire[27:0] addr_3500_6;

Selector_2 s3500_6(wires_875_5[0], addr_875_5, addr_positional[14003:14000], addr_3500_6);

wire[27:0] addr_3501_6;

Selector_2 s3501_6(wires_875_5[1], addr_875_5, addr_positional[14007:14004], addr_3501_6);

wire[27:0] addr_3502_6;

Selector_2 s3502_6(wires_875_5[2], addr_875_5, addr_positional[14011:14008], addr_3502_6);

wire[27:0] addr_3503_6;

Selector_2 s3503_6(wires_875_5[3], addr_875_5, addr_positional[14015:14012], addr_3503_6);

wire[27:0] addr_3504_6;

Selector_2 s3504_6(wires_876_5[0], addr_876_5, addr_positional[14019:14016], addr_3504_6);

wire[27:0] addr_3505_6;

Selector_2 s3505_6(wires_876_5[1], addr_876_5, addr_positional[14023:14020], addr_3505_6);

wire[27:0] addr_3506_6;

Selector_2 s3506_6(wires_876_5[2], addr_876_5, addr_positional[14027:14024], addr_3506_6);

wire[27:0] addr_3507_6;

Selector_2 s3507_6(wires_876_5[3], addr_876_5, addr_positional[14031:14028], addr_3507_6);

wire[27:0] addr_3508_6;

Selector_2 s3508_6(wires_877_5[0], addr_877_5, addr_positional[14035:14032], addr_3508_6);

wire[27:0] addr_3509_6;

Selector_2 s3509_6(wires_877_5[1], addr_877_5, addr_positional[14039:14036], addr_3509_6);

wire[27:0] addr_3510_6;

Selector_2 s3510_6(wires_877_5[2], addr_877_5, addr_positional[14043:14040], addr_3510_6);

wire[27:0] addr_3511_6;

Selector_2 s3511_6(wires_877_5[3], addr_877_5, addr_positional[14047:14044], addr_3511_6);

wire[27:0] addr_3512_6;

Selector_2 s3512_6(wires_878_5[0], addr_878_5, addr_positional[14051:14048], addr_3512_6);

wire[27:0] addr_3513_6;

Selector_2 s3513_6(wires_878_5[1], addr_878_5, addr_positional[14055:14052], addr_3513_6);

wire[27:0] addr_3514_6;

Selector_2 s3514_6(wires_878_5[2], addr_878_5, addr_positional[14059:14056], addr_3514_6);

wire[27:0] addr_3515_6;

Selector_2 s3515_6(wires_878_5[3], addr_878_5, addr_positional[14063:14060], addr_3515_6);

wire[27:0] addr_3516_6;

Selector_2 s3516_6(wires_879_5[0], addr_879_5, addr_positional[14067:14064], addr_3516_6);

wire[27:0] addr_3517_6;

Selector_2 s3517_6(wires_879_5[1], addr_879_5, addr_positional[14071:14068], addr_3517_6);

wire[27:0] addr_3518_6;

Selector_2 s3518_6(wires_879_5[2], addr_879_5, addr_positional[14075:14072], addr_3518_6);

wire[27:0] addr_3519_6;

Selector_2 s3519_6(wires_879_5[3], addr_879_5, addr_positional[14079:14076], addr_3519_6);

wire[27:0] addr_3520_6;

Selector_2 s3520_6(wires_880_5[0], addr_880_5, addr_positional[14083:14080], addr_3520_6);

wire[27:0] addr_3521_6;

Selector_2 s3521_6(wires_880_5[1], addr_880_5, addr_positional[14087:14084], addr_3521_6);

wire[27:0] addr_3522_6;

Selector_2 s3522_6(wires_880_5[2], addr_880_5, addr_positional[14091:14088], addr_3522_6);

wire[27:0] addr_3523_6;

Selector_2 s3523_6(wires_880_5[3], addr_880_5, addr_positional[14095:14092], addr_3523_6);

wire[27:0] addr_3524_6;

Selector_2 s3524_6(wires_881_5[0], addr_881_5, addr_positional[14099:14096], addr_3524_6);

wire[27:0] addr_3525_6;

Selector_2 s3525_6(wires_881_5[1], addr_881_5, addr_positional[14103:14100], addr_3525_6);

wire[27:0] addr_3526_6;

Selector_2 s3526_6(wires_881_5[2], addr_881_5, addr_positional[14107:14104], addr_3526_6);

wire[27:0] addr_3527_6;

Selector_2 s3527_6(wires_881_5[3], addr_881_5, addr_positional[14111:14108], addr_3527_6);

wire[27:0] addr_3528_6;

Selector_2 s3528_6(wires_882_5[0], addr_882_5, addr_positional[14115:14112], addr_3528_6);

wire[27:0] addr_3529_6;

Selector_2 s3529_6(wires_882_5[1], addr_882_5, addr_positional[14119:14116], addr_3529_6);

wire[27:0] addr_3530_6;

Selector_2 s3530_6(wires_882_5[2], addr_882_5, addr_positional[14123:14120], addr_3530_6);

wire[27:0] addr_3531_6;

Selector_2 s3531_6(wires_882_5[3], addr_882_5, addr_positional[14127:14124], addr_3531_6);

wire[27:0] addr_3532_6;

Selector_2 s3532_6(wires_883_5[0], addr_883_5, addr_positional[14131:14128], addr_3532_6);

wire[27:0] addr_3533_6;

Selector_2 s3533_6(wires_883_5[1], addr_883_5, addr_positional[14135:14132], addr_3533_6);

wire[27:0] addr_3534_6;

Selector_2 s3534_6(wires_883_5[2], addr_883_5, addr_positional[14139:14136], addr_3534_6);

wire[27:0] addr_3535_6;

Selector_2 s3535_6(wires_883_5[3], addr_883_5, addr_positional[14143:14140], addr_3535_6);

wire[27:0] addr_3536_6;

Selector_2 s3536_6(wires_884_5[0], addr_884_5, addr_positional[14147:14144], addr_3536_6);

wire[27:0] addr_3537_6;

Selector_2 s3537_6(wires_884_5[1], addr_884_5, addr_positional[14151:14148], addr_3537_6);

wire[27:0] addr_3538_6;

Selector_2 s3538_6(wires_884_5[2], addr_884_5, addr_positional[14155:14152], addr_3538_6);

wire[27:0] addr_3539_6;

Selector_2 s3539_6(wires_884_5[3], addr_884_5, addr_positional[14159:14156], addr_3539_6);

wire[27:0] addr_3540_6;

Selector_2 s3540_6(wires_885_5[0], addr_885_5, addr_positional[14163:14160], addr_3540_6);

wire[27:0] addr_3541_6;

Selector_2 s3541_6(wires_885_5[1], addr_885_5, addr_positional[14167:14164], addr_3541_6);

wire[27:0] addr_3542_6;

Selector_2 s3542_6(wires_885_5[2], addr_885_5, addr_positional[14171:14168], addr_3542_6);

wire[27:0] addr_3543_6;

Selector_2 s3543_6(wires_885_5[3], addr_885_5, addr_positional[14175:14172], addr_3543_6);

wire[27:0] addr_3544_6;

Selector_2 s3544_6(wires_886_5[0], addr_886_5, addr_positional[14179:14176], addr_3544_6);

wire[27:0] addr_3545_6;

Selector_2 s3545_6(wires_886_5[1], addr_886_5, addr_positional[14183:14180], addr_3545_6);

wire[27:0] addr_3546_6;

Selector_2 s3546_6(wires_886_5[2], addr_886_5, addr_positional[14187:14184], addr_3546_6);

wire[27:0] addr_3547_6;

Selector_2 s3547_6(wires_886_5[3], addr_886_5, addr_positional[14191:14188], addr_3547_6);

wire[27:0] addr_3548_6;

Selector_2 s3548_6(wires_887_5[0], addr_887_5, addr_positional[14195:14192], addr_3548_6);

wire[27:0] addr_3549_6;

Selector_2 s3549_6(wires_887_5[1], addr_887_5, addr_positional[14199:14196], addr_3549_6);

wire[27:0] addr_3550_6;

Selector_2 s3550_6(wires_887_5[2], addr_887_5, addr_positional[14203:14200], addr_3550_6);

wire[27:0] addr_3551_6;

Selector_2 s3551_6(wires_887_5[3], addr_887_5, addr_positional[14207:14204], addr_3551_6);

wire[27:0] addr_3552_6;

Selector_2 s3552_6(wires_888_5[0], addr_888_5, addr_positional[14211:14208], addr_3552_6);

wire[27:0] addr_3553_6;

Selector_2 s3553_6(wires_888_5[1], addr_888_5, addr_positional[14215:14212], addr_3553_6);

wire[27:0] addr_3554_6;

Selector_2 s3554_6(wires_888_5[2], addr_888_5, addr_positional[14219:14216], addr_3554_6);

wire[27:0] addr_3555_6;

Selector_2 s3555_6(wires_888_5[3], addr_888_5, addr_positional[14223:14220], addr_3555_6);

wire[27:0] addr_3556_6;

Selector_2 s3556_6(wires_889_5[0], addr_889_5, addr_positional[14227:14224], addr_3556_6);

wire[27:0] addr_3557_6;

Selector_2 s3557_6(wires_889_5[1], addr_889_5, addr_positional[14231:14228], addr_3557_6);

wire[27:0] addr_3558_6;

Selector_2 s3558_6(wires_889_5[2], addr_889_5, addr_positional[14235:14232], addr_3558_6);

wire[27:0] addr_3559_6;

Selector_2 s3559_6(wires_889_5[3], addr_889_5, addr_positional[14239:14236], addr_3559_6);

wire[27:0] addr_3560_6;

Selector_2 s3560_6(wires_890_5[0], addr_890_5, addr_positional[14243:14240], addr_3560_6);

wire[27:0] addr_3561_6;

Selector_2 s3561_6(wires_890_5[1], addr_890_5, addr_positional[14247:14244], addr_3561_6);

wire[27:0] addr_3562_6;

Selector_2 s3562_6(wires_890_5[2], addr_890_5, addr_positional[14251:14248], addr_3562_6);

wire[27:0] addr_3563_6;

Selector_2 s3563_6(wires_890_5[3], addr_890_5, addr_positional[14255:14252], addr_3563_6);

wire[27:0] addr_3564_6;

Selector_2 s3564_6(wires_891_5[0], addr_891_5, addr_positional[14259:14256], addr_3564_6);

wire[27:0] addr_3565_6;

Selector_2 s3565_6(wires_891_5[1], addr_891_5, addr_positional[14263:14260], addr_3565_6);

wire[27:0] addr_3566_6;

Selector_2 s3566_6(wires_891_5[2], addr_891_5, addr_positional[14267:14264], addr_3566_6);

wire[27:0] addr_3567_6;

Selector_2 s3567_6(wires_891_5[3], addr_891_5, addr_positional[14271:14268], addr_3567_6);

wire[27:0] addr_3568_6;

Selector_2 s3568_6(wires_892_5[0], addr_892_5, addr_positional[14275:14272], addr_3568_6);

wire[27:0] addr_3569_6;

Selector_2 s3569_6(wires_892_5[1], addr_892_5, addr_positional[14279:14276], addr_3569_6);

wire[27:0] addr_3570_6;

Selector_2 s3570_6(wires_892_5[2], addr_892_5, addr_positional[14283:14280], addr_3570_6);

wire[27:0] addr_3571_6;

Selector_2 s3571_6(wires_892_5[3], addr_892_5, addr_positional[14287:14284], addr_3571_6);

wire[27:0] addr_3572_6;

Selector_2 s3572_6(wires_893_5[0], addr_893_5, addr_positional[14291:14288], addr_3572_6);

wire[27:0] addr_3573_6;

Selector_2 s3573_6(wires_893_5[1], addr_893_5, addr_positional[14295:14292], addr_3573_6);

wire[27:0] addr_3574_6;

Selector_2 s3574_6(wires_893_5[2], addr_893_5, addr_positional[14299:14296], addr_3574_6);

wire[27:0] addr_3575_6;

Selector_2 s3575_6(wires_893_5[3], addr_893_5, addr_positional[14303:14300], addr_3575_6);

wire[27:0] addr_3576_6;

Selector_2 s3576_6(wires_894_5[0], addr_894_5, addr_positional[14307:14304], addr_3576_6);

wire[27:0] addr_3577_6;

Selector_2 s3577_6(wires_894_5[1], addr_894_5, addr_positional[14311:14308], addr_3577_6);

wire[27:0] addr_3578_6;

Selector_2 s3578_6(wires_894_5[2], addr_894_5, addr_positional[14315:14312], addr_3578_6);

wire[27:0] addr_3579_6;

Selector_2 s3579_6(wires_894_5[3], addr_894_5, addr_positional[14319:14316], addr_3579_6);

wire[27:0] addr_3580_6;

Selector_2 s3580_6(wires_895_5[0], addr_895_5, addr_positional[14323:14320], addr_3580_6);

wire[27:0] addr_3581_6;

Selector_2 s3581_6(wires_895_5[1], addr_895_5, addr_positional[14327:14324], addr_3581_6);

wire[27:0] addr_3582_6;

Selector_2 s3582_6(wires_895_5[2], addr_895_5, addr_positional[14331:14328], addr_3582_6);

wire[27:0] addr_3583_6;

Selector_2 s3583_6(wires_895_5[3], addr_895_5, addr_positional[14335:14332], addr_3583_6);

wire[27:0] addr_3584_6;

Selector_2 s3584_6(wires_896_5[0], addr_896_5, addr_positional[14339:14336], addr_3584_6);

wire[27:0] addr_3585_6;

Selector_2 s3585_6(wires_896_5[1], addr_896_5, addr_positional[14343:14340], addr_3585_6);

wire[27:0] addr_3586_6;

Selector_2 s3586_6(wires_896_5[2], addr_896_5, addr_positional[14347:14344], addr_3586_6);

wire[27:0] addr_3587_6;

Selector_2 s3587_6(wires_896_5[3], addr_896_5, addr_positional[14351:14348], addr_3587_6);

wire[27:0] addr_3588_6;

Selector_2 s3588_6(wires_897_5[0], addr_897_5, addr_positional[14355:14352], addr_3588_6);

wire[27:0] addr_3589_6;

Selector_2 s3589_6(wires_897_5[1], addr_897_5, addr_positional[14359:14356], addr_3589_6);

wire[27:0] addr_3590_6;

Selector_2 s3590_6(wires_897_5[2], addr_897_5, addr_positional[14363:14360], addr_3590_6);

wire[27:0] addr_3591_6;

Selector_2 s3591_6(wires_897_5[3], addr_897_5, addr_positional[14367:14364], addr_3591_6);

wire[27:0] addr_3592_6;

Selector_2 s3592_6(wires_898_5[0], addr_898_5, addr_positional[14371:14368], addr_3592_6);

wire[27:0] addr_3593_6;

Selector_2 s3593_6(wires_898_5[1], addr_898_5, addr_positional[14375:14372], addr_3593_6);

wire[27:0] addr_3594_6;

Selector_2 s3594_6(wires_898_5[2], addr_898_5, addr_positional[14379:14376], addr_3594_6);

wire[27:0] addr_3595_6;

Selector_2 s3595_6(wires_898_5[3], addr_898_5, addr_positional[14383:14380], addr_3595_6);

wire[27:0] addr_3596_6;

Selector_2 s3596_6(wires_899_5[0], addr_899_5, addr_positional[14387:14384], addr_3596_6);

wire[27:0] addr_3597_6;

Selector_2 s3597_6(wires_899_5[1], addr_899_5, addr_positional[14391:14388], addr_3597_6);

wire[27:0] addr_3598_6;

Selector_2 s3598_6(wires_899_5[2], addr_899_5, addr_positional[14395:14392], addr_3598_6);

wire[27:0] addr_3599_6;

Selector_2 s3599_6(wires_899_5[3], addr_899_5, addr_positional[14399:14396], addr_3599_6);

wire[27:0] addr_3600_6;

Selector_2 s3600_6(wires_900_5[0], addr_900_5, addr_positional[14403:14400], addr_3600_6);

wire[27:0] addr_3601_6;

Selector_2 s3601_6(wires_900_5[1], addr_900_5, addr_positional[14407:14404], addr_3601_6);

wire[27:0] addr_3602_6;

Selector_2 s3602_6(wires_900_5[2], addr_900_5, addr_positional[14411:14408], addr_3602_6);

wire[27:0] addr_3603_6;

Selector_2 s3603_6(wires_900_5[3], addr_900_5, addr_positional[14415:14412], addr_3603_6);

wire[27:0] addr_3604_6;

Selector_2 s3604_6(wires_901_5[0], addr_901_5, addr_positional[14419:14416], addr_3604_6);

wire[27:0] addr_3605_6;

Selector_2 s3605_6(wires_901_5[1], addr_901_5, addr_positional[14423:14420], addr_3605_6);

wire[27:0] addr_3606_6;

Selector_2 s3606_6(wires_901_5[2], addr_901_5, addr_positional[14427:14424], addr_3606_6);

wire[27:0] addr_3607_6;

Selector_2 s3607_6(wires_901_5[3], addr_901_5, addr_positional[14431:14428], addr_3607_6);

wire[27:0] addr_3608_6;

Selector_2 s3608_6(wires_902_5[0], addr_902_5, addr_positional[14435:14432], addr_3608_6);

wire[27:0] addr_3609_6;

Selector_2 s3609_6(wires_902_5[1], addr_902_5, addr_positional[14439:14436], addr_3609_6);

wire[27:0] addr_3610_6;

Selector_2 s3610_6(wires_902_5[2], addr_902_5, addr_positional[14443:14440], addr_3610_6);

wire[27:0] addr_3611_6;

Selector_2 s3611_6(wires_902_5[3], addr_902_5, addr_positional[14447:14444], addr_3611_6);

wire[27:0] addr_3612_6;

Selector_2 s3612_6(wires_903_5[0], addr_903_5, addr_positional[14451:14448], addr_3612_6);

wire[27:0] addr_3613_6;

Selector_2 s3613_6(wires_903_5[1], addr_903_5, addr_positional[14455:14452], addr_3613_6);

wire[27:0] addr_3614_6;

Selector_2 s3614_6(wires_903_5[2], addr_903_5, addr_positional[14459:14456], addr_3614_6);

wire[27:0] addr_3615_6;

Selector_2 s3615_6(wires_903_5[3], addr_903_5, addr_positional[14463:14460], addr_3615_6);

wire[27:0] addr_3616_6;

Selector_2 s3616_6(wires_904_5[0], addr_904_5, addr_positional[14467:14464], addr_3616_6);

wire[27:0] addr_3617_6;

Selector_2 s3617_6(wires_904_5[1], addr_904_5, addr_positional[14471:14468], addr_3617_6);

wire[27:0] addr_3618_6;

Selector_2 s3618_6(wires_904_5[2], addr_904_5, addr_positional[14475:14472], addr_3618_6);

wire[27:0] addr_3619_6;

Selector_2 s3619_6(wires_904_5[3], addr_904_5, addr_positional[14479:14476], addr_3619_6);

wire[27:0] addr_3620_6;

Selector_2 s3620_6(wires_905_5[0], addr_905_5, addr_positional[14483:14480], addr_3620_6);

wire[27:0] addr_3621_6;

Selector_2 s3621_6(wires_905_5[1], addr_905_5, addr_positional[14487:14484], addr_3621_6);

wire[27:0] addr_3622_6;

Selector_2 s3622_6(wires_905_5[2], addr_905_5, addr_positional[14491:14488], addr_3622_6);

wire[27:0] addr_3623_6;

Selector_2 s3623_6(wires_905_5[3], addr_905_5, addr_positional[14495:14492], addr_3623_6);

wire[27:0] addr_3624_6;

Selector_2 s3624_6(wires_906_5[0], addr_906_5, addr_positional[14499:14496], addr_3624_6);

wire[27:0] addr_3625_6;

Selector_2 s3625_6(wires_906_5[1], addr_906_5, addr_positional[14503:14500], addr_3625_6);

wire[27:0] addr_3626_6;

Selector_2 s3626_6(wires_906_5[2], addr_906_5, addr_positional[14507:14504], addr_3626_6);

wire[27:0] addr_3627_6;

Selector_2 s3627_6(wires_906_5[3], addr_906_5, addr_positional[14511:14508], addr_3627_6);

wire[27:0] addr_3628_6;

Selector_2 s3628_6(wires_907_5[0], addr_907_5, addr_positional[14515:14512], addr_3628_6);

wire[27:0] addr_3629_6;

Selector_2 s3629_6(wires_907_5[1], addr_907_5, addr_positional[14519:14516], addr_3629_6);

wire[27:0] addr_3630_6;

Selector_2 s3630_6(wires_907_5[2], addr_907_5, addr_positional[14523:14520], addr_3630_6);

wire[27:0] addr_3631_6;

Selector_2 s3631_6(wires_907_5[3], addr_907_5, addr_positional[14527:14524], addr_3631_6);

wire[27:0] addr_3632_6;

Selector_2 s3632_6(wires_908_5[0], addr_908_5, addr_positional[14531:14528], addr_3632_6);

wire[27:0] addr_3633_6;

Selector_2 s3633_6(wires_908_5[1], addr_908_5, addr_positional[14535:14532], addr_3633_6);

wire[27:0] addr_3634_6;

Selector_2 s3634_6(wires_908_5[2], addr_908_5, addr_positional[14539:14536], addr_3634_6);

wire[27:0] addr_3635_6;

Selector_2 s3635_6(wires_908_5[3], addr_908_5, addr_positional[14543:14540], addr_3635_6);

wire[27:0] addr_3636_6;

Selector_2 s3636_6(wires_909_5[0], addr_909_5, addr_positional[14547:14544], addr_3636_6);

wire[27:0] addr_3637_6;

Selector_2 s3637_6(wires_909_5[1], addr_909_5, addr_positional[14551:14548], addr_3637_6);

wire[27:0] addr_3638_6;

Selector_2 s3638_6(wires_909_5[2], addr_909_5, addr_positional[14555:14552], addr_3638_6);

wire[27:0] addr_3639_6;

Selector_2 s3639_6(wires_909_5[3], addr_909_5, addr_positional[14559:14556], addr_3639_6);

wire[27:0] addr_3640_6;

Selector_2 s3640_6(wires_910_5[0], addr_910_5, addr_positional[14563:14560], addr_3640_6);

wire[27:0] addr_3641_6;

Selector_2 s3641_6(wires_910_5[1], addr_910_5, addr_positional[14567:14564], addr_3641_6);

wire[27:0] addr_3642_6;

Selector_2 s3642_6(wires_910_5[2], addr_910_5, addr_positional[14571:14568], addr_3642_6);

wire[27:0] addr_3643_6;

Selector_2 s3643_6(wires_910_5[3], addr_910_5, addr_positional[14575:14572], addr_3643_6);

wire[27:0] addr_3644_6;

Selector_2 s3644_6(wires_911_5[0], addr_911_5, addr_positional[14579:14576], addr_3644_6);

wire[27:0] addr_3645_6;

Selector_2 s3645_6(wires_911_5[1], addr_911_5, addr_positional[14583:14580], addr_3645_6);

wire[27:0] addr_3646_6;

Selector_2 s3646_6(wires_911_5[2], addr_911_5, addr_positional[14587:14584], addr_3646_6);

wire[27:0] addr_3647_6;

Selector_2 s3647_6(wires_911_5[3], addr_911_5, addr_positional[14591:14588], addr_3647_6);

wire[27:0] addr_3648_6;

Selector_2 s3648_6(wires_912_5[0], addr_912_5, addr_positional[14595:14592], addr_3648_6);

wire[27:0] addr_3649_6;

Selector_2 s3649_6(wires_912_5[1], addr_912_5, addr_positional[14599:14596], addr_3649_6);

wire[27:0] addr_3650_6;

Selector_2 s3650_6(wires_912_5[2], addr_912_5, addr_positional[14603:14600], addr_3650_6);

wire[27:0] addr_3651_6;

Selector_2 s3651_6(wires_912_5[3], addr_912_5, addr_positional[14607:14604], addr_3651_6);

wire[27:0] addr_3652_6;

Selector_2 s3652_6(wires_913_5[0], addr_913_5, addr_positional[14611:14608], addr_3652_6);

wire[27:0] addr_3653_6;

Selector_2 s3653_6(wires_913_5[1], addr_913_5, addr_positional[14615:14612], addr_3653_6);

wire[27:0] addr_3654_6;

Selector_2 s3654_6(wires_913_5[2], addr_913_5, addr_positional[14619:14616], addr_3654_6);

wire[27:0] addr_3655_6;

Selector_2 s3655_6(wires_913_5[3], addr_913_5, addr_positional[14623:14620], addr_3655_6);

wire[27:0] addr_3656_6;

Selector_2 s3656_6(wires_914_5[0], addr_914_5, addr_positional[14627:14624], addr_3656_6);

wire[27:0] addr_3657_6;

Selector_2 s3657_6(wires_914_5[1], addr_914_5, addr_positional[14631:14628], addr_3657_6);

wire[27:0] addr_3658_6;

Selector_2 s3658_6(wires_914_5[2], addr_914_5, addr_positional[14635:14632], addr_3658_6);

wire[27:0] addr_3659_6;

Selector_2 s3659_6(wires_914_5[3], addr_914_5, addr_positional[14639:14636], addr_3659_6);

wire[27:0] addr_3660_6;

Selector_2 s3660_6(wires_915_5[0], addr_915_5, addr_positional[14643:14640], addr_3660_6);

wire[27:0] addr_3661_6;

Selector_2 s3661_6(wires_915_5[1], addr_915_5, addr_positional[14647:14644], addr_3661_6);

wire[27:0] addr_3662_6;

Selector_2 s3662_6(wires_915_5[2], addr_915_5, addr_positional[14651:14648], addr_3662_6);

wire[27:0] addr_3663_6;

Selector_2 s3663_6(wires_915_5[3], addr_915_5, addr_positional[14655:14652], addr_3663_6);

wire[27:0] addr_3664_6;

Selector_2 s3664_6(wires_916_5[0], addr_916_5, addr_positional[14659:14656], addr_3664_6);

wire[27:0] addr_3665_6;

Selector_2 s3665_6(wires_916_5[1], addr_916_5, addr_positional[14663:14660], addr_3665_6);

wire[27:0] addr_3666_6;

Selector_2 s3666_6(wires_916_5[2], addr_916_5, addr_positional[14667:14664], addr_3666_6);

wire[27:0] addr_3667_6;

Selector_2 s3667_6(wires_916_5[3], addr_916_5, addr_positional[14671:14668], addr_3667_6);

wire[27:0] addr_3668_6;

Selector_2 s3668_6(wires_917_5[0], addr_917_5, addr_positional[14675:14672], addr_3668_6);

wire[27:0] addr_3669_6;

Selector_2 s3669_6(wires_917_5[1], addr_917_5, addr_positional[14679:14676], addr_3669_6);

wire[27:0] addr_3670_6;

Selector_2 s3670_6(wires_917_5[2], addr_917_5, addr_positional[14683:14680], addr_3670_6);

wire[27:0] addr_3671_6;

Selector_2 s3671_6(wires_917_5[3], addr_917_5, addr_positional[14687:14684], addr_3671_6);

wire[27:0] addr_3672_6;

Selector_2 s3672_6(wires_918_5[0], addr_918_5, addr_positional[14691:14688], addr_3672_6);

wire[27:0] addr_3673_6;

Selector_2 s3673_6(wires_918_5[1], addr_918_5, addr_positional[14695:14692], addr_3673_6);

wire[27:0] addr_3674_6;

Selector_2 s3674_6(wires_918_5[2], addr_918_5, addr_positional[14699:14696], addr_3674_6);

wire[27:0] addr_3675_6;

Selector_2 s3675_6(wires_918_5[3], addr_918_5, addr_positional[14703:14700], addr_3675_6);

wire[27:0] addr_3676_6;

Selector_2 s3676_6(wires_919_5[0], addr_919_5, addr_positional[14707:14704], addr_3676_6);

wire[27:0] addr_3677_6;

Selector_2 s3677_6(wires_919_5[1], addr_919_5, addr_positional[14711:14708], addr_3677_6);

wire[27:0] addr_3678_6;

Selector_2 s3678_6(wires_919_5[2], addr_919_5, addr_positional[14715:14712], addr_3678_6);

wire[27:0] addr_3679_6;

Selector_2 s3679_6(wires_919_5[3], addr_919_5, addr_positional[14719:14716], addr_3679_6);

wire[27:0] addr_3680_6;

Selector_2 s3680_6(wires_920_5[0], addr_920_5, addr_positional[14723:14720], addr_3680_6);

wire[27:0] addr_3681_6;

Selector_2 s3681_6(wires_920_5[1], addr_920_5, addr_positional[14727:14724], addr_3681_6);

wire[27:0] addr_3682_6;

Selector_2 s3682_6(wires_920_5[2], addr_920_5, addr_positional[14731:14728], addr_3682_6);

wire[27:0] addr_3683_6;

Selector_2 s3683_6(wires_920_5[3], addr_920_5, addr_positional[14735:14732], addr_3683_6);

wire[27:0] addr_3684_6;

Selector_2 s3684_6(wires_921_5[0], addr_921_5, addr_positional[14739:14736], addr_3684_6);

wire[27:0] addr_3685_6;

Selector_2 s3685_6(wires_921_5[1], addr_921_5, addr_positional[14743:14740], addr_3685_6);

wire[27:0] addr_3686_6;

Selector_2 s3686_6(wires_921_5[2], addr_921_5, addr_positional[14747:14744], addr_3686_6);

wire[27:0] addr_3687_6;

Selector_2 s3687_6(wires_921_5[3], addr_921_5, addr_positional[14751:14748], addr_3687_6);

wire[27:0] addr_3688_6;

Selector_2 s3688_6(wires_922_5[0], addr_922_5, addr_positional[14755:14752], addr_3688_6);

wire[27:0] addr_3689_6;

Selector_2 s3689_6(wires_922_5[1], addr_922_5, addr_positional[14759:14756], addr_3689_6);

wire[27:0] addr_3690_6;

Selector_2 s3690_6(wires_922_5[2], addr_922_5, addr_positional[14763:14760], addr_3690_6);

wire[27:0] addr_3691_6;

Selector_2 s3691_6(wires_922_5[3], addr_922_5, addr_positional[14767:14764], addr_3691_6);

wire[27:0] addr_3692_6;

Selector_2 s3692_6(wires_923_5[0], addr_923_5, addr_positional[14771:14768], addr_3692_6);

wire[27:0] addr_3693_6;

Selector_2 s3693_6(wires_923_5[1], addr_923_5, addr_positional[14775:14772], addr_3693_6);

wire[27:0] addr_3694_6;

Selector_2 s3694_6(wires_923_5[2], addr_923_5, addr_positional[14779:14776], addr_3694_6);

wire[27:0] addr_3695_6;

Selector_2 s3695_6(wires_923_5[3], addr_923_5, addr_positional[14783:14780], addr_3695_6);

wire[27:0] addr_3696_6;

Selector_2 s3696_6(wires_924_5[0], addr_924_5, addr_positional[14787:14784], addr_3696_6);

wire[27:0] addr_3697_6;

Selector_2 s3697_6(wires_924_5[1], addr_924_5, addr_positional[14791:14788], addr_3697_6);

wire[27:0] addr_3698_6;

Selector_2 s3698_6(wires_924_5[2], addr_924_5, addr_positional[14795:14792], addr_3698_6);

wire[27:0] addr_3699_6;

Selector_2 s3699_6(wires_924_5[3], addr_924_5, addr_positional[14799:14796], addr_3699_6);

wire[27:0] addr_3700_6;

Selector_2 s3700_6(wires_925_5[0], addr_925_5, addr_positional[14803:14800], addr_3700_6);

wire[27:0] addr_3701_6;

Selector_2 s3701_6(wires_925_5[1], addr_925_5, addr_positional[14807:14804], addr_3701_6);

wire[27:0] addr_3702_6;

Selector_2 s3702_6(wires_925_5[2], addr_925_5, addr_positional[14811:14808], addr_3702_6);

wire[27:0] addr_3703_6;

Selector_2 s3703_6(wires_925_5[3], addr_925_5, addr_positional[14815:14812], addr_3703_6);

wire[27:0] addr_3704_6;

Selector_2 s3704_6(wires_926_5[0], addr_926_5, addr_positional[14819:14816], addr_3704_6);

wire[27:0] addr_3705_6;

Selector_2 s3705_6(wires_926_5[1], addr_926_5, addr_positional[14823:14820], addr_3705_6);

wire[27:0] addr_3706_6;

Selector_2 s3706_6(wires_926_5[2], addr_926_5, addr_positional[14827:14824], addr_3706_6);

wire[27:0] addr_3707_6;

Selector_2 s3707_6(wires_926_5[3], addr_926_5, addr_positional[14831:14828], addr_3707_6);

wire[27:0] addr_3708_6;

Selector_2 s3708_6(wires_927_5[0], addr_927_5, addr_positional[14835:14832], addr_3708_6);

wire[27:0] addr_3709_6;

Selector_2 s3709_6(wires_927_5[1], addr_927_5, addr_positional[14839:14836], addr_3709_6);

wire[27:0] addr_3710_6;

Selector_2 s3710_6(wires_927_5[2], addr_927_5, addr_positional[14843:14840], addr_3710_6);

wire[27:0] addr_3711_6;

Selector_2 s3711_6(wires_927_5[3], addr_927_5, addr_positional[14847:14844], addr_3711_6);

wire[27:0] addr_3712_6;

Selector_2 s3712_6(wires_928_5[0], addr_928_5, addr_positional[14851:14848], addr_3712_6);

wire[27:0] addr_3713_6;

Selector_2 s3713_6(wires_928_5[1], addr_928_5, addr_positional[14855:14852], addr_3713_6);

wire[27:0] addr_3714_6;

Selector_2 s3714_6(wires_928_5[2], addr_928_5, addr_positional[14859:14856], addr_3714_6);

wire[27:0] addr_3715_6;

Selector_2 s3715_6(wires_928_5[3], addr_928_5, addr_positional[14863:14860], addr_3715_6);

wire[27:0] addr_3716_6;

Selector_2 s3716_6(wires_929_5[0], addr_929_5, addr_positional[14867:14864], addr_3716_6);

wire[27:0] addr_3717_6;

Selector_2 s3717_6(wires_929_5[1], addr_929_5, addr_positional[14871:14868], addr_3717_6);

wire[27:0] addr_3718_6;

Selector_2 s3718_6(wires_929_5[2], addr_929_5, addr_positional[14875:14872], addr_3718_6);

wire[27:0] addr_3719_6;

Selector_2 s3719_6(wires_929_5[3], addr_929_5, addr_positional[14879:14876], addr_3719_6);

wire[27:0] addr_3720_6;

Selector_2 s3720_6(wires_930_5[0], addr_930_5, addr_positional[14883:14880], addr_3720_6);

wire[27:0] addr_3721_6;

Selector_2 s3721_6(wires_930_5[1], addr_930_5, addr_positional[14887:14884], addr_3721_6);

wire[27:0] addr_3722_6;

Selector_2 s3722_6(wires_930_5[2], addr_930_5, addr_positional[14891:14888], addr_3722_6);

wire[27:0] addr_3723_6;

Selector_2 s3723_6(wires_930_5[3], addr_930_5, addr_positional[14895:14892], addr_3723_6);

wire[27:0] addr_3724_6;

Selector_2 s3724_6(wires_931_5[0], addr_931_5, addr_positional[14899:14896], addr_3724_6);

wire[27:0] addr_3725_6;

Selector_2 s3725_6(wires_931_5[1], addr_931_5, addr_positional[14903:14900], addr_3725_6);

wire[27:0] addr_3726_6;

Selector_2 s3726_6(wires_931_5[2], addr_931_5, addr_positional[14907:14904], addr_3726_6);

wire[27:0] addr_3727_6;

Selector_2 s3727_6(wires_931_5[3], addr_931_5, addr_positional[14911:14908], addr_3727_6);

wire[27:0] addr_3728_6;

Selector_2 s3728_6(wires_932_5[0], addr_932_5, addr_positional[14915:14912], addr_3728_6);

wire[27:0] addr_3729_6;

Selector_2 s3729_6(wires_932_5[1], addr_932_5, addr_positional[14919:14916], addr_3729_6);

wire[27:0] addr_3730_6;

Selector_2 s3730_6(wires_932_5[2], addr_932_5, addr_positional[14923:14920], addr_3730_6);

wire[27:0] addr_3731_6;

Selector_2 s3731_6(wires_932_5[3], addr_932_5, addr_positional[14927:14924], addr_3731_6);

wire[27:0] addr_3732_6;

Selector_2 s3732_6(wires_933_5[0], addr_933_5, addr_positional[14931:14928], addr_3732_6);

wire[27:0] addr_3733_6;

Selector_2 s3733_6(wires_933_5[1], addr_933_5, addr_positional[14935:14932], addr_3733_6);

wire[27:0] addr_3734_6;

Selector_2 s3734_6(wires_933_5[2], addr_933_5, addr_positional[14939:14936], addr_3734_6);

wire[27:0] addr_3735_6;

Selector_2 s3735_6(wires_933_5[3], addr_933_5, addr_positional[14943:14940], addr_3735_6);

wire[27:0] addr_3736_6;

Selector_2 s3736_6(wires_934_5[0], addr_934_5, addr_positional[14947:14944], addr_3736_6);

wire[27:0] addr_3737_6;

Selector_2 s3737_6(wires_934_5[1], addr_934_5, addr_positional[14951:14948], addr_3737_6);

wire[27:0] addr_3738_6;

Selector_2 s3738_6(wires_934_5[2], addr_934_5, addr_positional[14955:14952], addr_3738_6);

wire[27:0] addr_3739_6;

Selector_2 s3739_6(wires_934_5[3], addr_934_5, addr_positional[14959:14956], addr_3739_6);

wire[27:0] addr_3740_6;

Selector_2 s3740_6(wires_935_5[0], addr_935_5, addr_positional[14963:14960], addr_3740_6);

wire[27:0] addr_3741_6;

Selector_2 s3741_6(wires_935_5[1], addr_935_5, addr_positional[14967:14964], addr_3741_6);

wire[27:0] addr_3742_6;

Selector_2 s3742_6(wires_935_5[2], addr_935_5, addr_positional[14971:14968], addr_3742_6);

wire[27:0] addr_3743_6;

Selector_2 s3743_6(wires_935_5[3], addr_935_5, addr_positional[14975:14972], addr_3743_6);

wire[27:0] addr_3744_6;

Selector_2 s3744_6(wires_936_5[0], addr_936_5, addr_positional[14979:14976], addr_3744_6);

wire[27:0] addr_3745_6;

Selector_2 s3745_6(wires_936_5[1], addr_936_5, addr_positional[14983:14980], addr_3745_6);

wire[27:0] addr_3746_6;

Selector_2 s3746_6(wires_936_5[2], addr_936_5, addr_positional[14987:14984], addr_3746_6);

wire[27:0] addr_3747_6;

Selector_2 s3747_6(wires_936_5[3], addr_936_5, addr_positional[14991:14988], addr_3747_6);

wire[27:0] addr_3748_6;

Selector_2 s3748_6(wires_937_5[0], addr_937_5, addr_positional[14995:14992], addr_3748_6);

wire[27:0] addr_3749_6;

Selector_2 s3749_6(wires_937_5[1], addr_937_5, addr_positional[14999:14996], addr_3749_6);

wire[27:0] addr_3750_6;

Selector_2 s3750_6(wires_937_5[2], addr_937_5, addr_positional[15003:15000], addr_3750_6);

wire[27:0] addr_3751_6;

Selector_2 s3751_6(wires_937_5[3], addr_937_5, addr_positional[15007:15004], addr_3751_6);

wire[27:0] addr_3752_6;

Selector_2 s3752_6(wires_938_5[0], addr_938_5, addr_positional[15011:15008], addr_3752_6);

wire[27:0] addr_3753_6;

Selector_2 s3753_6(wires_938_5[1], addr_938_5, addr_positional[15015:15012], addr_3753_6);

wire[27:0] addr_3754_6;

Selector_2 s3754_6(wires_938_5[2], addr_938_5, addr_positional[15019:15016], addr_3754_6);

wire[27:0] addr_3755_6;

Selector_2 s3755_6(wires_938_5[3], addr_938_5, addr_positional[15023:15020], addr_3755_6);

wire[27:0] addr_3756_6;

Selector_2 s3756_6(wires_939_5[0], addr_939_5, addr_positional[15027:15024], addr_3756_6);

wire[27:0] addr_3757_6;

Selector_2 s3757_6(wires_939_5[1], addr_939_5, addr_positional[15031:15028], addr_3757_6);

wire[27:0] addr_3758_6;

Selector_2 s3758_6(wires_939_5[2], addr_939_5, addr_positional[15035:15032], addr_3758_6);

wire[27:0] addr_3759_6;

Selector_2 s3759_6(wires_939_5[3], addr_939_5, addr_positional[15039:15036], addr_3759_6);

wire[27:0] addr_3760_6;

Selector_2 s3760_6(wires_940_5[0], addr_940_5, addr_positional[15043:15040], addr_3760_6);

wire[27:0] addr_3761_6;

Selector_2 s3761_6(wires_940_5[1], addr_940_5, addr_positional[15047:15044], addr_3761_6);

wire[27:0] addr_3762_6;

Selector_2 s3762_6(wires_940_5[2], addr_940_5, addr_positional[15051:15048], addr_3762_6);

wire[27:0] addr_3763_6;

Selector_2 s3763_6(wires_940_5[3], addr_940_5, addr_positional[15055:15052], addr_3763_6);

wire[27:0] addr_3764_6;

Selector_2 s3764_6(wires_941_5[0], addr_941_5, addr_positional[15059:15056], addr_3764_6);

wire[27:0] addr_3765_6;

Selector_2 s3765_6(wires_941_5[1], addr_941_5, addr_positional[15063:15060], addr_3765_6);

wire[27:0] addr_3766_6;

Selector_2 s3766_6(wires_941_5[2], addr_941_5, addr_positional[15067:15064], addr_3766_6);

wire[27:0] addr_3767_6;

Selector_2 s3767_6(wires_941_5[3], addr_941_5, addr_positional[15071:15068], addr_3767_6);

wire[27:0] addr_3768_6;

Selector_2 s3768_6(wires_942_5[0], addr_942_5, addr_positional[15075:15072], addr_3768_6);

wire[27:0] addr_3769_6;

Selector_2 s3769_6(wires_942_5[1], addr_942_5, addr_positional[15079:15076], addr_3769_6);

wire[27:0] addr_3770_6;

Selector_2 s3770_6(wires_942_5[2], addr_942_5, addr_positional[15083:15080], addr_3770_6);

wire[27:0] addr_3771_6;

Selector_2 s3771_6(wires_942_5[3], addr_942_5, addr_positional[15087:15084], addr_3771_6);

wire[27:0] addr_3772_6;

Selector_2 s3772_6(wires_943_5[0], addr_943_5, addr_positional[15091:15088], addr_3772_6);

wire[27:0] addr_3773_6;

Selector_2 s3773_6(wires_943_5[1], addr_943_5, addr_positional[15095:15092], addr_3773_6);

wire[27:0] addr_3774_6;

Selector_2 s3774_6(wires_943_5[2], addr_943_5, addr_positional[15099:15096], addr_3774_6);

wire[27:0] addr_3775_6;

Selector_2 s3775_6(wires_943_5[3], addr_943_5, addr_positional[15103:15100], addr_3775_6);

wire[27:0] addr_3776_6;

Selector_2 s3776_6(wires_944_5[0], addr_944_5, addr_positional[15107:15104], addr_3776_6);

wire[27:0] addr_3777_6;

Selector_2 s3777_6(wires_944_5[1], addr_944_5, addr_positional[15111:15108], addr_3777_6);

wire[27:0] addr_3778_6;

Selector_2 s3778_6(wires_944_5[2], addr_944_5, addr_positional[15115:15112], addr_3778_6);

wire[27:0] addr_3779_6;

Selector_2 s3779_6(wires_944_5[3], addr_944_5, addr_positional[15119:15116], addr_3779_6);

wire[27:0] addr_3780_6;

Selector_2 s3780_6(wires_945_5[0], addr_945_5, addr_positional[15123:15120], addr_3780_6);

wire[27:0] addr_3781_6;

Selector_2 s3781_6(wires_945_5[1], addr_945_5, addr_positional[15127:15124], addr_3781_6);

wire[27:0] addr_3782_6;

Selector_2 s3782_6(wires_945_5[2], addr_945_5, addr_positional[15131:15128], addr_3782_6);

wire[27:0] addr_3783_6;

Selector_2 s3783_6(wires_945_5[3], addr_945_5, addr_positional[15135:15132], addr_3783_6);

wire[27:0] addr_3784_6;

Selector_2 s3784_6(wires_946_5[0], addr_946_5, addr_positional[15139:15136], addr_3784_6);

wire[27:0] addr_3785_6;

Selector_2 s3785_6(wires_946_5[1], addr_946_5, addr_positional[15143:15140], addr_3785_6);

wire[27:0] addr_3786_6;

Selector_2 s3786_6(wires_946_5[2], addr_946_5, addr_positional[15147:15144], addr_3786_6);

wire[27:0] addr_3787_6;

Selector_2 s3787_6(wires_946_5[3], addr_946_5, addr_positional[15151:15148], addr_3787_6);

wire[27:0] addr_3788_6;

Selector_2 s3788_6(wires_947_5[0], addr_947_5, addr_positional[15155:15152], addr_3788_6);

wire[27:0] addr_3789_6;

Selector_2 s3789_6(wires_947_5[1], addr_947_5, addr_positional[15159:15156], addr_3789_6);

wire[27:0] addr_3790_6;

Selector_2 s3790_6(wires_947_5[2], addr_947_5, addr_positional[15163:15160], addr_3790_6);

wire[27:0] addr_3791_6;

Selector_2 s3791_6(wires_947_5[3], addr_947_5, addr_positional[15167:15164], addr_3791_6);

wire[27:0] addr_3792_6;

Selector_2 s3792_6(wires_948_5[0], addr_948_5, addr_positional[15171:15168], addr_3792_6);

wire[27:0] addr_3793_6;

Selector_2 s3793_6(wires_948_5[1], addr_948_5, addr_positional[15175:15172], addr_3793_6);

wire[27:0] addr_3794_6;

Selector_2 s3794_6(wires_948_5[2], addr_948_5, addr_positional[15179:15176], addr_3794_6);

wire[27:0] addr_3795_6;

Selector_2 s3795_6(wires_948_5[3], addr_948_5, addr_positional[15183:15180], addr_3795_6);

wire[27:0] addr_3796_6;

Selector_2 s3796_6(wires_949_5[0], addr_949_5, addr_positional[15187:15184], addr_3796_6);

wire[27:0] addr_3797_6;

Selector_2 s3797_6(wires_949_5[1], addr_949_5, addr_positional[15191:15188], addr_3797_6);

wire[27:0] addr_3798_6;

Selector_2 s3798_6(wires_949_5[2], addr_949_5, addr_positional[15195:15192], addr_3798_6);

wire[27:0] addr_3799_6;

Selector_2 s3799_6(wires_949_5[3], addr_949_5, addr_positional[15199:15196], addr_3799_6);

wire[27:0] addr_3800_6;

Selector_2 s3800_6(wires_950_5[0], addr_950_5, addr_positional[15203:15200], addr_3800_6);

wire[27:0] addr_3801_6;

Selector_2 s3801_6(wires_950_5[1], addr_950_5, addr_positional[15207:15204], addr_3801_6);

wire[27:0] addr_3802_6;

Selector_2 s3802_6(wires_950_5[2], addr_950_5, addr_positional[15211:15208], addr_3802_6);

wire[27:0] addr_3803_6;

Selector_2 s3803_6(wires_950_5[3], addr_950_5, addr_positional[15215:15212], addr_3803_6);

wire[27:0] addr_3804_6;

Selector_2 s3804_6(wires_951_5[0], addr_951_5, addr_positional[15219:15216], addr_3804_6);

wire[27:0] addr_3805_6;

Selector_2 s3805_6(wires_951_5[1], addr_951_5, addr_positional[15223:15220], addr_3805_6);

wire[27:0] addr_3806_6;

Selector_2 s3806_6(wires_951_5[2], addr_951_5, addr_positional[15227:15224], addr_3806_6);

wire[27:0] addr_3807_6;

Selector_2 s3807_6(wires_951_5[3], addr_951_5, addr_positional[15231:15228], addr_3807_6);

wire[27:0] addr_3808_6;

Selector_2 s3808_6(wires_952_5[0], addr_952_5, addr_positional[15235:15232], addr_3808_6);

wire[27:0] addr_3809_6;

Selector_2 s3809_6(wires_952_5[1], addr_952_5, addr_positional[15239:15236], addr_3809_6);

wire[27:0] addr_3810_6;

Selector_2 s3810_6(wires_952_5[2], addr_952_5, addr_positional[15243:15240], addr_3810_6);

wire[27:0] addr_3811_6;

Selector_2 s3811_6(wires_952_5[3], addr_952_5, addr_positional[15247:15244], addr_3811_6);

wire[27:0] addr_3812_6;

Selector_2 s3812_6(wires_953_5[0], addr_953_5, addr_positional[15251:15248], addr_3812_6);

wire[27:0] addr_3813_6;

Selector_2 s3813_6(wires_953_5[1], addr_953_5, addr_positional[15255:15252], addr_3813_6);

wire[27:0] addr_3814_6;

Selector_2 s3814_6(wires_953_5[2], addr_953_5, addr_positional[15259:15256], addr_3814_6);

wire[27:0] addr_3815_6;

Selector_2 s3815_6(wires_953_5[3], addr_953_5, addr_positional[15263:15260], addr_3815_6);

wire[27:0] addr_3816_6;

Selector_2 s3816_6(wires_954_5[0], addr_954_5, addr_positional[15267:15264], addr_3816_6);

wire[27:0] addr_3817_6;

Selector_2 s3817_6(wires_954_5[1], addr_954_5, addr_positional[15271:15268], addr_3817_6);

wire[27:0] addr_3818_6;

Selector_2 s3818_6(wires_954_5[2], addr_954_5, addr_positional[15275:15272], addr_3818_6);

wire[27:0] addr_3819_6;

Selector_2 s3819_6(wires_954_5[3], addr_954_5, addr_positional[15279:15276], addr_3819_6);

wire[27:0] addr_3820_6;

Selector_2 s3820_6(wires_955_5[0], addr_955_5, addr_positional[15283:15280], addr_3820_6);

wire[27:0] addr_3821_6;

Selector_2 s3821_6(wires_955_5[1], addr_955_5, addr_positional[15287:15284], addr_3821_6);

wire[27:0] addr_3822_6;

Selector_2 s3822_6(wires_955_5[2], addr_955_5, addr_positional[15291:15288], addr_3822_6);

wire[27:0] addr_3823_6;

Selector_2 s3823_6(wires_955_5[3], addr_955_5, addr_positional[15295:15292], addr_3823_6);

wire[27:0] addr_3824_6;

Selector_2 s3824_6(wires_956_5[0], addr_956_5, addr_positional[15299:15296], addr_3824_6);

wire[27:0] addr_3825_6;

Selector_2 s3825_6(wires_956_5[1], addr_956_5, addr_positional[15303:15300], addr_3825_6);

wire[27:0] addr_3826_6;

Selector_2 s3826_6(wires_956_5[2], addr_956_5, addr_positional[15307:15304], addr_3826_6);

wire[27:0] addr_3827_6;

Selector_2 s3827_6(wires_956_5[3], addr_956_5, addr_positional[15311:15308], addr_3827_6);

wire[27:0] addr_3828_6;

Selector_2 s3828_6(wires_957_5[0], addr_957_5, addr_positional[15315:15312], addr_3828_6);

wire[27:0] addr_3829_6;

Selector_2 s3829_6(wires_957_5[1], addr_957_5, addr_positional[15319:15316], addr_3829_6);

wire[27:0] addr_3830_6;

Selector_2 s3830_6(wires_957_5[2], addr_957_5, addr_positional[15323:15320], addr_3830_6);

wire[27:0] addr_3831_6;

Selector_2 s3831_6(wires_957_5[3], addr_957_5, addr_positional[15327:15324], addr_3831_6);

wire[27:0] addr_3832_6;

Selector_2 s3832_6(wires_958_5[0], addr_958_5, addr_positional[15331:15328], addr_3832_6);

wire[27:0] addr_3833_6;

Selector_2 s3833_6(wires_958_5[1], addr_958_5, addr_positional[15335:15332], addr_3833_6);

wire[27:0] addr_3834_6;

Selector_2 s3834_6(wires_958_5[2], addr_958_5, addr_positional[15339:15336], addr_3834_6);

wire[27:0] addr_3835_6;

Selector_2 s3835_6(wires_958_5[3], addr_958_5, addr_positional[15343:15340], addr_3835_6);

wire[27:0] addr_3836_6;

Selector_2 s3836_6(wires_959_5[0], addr_959_5, addr_positional[15347:15344], addr_3836_6);

wire[27:0] addr_3837_6;

Selector_2 s3837_6(wires_959_5[1], addr_959_5, addr_positional[15351:15348], addr_3837_6);

wire[27:0] addr_3838_6;

Selector_2 s3838_6(wires_959_5[2], addr_959_5, addr_positional[15355:15352], addr_3838_6);

wire[27:0] addr_3839_6;

Selector_2 s3839_6(wires_959_5[3], addr_959_5, addr_positional[15359:15356], addr_3839_6);

wire[27:0] addr_3840_6;

Selector_2 s3840_6(wires_960_5[0], addr_960_5, addr_positional[15363:15360], addr_3840_6);

wire[27:0] addr_3841_6;

Selector_2 s3841_6(wires_960_5[1], addr_960_5, addr_positional[15367:15364], addr_3841_6);

wire[27:0] addr_3842_6;

Selector_2 s3842_6(wires_960_5[2], addr_960_5, addr_positional[15371:15368], addr_3842_6);

wire[27:0] addr_3843_6;

Selector_2 s3843_6(wires_960_5[3], addr_960_5, addr_positional[15375:15372], addr_3843_6);

wire[27:0] addr_3844_6;

Selector_2 s3844_6(wires_961_5[0], addr_961_5, addr_positional[15379:15376], addr_3844_6);

wire[27:0] addr_3845_6;

Selector_2 s3845_6(wires_961_5[1], addr_961_5, addr_positional[15383:15380], addr_3845_6);

wire[27:0] addr_3846_6;

Selector_2 s3846_6(wires_961_5[2], addr_961_5, addr_positional[15387:15384], addr_3846_6);

wire[27:0] addr_3847_6;

Selector_2 s3847_6(wires_961_5[3], addr_961_5, addr_positional[15391:15388], addr_3847_6);

wire[27:0] addr_3848_6;

Selector_2 s3848_6(wires_962_5[0], addr_962_5, addr_positional[15395:15392], addr_3848_6);

wire[27:0] addr_3849_6;

Selector_2 s3849_6(wires_962_5[1], addr_962_5, addr_positional[15399:15396], addr_3849_6);

wire[27:0] addr_3850_6;

Selector_2 s3850_6(wires_962_5[2], addr_962_5, addr_positional[15403:15400], addr_3850_6);

wire[27:0] addr_3851_6;

Selector_2 s3851_6(wires_962_5[3], addr_962_5, addr_positional[15407:15404], addr_3851_6);

wire[27:0] addr_3852_6;

Selector_2 s3852_6(wires_963_5[0], addr_963_5, addr_positional[15411:15408], addr_3852_6);

wire[27:0] addr_3853_6;

Selector_2 s3853_6(wires_963_5[1], addr_963_5, addr_positional[15415:15412], addr_3853_6);

wire[27:0] addr_3854_6;

Selector_2 s3854_6(wires_963_5[2], addr_963_5, addr_positional[15419:15416], addr_3854_6);

wire[27:0] addr_3855_6;

Selector_2 s3855_6(wires_963_5[3], addr_963_5, addr_positional[15423:15420], addr_3855_6);

wire[27:0] addr_3856_6;

Selector_2 s3856_6(wires_964_5[0], addr_964_5, addr_positional[15427:15424], addr_3856_6);

wire[27:0] addr_3857_6;

Selector_2 s3857_6(wires_964_5[1], addr_964_5, addr_positional[15431:15428], addr_3857_6);

wire[27:0] addr_3858_6;

Selector_2 s3858_6(wires_964_5[2], addr_964_5, addr_positional[15435:15432], addr_3858_6);

wire[27:0] addr_3859_6;

Selector_2 s3859_6(wires_964_5[3], addr_964_5, addr_positional[15439:15436], addr_3859_6);

wire[27:0] addr_3860_6;

Selector_2 s3860_6(wires_965_5[0], addr_965_5, addr_positional[15443:15440], addr_3860_6);

wire[27:0] addr_3861_6;

Selector_2 s3861_6(wires_965_5[1], addr_965_5, addr_positional[15447:15444], addr_3861_6);

wire[27:0] addr_3862_6;

Selector_2 s3862_6(wires_965_5[2], addr_965_5, addr_positional[15451:15448], addr_3862_6);

wire[27:0] addr_3863_6;

Selector_2 s3863_6(wires_965_5[3], addr_965_5, addr_positional[15455:15452], addr_3863_6);

wire[27:0] addr_3864_6;

Selector_2 s3864_6(wires_966_5[0], addr_966_5, addr_positional[15459:15456], addr_3864_6);

wire[27:0] addr_3865_6;

Selector_2 s3865_6(wires_966_5[1], addr_966_5, addr_positional[15463:15460], addr_3865_6);

wire[27:0] addr_3866_6;

Selector_2 s3866_6(wires_966_5[2], addr_966_5, addr_positional[15467:15464], addr_3866_6);

wire[27:0] addr_3867_6;

Selector_2 s3867_6(wires_966_5[3], addr_966_5, addr_positional[15471:15468], addr_3867_6);

wire[27:0] addr_3868_6;

Selector_2 s3868_6(wires_967_5[0], addr_967_5, addr_positional[15475:15472], addr_3868_6);

wire[27:0] addr_3869_6;

Selector_2 s3869_6(wires_967_5[1], addr_967_5, addr_positional[15479:15476], addr_3869_6);

wire[27:0] addr_3870_6;

Selector_2 s3870_6(wires_967_5[2], addr_967_5, addr_positional[15483:15480], addr_3870_6);

wire[27:0] addr_3871_6;

Selector_2 s3871_6(wires_967_5[3], addr_967_5, addr_positional[15487:15484], addr_3871_6);

wire[27:0] addr_3872_6;

Selector_2 s3872_6(wires_968_5[0], addr_968_5, addr_positional[15491:15488], addr_3872_6);

wire[27:0] addr_3873_6;

Selector_2 s3873_6(wires_968_5[1], addr_968_5, addr_positional[15495:15492], addr_3873_6);

wire[27:0] addr_3874_6;

Selector_2 s3874_6(wires_968_5[2], addr_968_5, addr_positional[15499:15496], addr_3874_6);

wire[27:0] addr_3875_6;

Selector_2 s3875_6(wires_968_5[3], addr_968_5, addr_positional[15503:15500], addr_3875_6);

wire[27:0] addr_3876_6;

Selector_2 s3876_6(wires_969_5[0], addr_969_5, addr_positional[15507:15504], addr_3876_6);

wire[27:0] addr_3877_6;

Selector_2 s3877_6(wires_969_5[1], addr_969_5, addr_positional[15511:15508], addr_3877_6);

wire[27:0] addr_3878_6;

Selector_2 s3878_6(wires_969_5[2], addr_969_5, addr_positional[15515:15512], addr_3878_6);

wire[27:0] addr_3879_6;

Selector_2 s3879_6(wires_969_5[3], addr_969_5, addr_positional[15519:15516], addr_3879_6);

wire[27:0] addr_3880_6;

Selector_2 s3880_6(wires_970_5[0], addr_970_5, addr_positional[15523:15520], addr_3880_6);

wire[27:0] addr_3881_6;

Selector_2 s3881_6(wires_970_5[1], addr_970_5, addr_positional[15527:15524], addr_3881_6);

wire[27:0] addr_3882_6;

Selector_2 s3882_6(wires_970_5[2], addr_970_5, addr_positional[15531:15528], addr_3882_6);

wire[27:0] addr_3883_6;

Selector_2 s3883_6(wires_970_5[3], addr_970_5, addr_positional[15535:15532], addr_3883_6);

wire[27:0] addr_3884_6;

Selector_2 s3884_6(wires_971_5[0], addr_971_5, addr_positional[15539:15536], addr_3884_6);

wire[27:0] addr_3885_6;

Selector_2 s3885_6(wires_971_5[1], addr_971_5, addr_positional[15543:15540], addr_3885_6);

wire[27:0] addr_3886_6;

Selector_2 s3886_6(wires_971_5[2], addr_971_5, addr_positional[15547:15544], addr_3886_6);

wire[27:0] addr_3887_6;

Selector_2 s3887_6(wires_971_5[3], addr_971_5, addr_positional[15551:15548], addr_3887_6);

wire[27:0] addr_3888_6;

Selector_2 s3888_6(wires_972_5[0], addr_972_5, addr_positional[15555:15552], addr_3888_6);

wire[27:0] addr_3889_6;

Selector_2 s3889_6(wires_972_5[1], addr_972_5, addr_positional[15559:15556], addr_3889_6);

wire[27:0] addr_3890_6;

Selector_2 s3890_6(wires_972_5[2], addr_972_5, addr_positional[15563:15560], addr_3890_6);

wire[27:0] addr_3891_6;

Selector_2 s3891_6(wires_972_5[3], addr_972_5, addr_positional[15567:15564], addr_3891_6);

wire[27:0] addr_3892_6;

Selector_2 s3892_6(wires_973_5[0], addr_973_5, addr_positional[15571:15568], addr_3892_6);

wire[27:0] addr_3893_6;

Selector_2 s3893_6(wires_973_5[1], addr_973_5, addr_positional[15575:15572], addr_3893_6);

wire[27:0] addr_3894_6;

Selector_2 s3894_6(wires_973_5[2], addr_973_5, addr_positional[15579:15576], addr_3894_6);

wire[27:0] addr_3895_6;

Selector_2 s3895_6(wires_973_5[3], addr_973_5, addr_positional[15583:15580], addr_3895_6);

wire[27:0] addr_3896_6;

Selector_2 s3896_6(wires_974_5[0], addr_974_5, addr_positional[15587:15584], addr_3896_6);

wire[27:0] addr_3897_6;

Selector_2 s3897_6(wires_974_5[1], addr_974_5, addr_positional[15591:15588], addr_3897_6);

wire[27:0] addr_3898_6;

Selector_2 s3898_6(wires_974_5[2], addr_974_5, addr_positional[15595:15592], addr_3898_6);

wire[27:0] addr_3899_6;

Selector_2 s3899_6(wires_974_5[3], addr_974_5, addr_positional[15599:15596], addr_3899_6);

wire[27:0] addr_3900_6;

Selector_2 s3900_6(wires_975_5[0], addr_975_5, addr_positional[15603:15600], addr_3900_6);

wire[27:0] addr_3901_6;

Selector_2 s3901_6(wires_975_5[1], addr_975_5, addr_positional[15607:15604], addr_3901_6);

wire[27:0] addr_3902_6;

Selector_2 s3902_6(wires_975_5[2], addr_975_5, addr_positional[15611:15608], addr_3902_6);

wire[27:0] addr_3903_6;

Selector_2 s3903_6(wires_975_5[3], addr_975_5, addr_positional[15615:15612], addr_3903_6);

wire[27:0] addr_3904_6;

Selector_2 s3904_6(wires_976_5[0], addr_976_5, addr_positional[15619:15616], addr_3904_6);

wire[27:0] addr_3905_6;

Selector_2 s3905_6(wires_976_5[1], addr_976_5, addr_positional[15623:15620], addr_3905_6);

wire[27:0] addr_3906_6;

Selector_2 s3906_6(wires_976_5[2], addr_976_5, addr_positional[15627:15624], addr_3906_6);

wire[27:0] addr_3907_6;

Selector_2 s3907_6(wires_976_5[3], addr_976_5, addr_positional[15631:15628], addr_3907_6);

wire[27:0] addr_3908_6;

Selector_2 s3908_6(wires_977_5[0], addr_977_5, addr_positional[15635:15632], addr_3908_6);

wire[27:0] addr_3909_6;

Selector_2 s3909_6(wires_977_5[1], addr_977_5, addr_positional[15639:15636], addr_3909_6);

wire[27:0] addr_3910_6;

Selector_2 s3910_6(wires_977_5[2], addr_977_5, addr_positional[15643:15640], addr_3910_6);

wire[27:0] addr_3911_6;

Selector_2 s3911_6(wires_977_5[3], addr_977_5, addr_positional[15647:15644], addr_3911_6);

wire[27:0] addr_3912_6;

Selector_2 s3912_6(wires_978_5[0], addr_978_5, addr_positional[15651:15648], addr_3912_6);

wire[27:0] addr_3913_6;

Selector_2 s3913_6(wires_978_5[1], addr_978_5, addr_positional[15655:15652], addr_3913_6);

wire[27:0] addr_3914_6;

Selector_2 s3914_6(wires_978_5[2], addr_978_5, addr_positional[15659:15656], addr_3914_6);

wire[27:0] addr_3915_6;

Selector_2 s3915_6(wires_978_5[3], addr_978_5, addr_positional[15663:15660], addr_3915_6);

wire[27:0] addr_3916_6;

Selector_2 s3916_6(wires_979_5[0], addr_979_5, addr_positional[15667:15664], addr_3916_6);

wire[27:0] addr_3917_6;

Selector_2 s3917_6(wires_979_5[1], addr_979_5, addr_positional[15671:15668], addr_3917_6);

wire[27:0] addr_3918_6;

Selector_2 s3918_6(wires_979_5[2], addr_979_5, addr_positional[15675:15672], addr_3918_6);

wire[27:0] addr_3919_6;

Selector_2 s3919_6(wires_979_5[3], addr_979_5, addr_positional[15679:15676], addr_3919_6);

wire[27:0] addr_3920_6;

Selector_2 s3920_6(wires_980_5[0], addr_980_5, addr_positional[15683:15680], addr_3920_6);

wire[27:0] addr_3921_6;

Selector_2 s3921_6(wires_980_5[1], addr_980_5, addr_positional[15687:15684], addr_3921_6);

wire[27:0] addr_3922_6;

Selector_2 s3922_6(wires_980_5[2], addr_980_5, addr_positional[15691:15688], addr_3922_6);

wire[27:0] addr_3923_6;

Selector_2 s3923_6(wires_980_5[3], addr_980_5, addr_positional[15695:15692], addr_3923_6);

wire[27:0] addr_3924_6;

Selector_2 s3924_6(wires_981_5[0], addr_981_5, addr_positional[15699:15696], addr_3924_6);

wire[27:0] addr_3925_6;

Selector_2 s3925_6(wires_981_5[1], addr_981_5, addr_positional[15703:15700], addr_3925_6);

wire[27:0] addr_3926_6;

Selector_2 s3926_6(wires_981_5[2], addr_981_5, addr_positional[15707:15704], addr_3926_6);

wire[27:0] addr_3927_6;

Selector_2 s3927_6(wires_981_5[3], addr_981_5, addr_positional[15711:15708], addr_3927_6);

wire[27:0] addr_3928_6;

Selector_2 s3928_6(wires_982_5[0], addr_982_5, addr_positional[15715:15712], addr_3928_6);

wire[27:0] addr_3929_6;

Selector_2 s3929_6(wires_982_5[1], addr_982_5, addr_positional[15719:15716], addr_3929_6);

wire[27:0] addr_3930_6;

Selector_2 s3930_6(wires_982_5[2], addr_982_5, addr_positional[15723:15720], addr_3930_6);

wire[27:0] addr_3931_6;

Selector_2 s3931_6(wires_982_5[3], addr_982_5, addr_positional[15727:15724], addr_3931_6);

wire[27:0] addr_3932_6;

Selector_2 s3932_6(wires_983_5[0], addr_983_5, addr_positional[15731:15728], addr_3932_6);

wire[27:0] addr_3933_6;

Selector_2 s3933_6(wires_983_5[1], addr_983_5, addr_positional[15735:15732], addr_3933_6);

wire[27:0] addr_3934_6;

Selector_2 s3934_6(wires_983_5[2], addr_983_5, addr_positional[15739:15736], addr_3934_6);

wire[27:0] addr_3935_6;

Selector_2 s3935_6(wires_983_5[3], addr_983_5, addr_positional[15743:15740], addr_3935_6);

wire[27:0] addr_3936_6;

Selector_2 s3936_6(wires_984_5[0], addr_984_5, addr_positional[15747:15744], addr_3936_6);

wire[27:0] addr_3937_6;

Selector_2 s3937_6(wires_984_5[1], addr_984_5, addr_positional[15751:15748], addr_3937_6);

wire[27:0] addr_3938_6;

Selector_2 s3938_6(wires_984_5[2], addr_984_5, addr_positional[15755:15752], addr_3938_6);

wire[27:0] addr_3939_6;

Selector_2 s3939_6(wires_984_5[3], addr_984_5, addr_positional[15759:15756], addr_3939_6);

wire[27:0] addr_3940_6;

Selector_2 s3940_6(wires_985_5[0], addr_985_5, addr_positional[15763:15760], addr_3940_6);

wire[27:0] addr_3941_6;

Selector_2 s3941_6(wires_985_5[1], addr_985_5, addr_positional[15767:15764], addr_3941_6);

wire[27:0] addr_3942_6;

Selector_2 s3942_6(wires_985_5[2], addr_985_5, addr_positional[15771:15768], addr_3942_6);

wire[27:0] addr_3943_6;

Selector_2 s3943_6(wires_985_5[3], addr_985_5, addr_positional[15775:15772], addr_3943_6);

wire[27:0] addr_3944_6;

Selector_2 s3944_6(wires_986_5[0], addr_986_5, addr_positional[15779:15776], addr_3944_6);

wire[27:0] addr_3945_6;

Selector_2 s3945_6(wires_986_5[1], addr_986_5, addr_positional[15783:15780], addr_3945_6);

wire[27:0] addr_3946_6;

Selector_2 s3946_6(wires_986_5[2], addr_986_5, addr_positional[15787:15784], addr_3946_6);

wire[27:0] addr_3947_6;

Selector_2 s3947_6(wires_986_5[3], addr_986_5, addr_positional[15791:15788], addr_3947_6);

wire[27:0] addr_3948_6;

Selector_2 s3948_6(wires_987_5[0], addr_987_5, addr_positional[15795:15792], addr_3948_6);

wire[27:0] addr_3949_6;

Selector_2 s3949_6(wires_987_5[1], addr_987_5, addr_positional[15799:15796], addr_3949_6);

wire[27:0] addr_3950_6;

Selector_2 s3950_6(wires_987_5[2], addr_987_5, addr_positional[15803:15800], addr_3950_6);

wire[27:0] addr_3951_6;

Selector_2 s3951_6(wires_987_5[3], addr_987_5, addr_positional[15807:15804], addr_3951_6);

wire[27:0] addr_3952_6;

Selector_2 s3952_6(wires_988_5[0], addr_988_5, addr_positional[15811:15808], addr_3952_6);

wire[27:0] addr_3953_6;

Selector_2 s3953_6(wires_988_5[1], addr_988_5, addr_positional[15815:15812], addr_3953_6);

wire[27:0] addr_3954_6;

Selector_2 s3954_6(wires_988_5[2], addr_988_5, addr_positional[15819:15816], addr_3954_6);

wire[27:0] addr_3955_6;

Selector_2 s3955_6(wires_988_5[3], addr_988_5, addr_positional[15823:15820], addr_3955_6);

wire[27:0] addr_3956_6;

Selector_2 s3956_6(wires_989_5[0], addr_989_5, addr_positional[15827:15824], addr_3956_6);

wire[27:0] addr_3957_6;

Selector_2 s3957_6(wires_989_5[1], addr_989_5, addr_positional[15831:15828], addr_3957_6);

wire[27:0] addr_3958_6;

Selector_2 s3958_6(wires_989_5[2], addr_989_5, addr_positional[15835:15832], addr_3958_6);

wire[27:0] addr_3959_6;

Selector_2 s3959_6(wires_989_5[3], addr_989_5, addr_positional[15839:15836], addr_3959_6);

wire[27:0] addr_3960_6;

Selector_2 s3960_6(wires_990_5[0], addr_990_5, addr_positional[15843:15840], addr_3960_6);

wire[27:0] addr_3961_6;

Selector_2 s3961_6(wires_990_5[1], addr_990_5, addr_positional[15847:15844], addr_3961_6);

wire[27:0] addr_3962_6;

Selector_2 s3962_6(wires_990_5[2], addr_990_5, addr_positional[15851:15848], addr_3962_6);

wire[27:0] addr_3963_6;

Selector_2 s3963_6(wires_990_5[3], addr_990_5, addr_positional[15855:15852], addr_3963_6);

wire[27:0] addr_3964_6;

Selector_2 s3964_6(wires_991_5[0], addr_991_5, addr_positional[15859:15856], addr_3964_6);

wire[27:0] addr_3965_6;

Selector_2 s3965_6(wires_991_5[1], addr_991_5, addr_positional[15863:15860], addr_3965_6);

wire[27:0] addr_3966_6;

Selector_2 s3966_6(wires_991_5[2], addr_991_5, addr_positional[15867:15864], addr_3966_6);

wire[27:0] addr_3967_6;

Selector_2 s3967_6(wires_991_5[3], addr_991_5, addr_positional[15871:15868], addr_3967_6);

wire[27:0] addr_3968_6;

Selector_2 s3968_6(wires_992_5[0], addr_992_5, addr_positional[15875:15872], addr_3968_6);

wire[27:0] addr_3969_6;

Selector_2 s3969_6(wires_992_5[1], addr_992_5, addr_positional[15879:15876], addr_3969_6);

wire[27:0] addr_3970_6;

Selector_2 s3970_6(wires_992_5[2], addr_992_5, addr_positional[15883:15880], addr_3970_6);

wire[27:0] addr_3971_6;

Selector_2 s3971_6(wires_992_5[3], addr_992_5, addr_positional[15887:15884], addr_3971_6);

wire[27:0] addr_3972_6;

Selector_2 s3972_6(wires_993_5[0], addr_993_5, addr_positional[15891:15888], addr_3972_6);

wire[27:0] addr_3973_6;

Selector_2 s3973_6(wires_993_5[1], addr_993_5, addr_positional[15895:15892], addr_3973_6);

wire[27:0] addr_3974_6;

Selector_2 s3974_6(wires_993_5[2], addr_993_5, addr_positional[15899:15896], addr_3974_6);

wire[27:0] addr_3975_6;

Selector_2 s3975_6(wires_993_5[3], addr_993_5, addr_positional[15903:15900], addr_3975_6);

wire[27:0] addr_3976_6;

Selector_2 s3976_6(wires_994_5[0], addr_994_5, addr_positional[15907:15904], addr_3976_6);

wire[27:0] addr_3977_6;

Selector_2 s3977_6(wires_994_5[1], addr_994_5, addr_positional[15911:15908], addr_3977_6);

wire[27:0] addr_3978_6;

Selector_2 s3978_6(wires_994_5[2], addr_994_5, addr_positional[15915:15912], addr_3978_6);

wire[27:0] addr_3979_6;

Selector_2 s3979_6(wires_994_5[3], addr_994_5, addr_positional[15919:15916], addr_3979_6);

wire[27:0] addr_3980_6;

Selector_2 s3980_6(wires_995_5[0], addr_995_5, addr_positional[15923:15920], addr_3980_6);

wire[27:0] addr_3981_6;

Selector_2 s3981_6(wires_995_5[1], addr_995_5, addr_positional[15927:15924], addr_3981_6);

wire[27:0] addr_3982_6;

Selector_2 s3982_6(wires_995_5[2], addr_995_5, addr_positional[15931:15928], addr_3982_6);

wire[27:0] addr_3983_6;

Selector_2 s3983_6(wires_995_5[3], addr_995_5, addr_positional[15935:15932], addr_3983_6);

wire[27:0] addr_3984_6;

Selector_2 s3984_6(wires_996_5[0], addr_996_5, addr_positional[15939:15936], addr_3984_6);

wire[27:0] addr_3985_6;

Selector_2 s3985_6(wires_996_5[1], addr_996_5, addr_positional[15943:15940], addr_3985_6);

wire[27:0] addr_3986_6;

Selector_2 s3986_6(wires_996_5[2], addr_996_5, addr_positional[15947:15944], addr_3986_6);

wire[27:0] addr_3987_6;

Selector_2 s3987_6(wires_996_5[3], addr_996_5, addr_positional[15951:15948], addr_3987_6);

wire[27:0] addr_3988_6;

Selector_2 s3988_6(wires_997_5[0], addr_997_5, addr_positional[15955:15952], addr_3988_6);

wire[27:0] addr_3989_6;

Selector_2 s3989_6(wires_997_5[1], addr_997_5, addr_positional[15959:15956], addr_3989_6);

wire[27:0] addr_3990_6;

Selector_2 s3990_6(wires_997_5[2], addr_997_5, addr_positional[15963:15960], addr_3990_6);

wire[27:0] addr_3991_6;

Selector_2 s3991_6(wires_997_5[3], addr_997_5, addr_positional[15967:15964], addr_3991_6);

wire[27:0] addr_3992_6;

Selector_2 s3992_6(wires_998_5[0], addr_998_5, addr_positional[15971:15968], addr_3992_6);

wire[27:0] addr_3993_6;

Selector_2 s3993_6(wires_998_5[1], addr_998_5, addr_positional[15975:15972], addr_3993_6);

wire[27:0] addr_3994_6;

Selector_2 s3994_6(wires_998_5[2], addr_998_5, addr_positional[15979:15976], addr_3994_6);

wire[27:0] addr_3995_6;

Selector_2 s3995_6(wires_998_5[3], addr_998_5, addr_positional[15983:15980], addr_3995_6);

wire[27:0] addr_3996_6;

Selector_2 s3996_6(wires_999_5[0], addr_999_5, addr_positional[15987:15984], addr_3996_6);

wire[27:0] addr_3997_6;

Selector_2 s3997_6(wires_999_5[1], addr_999_5, addr_positional[15991:15988], addr_3997_6);

wire[27:0] addr_3998_6;

Selector_2 s3998_6(wires_999_5[2], addr_999_5, addr_positional[15995:15992], addr_3998_6);

wire[27:0] addr_3999_6;

Selector_2 s3999_6(wires_999_5[3], addr_999_5, addr_positional[15999:15996], addr_3999_6);

wire[27:0] addr_4000_6;

Selector_2 s4000_6(wires_1000_5[0], addr_1000_5, addr_positional[16003:16000], addr_4000_6);

wire[27:0] addr_4001_6;

Selector_2 s4001_6(wires_1000_5[1], addr_1000_5, addr_positional[16007:16004], addr_4001_6);

wire[27:0] addr_4002_6;

Selector_2 s4002_6(wires_1000_5[2], addr_1000_5, addr_positional[16011:16008], addr_4002_6);

wire[27:0] addr_4003_6;

Selector_2 s4003_6(wires_1000_5[3], addr_1000_5, addr_positional[16015:16012], addr_4003_6);

wire[27:0] addr_4004_6;

Selector_2 s4004_6(wires_1001_5[0], addr_1001_5, addr_positional[16019:16016], addr_4004_6);

wire[27:0] addr_4005_6;

Selector_2 s4005_6(wires_1001_5[1], addr_1001_5, addr_positional[16023:16020], addr_4005_6);

wire[27:0] addr_4006_6;

Selector_2 s4006_6(wires_1001_5[2], addr_1001_5, addr_positional[16027:16024], addr_4006_6);

wire[27:0] addr_4007_6;

Selector_2 s4007_6(wires_1001_5[3], addr_1001_5, addr_positional[16031:16028], addr_4007_6);

wire[27:0] addr_4008_6;

Selector_2 s4008_6(wires_1002_5[0], addr_1002_5, addr_positional[16035:16032], addr_4008_6);

wire[27:0] addr_4009_6;

Selector_2 s4009_6(wires_1002_5[1], addr_1002_5, addr_positional[16039:16036], addr_4009_6);

wire[27:0] addr_4010_6;

Selector_2 s4010_6(wires_1002_5[2], addr_1002_5, addr_positional[16043:16040], addr_4010_6);

wire[27:0] addr_4011_6;

Selector_2 s4011_6(wires_1002_5[3], addr_1002_5, addr_positional[16047:16044], addr_4011_6);

wire[27:0] addr_4012_6;

Selector_2 s4012_6(wires_1003_5[0], addr_1003_5, addr_positional[16051:16048], addr_4012_6);

wire[27:0] addr_4013_6;

Selector_2 s4013_6(wires_1003_5[1], addr_1003_5, addr_positional[16055:16052], addr_4013_6);

wire[27:0] addr_4014_6;

Selector_2 s4014_6(wires_1003_5[2], addr_1003_5, addr_positional[16059:16056], addr_4014_6);

wire[27:0] addr_4015_6;

Selector_2 s4015_6(wires_1003_5[3], addr_1003_5, addr_positional[16063:16060], addr_4015_6);

wire[27:0] addr_4016_6;

Selector_2 s4016_6(wires_1004_5[0], addr_1004_5, addr_positional[16067:16064], addr_4016_6);

wire[27:0] addr_4017_6;

Selector_2 s4017_6(wires_1004_5[1], addr_1004_5, addr_positional[16071:16068], addr_4017_6);

wire[27:0] addr_4018_6;

Selector_2 s4018_6(wires_1004_5[2], addr_1004_5, addr_positional[16075:16072], addr_4018_6);

wire[27:0] addr_4019_6;

Selector_2 s4019_6(wires_1004_5[3], addr_1004_5, addr_positional[16079:16076], addr_4019_6);

wire[27:0] addr_4020_6;

Selector_2 s4020_6(wires_1005_5[0], addr_1005_5, addr_positional[16083:16080], addr_4020_6);

wire[27:0] addr_4021_6;

Selector_2 s4021_6(wires_1005_5[1], addr_1005_5, addr_positional[16087:16084], addr_4021_6);

wire[27:0] addr_4022_6;

Selector_2 s4022_6(wires_1005_5[2], addr_1005_5, addr_positional[16091:16088], addr_4022_6);

wire[27:0] addr_4023_6;

Selector_2 s4023_6(wires_1005_5[3], addr_1005_5, addr_positional[16095:16092], addr_4023_6);

wire[27:0] addr_4024_6;

Selector_2 s4024_6(wires_1006_5[0], addr_1006_5, addr_positional[16099:16096], addr_4024_6);

wire[27:0] addr_4025_6;

Selector_2 s4025_6(wires_1006_5[1], addr_1006_5, addr_positional[16103:16100], addr_4025_6);

wire[27:0] addr_4026_6;

Selector_2 s4026_6(wires_1006_5[2], addr_1006_5, addr_positional[16107:16104], addr_4026_6);

wire[27:0] addr_4027_6;

Selector_2 s4027_6(wires_1006_5[3], addr_1006_5, addr_positional[16111:16108], addr_4027_6);

wire[27:0] addr_4028_6;

Selector_2 s4028_6(wires_1007_5[0], addr_1007_5, addr_positional[16115:16112], addr_4028_6);

wire[27:0] addr_4029_6;

Selector_2 s4029_6(wires_1007_5[1], addr_1007_5, addr_positional[16119:16116], addr_4029_6);

wire[27:0] addr_4030_6;

Selector_2 s4030_6(wires_1007_5[2], addr_1007_5, addr_positional[16123:16120], addr_4030_6);

wire[27:0] addr_4031_6;

Selector_2 s4031_6(wires_1007_5[3], addr_1007_5, addr_positional[16127:16124], addr_4031_6);

wire[27:0] addr_4032_6;

Selector_2 s4032_6(wires_1008_5[0], addr_1008_5, addr_positional[16131:16128], addr_4032_6);

wire[27:0] addr_4033_6;

Selector_2 s4033_6(wires_1008_5[1], addr_1008_5, addr_positional[16135:16132], addr_4033_6);

wire[27:0] addr_4034_6;

Selector_2 s4034_6(wires_1008_5[2], addr_1008_5, addr_positional[16139:16136], addr_4034_6);

wire[27:0] addr_4035_6;

Selector_2 s4035_6(wires_1008_5[3], addr_1008_5, addr_positional[16143:16140], addr_4035_6);

wire[27:0] addr_4036_6;

Selector_2 s4036_6(wires_1009_5[0], addr_1009_5, addr_positional[16147:16144], addr_4036_6);

wire[27:0] addr_4037_6;

Selector_2 s4037_6(wires_1009_5[1], addr_1009_5, addr_positional[16151:16148], addr_4037_6);

wire[27:0] addr_4038_6;

Selector_2 s4038_6(wires_1009_5[2], addr_1009_5, addr_positional[16155:16152], addr_4038_6);

wire[27:0] addr_4039_6;

Selector_2 s4039_6(wires_1009_5[3], addr_1009_5, addr_positional[16159:16156], addr_4039_6);

wire[27:0] addr_4040_6;

Selector_2 s4040_6(wires_1010_5[0], addr_1010_5, addr_positional[16163:16160], addr_4040_6);

wire[27:0] addr_4041_6;

Selector_2 s4041_6(wires_1010_5[1], addr_1010_5, addr_positional[16167:16164], addr_4041_6);

wire[27:0] addr_4042_6;

Selector_2 s4042_6(wires_1010_5[2], addr_1010_5, addr_positional[16171:16168], addr_4042_6);

wire[27:0] addr_4043_6;

Selector_2 s4043_6(wires_1010_5[3], addr_1010_5, addr_positional[16175:16172], addr_4043_6);

wire[27:0] addr_4044_6;

Selector_2 s4044_6(wires_1011_5[0], addr_1011_5, addr_positional[16179:16176], addr_4044_6);

wire[27:0] addr_4045_6;

Selector_2 s4045_6(wires_1011_5[1], addr_1011_5, addr_positional[16183:16180], addr_4045_6);

wire[27:0] addr_4046_6;

Selector_2 s4046_6(wires_1011_5[2], addr_1011_5, addr_positional[16187:16184], addr_4046_6);

wire[27:0] addr_4047_6;

Selector_2 s4047_6(wires_1011_5[3], addr_1011_5, addr_positional[16191:16188], addr_4047_6);

wire[27:0] addr_4048_6;

Selector_2 s4048_6(wires_1012_5[0], addr_1012_5, addr_positional[16195:16192], addr_4048_6);

wire[27:0] addr_4049_6;

Selector_2 s4049_6(wires_1012_5[1], addr_1012_5, addr_positional[16199:16196], addr_4049_6);

wire[27:0] addr_4050_6;

Selector_2 s4050_6(wires_1012_5[2], addr_1012_5, addr_positional[16203:16200], addr_4050_6);

wire[27:0] addr_4051_6;

Selector_2 s4051_6(wires_1012_5[3], addr_1012_5, addr_positional[16207:16204], addr_4051_6);

wire[27:0] addr_4052_6;

Selector_2 s4052_6(wires_1013_5[0], addr_1013_5, addr_positional[16211:16208], addr_4052_6);

wire[27:0] addr_4053_6;

Selector_2 s4053_6(wires_1013_5[1], addr_1013_5, addr_positional[16215:16212], addr_4053_6);

wire[27:0] addr_4054_6;

Selector_2 s4054_6(wires_1013_5[2], addr_1013_5, addr_positional[16219:16216], addr_4054_6);

wire[27:0] addr_4055_6;

Selector_2 s4055_6(wires_1013_5[3], addr_1013_5, addr_positional[16223:16220], addr_4055_6);

wire[27:0] addr_4056_6;

Selector_2 s4056_6(wires_1014_5[0], addr_1014_5, addr_positional[16227:16224], addr_4056_6);

wire[27:0] addr_4057_6;

Selector_2 s4057_6(wires_1014_5[1], addr_1014_5, addr_positional[16231:16228], addr_4057_6);

wire[27:0] addr_4058_6;

Selector_2 s4058_6(wires_1014_5[2], addr_1014_5, addr_positional[16235:16232], addr_4058_6);

wire[27:0] addr_4059_6;

Selector_2 s4059_6(wires_1014_5[3], addr_1014_5, addr_positional[16239:16236], addr_4059_6);

wire[27:0] addr_4060_6;

Selector_2 s4060_6(wires_1015_5[0], addr_1015_5, addr_positional[16243:16240], addr_4060_6);

wire[27:0] addr_4061_6;

Selector_2 s4061_6(wires_1015_5[1], addr_1015_5, addr_positional[16247:16244], addr_4061_6);

wire[27:0] addr_4062_6;

Selector_2 s4062_6(wires_1015_5[2], addr_1015_5, addr_positional[16251:16248], addr_4062_6);

wire[27:0] addr_4063_6;

Selector_2 s4063_6(wires_1015_5[3], addr_1015_5, addr_positional[16255:16252], addr_4063_6);

wire[27:0] addr_4064_6;

Selector_2 s4064_6(wires_1016_5[0], addr_1016_5, addr_positional[16259:16256], addr_4064_6);

wire[27:0] addr_4065_6;

Selector_2 s4065_6(wires_1016_5[1], addr_1016_5, addr_positional[16263:16260], addr_4065_6);

wire[27:0] addr_4066_6;

Selector_2 s4066_6(wires_1016_5[2], addr_1016_5, addr_positional[16267:16264], addr_4066_6);

wire[27:0] addr_4067_6;

Selector_2 s4067_6(wires_1016_5[3], addr_1016_5, addr_positional[16271:16268], addr_4067_6);

wire[27:0] addr_4068_6;

Selector_2 s4068_6(wires_1017_5[0], addr_1017_5, addr_positional[16275:16272], addr_4068_6);

wire[27:0] addr_4069_6;

Selector_2 s4069_6(wires_1017_5[1], addr_1017_5, addr_positional[16279:16276], addr_4069_6);

wire[27:0] addr_4070_6;

Selector_2 s4070_6(wires_1017_5[2], addr_1017_5, addr_positional[16283:16280], addr_4070_6);

wire[27:0] addr_4071_6;

Selector_2 s4071_6(wires_1017_5[3], addr_1017_5, addr_positional[16287:16284], addr_4071_6);

wire[27:0] addr_4072_6;

Selector_2 s4072_6(wires_1018_5[0], addr_1018_5, addr_positional[16291:16288], addr_4072_6);

wire[27:0] addr_4073_6;

Selector_2 s4073_6(wires_1018_5[1], addr_1018_5, addr_positional[16295:16292], addr_4073_6);

wire[27:0] addr_4074_6;

Selector_2 s4074_6(wires_1018_5[2], addr_1018_5, addr_positional[16299:16296], addr_4074_6);

wire[27:0] addr_4075_6;

Selector_2 s4075_6(wires_1018_5[3], addr_1018_5, addr_positional[16303:16300], addr_4075_6);

wire[27:0] addr_4076_6;

Selector_2 s4076_6(wires_1019_5[0], addr_1019_5, addr_positional[16307:16304], addr_4076_6);

wire[27:0] addr_4077_6;

Selector_2 s4077_6(wires_1019_5[1], addr_1019_5, addr_positional[16311:16308], addr_4077_6);

wire[27:0] addr_4078_6;

Selector_2 s4078_6(wires_1019_5[2], addr_1019_5, addr_positional[16315:16312], addr_4078_6);

wire[27:0] addr_4079_6;

Selector_2 s4079_6(wires_1019_5[3], addr_1019_5, addr_positional[16319:16316], addr_4079_6);

wire[27:0] addr_4080_6;

Selector_2 s4080_6(wires_1020_5[0], addr_1020_5, addr_positional[16323:16320], addr_4080_6);

wire[27:0] addr_4081_6;

Selector_2 s4081_6(wires_1020_5[1], addr_1020_5, addr_positional[16327:16324], addr_4081_6);

wire[27:0] addr_4082_6;

Selector_2 s4082_6(wires_1020_5[2], addr_1020_5, addr_positional[16331:16328], addr_4082_6);

wire[27:0] addr_4083_6;

Selector_2 s4083_6(wires_1020_5[3], addr_1020_5, addr_positional[16335:16332], addr_4083_6);

wire[27:0] addr_4084_6;

Selector_2 s4084_6(wires_1021_5[0], addr_1021_5, addr_positional[16339:16336], addr_4084_6);

wire[27:0] addr_4085_6;

Selector_2 s4085_6(wires_1021_5[1], addr_1021_5, addr_positional[16343:16340], addr_4085_6);

wire[27:0] addr_4086_6;

Selector_2 s4086_6(wires_1021_5[2], addr_1021_5, addr_positional[16347:16344], addr_4086_6);

wire[27:0] addr_4087_6;

Selector_2 s4087_6(wires_1021_5[3], addr_1021_5, addr_positional[16351:16348], addr_4087_6);

wire[27:0] addr_4088_6;

Selector_2 s4088_6(wires_1022_5[0], addr_1022_5, addr_positional[16355:16352], addr_4088_6);

wire[27:0] addr_4089_6;

Selector_2 s4089_6(wires_1022_5[1], addr_1022_5, addr_positional[16359:16356], addr_4089_6);

wire[27:0] addr_4090_6;

Selector_2 s4090_6(wires_1022_5[2], addr_1022_5, addr_positional[16363:16360], addr_4090_6);

wire[27:0] addr_4091_6;

Selector_2 s4091_6(wires_1022_5[3], addr_1022_5, addr_positional[16367:16364], addr_4091_6);

wire[27:0] addr_4092_6;

Selector_2 s4092_6(wires_1023_5[0], addr_1023_5, addr_positional[16371:16368], addr_4092_6);

wire[27:0] addr_4093_6;

Selector_2 s4093_6(wires_1023_5[1], addr_1023_5, addr_positional[16375:16372], addr_4093_6);

wire[27:0] addr_4094_6;

Selector_2 s4094_6(wires_1023_5[2], addr_1023_5, addr_positional[16379:16376], addr_4094_6);

wire[27:0] addr_4095_6;

Selector_2 s4095_6(wires_1023_5[3], addr_1023_5, addr_positional[16383:16380], addr_4095_6);



endmodule

