module address_decode_2
(

    input wire[1:0] addr_src,

    output wire[3:0] addr_positional
);



assign addr_positional[3] = (addr_src==2'b11) ?1'b1:1'b0;

assign addr_positional[2] = (addr_src==2'b10) ?1'b1:1'b0;

assign addr_positional[1] = (addr_src==2'b01) ?1'b1:1'b0;

assign addr_positional[0] = (addr_src==2'b00) ?1'b1:1'b0;



endmodule

module address_decode_16
(

    input wire[15:0] addr_src,

    output wire[31:0] addr_positional
);



address_decode_2 enc0(addr_src[1:0], addr_positional[31:28]);

address_decode_2 enc1(addr_src[3:2], addr_positional[27:24]);

address_decode_2 enc2(addr_src[5:4], addr_positional[23:20]);

address_decode_2 enc3(addr_src[7:6], addr_positional[19:16]);

address_decode_2 enc4(addr_src[9:8], addr_positional[15:12]);

address_decode_2 enc5(addr_src[11:10], addr_positional[11:8]);

address_decode_2 enc6(addr_src[13:12], addr_positional[7:4]);

address_decode_2 enc7(addr_src[15:14], addr_positional[3:0]);



endmodule

module Selector_2
(

    input wire selector_enabled,

    input wire[31:0] addr_src,

    output wire[3:0] addr_positional,

    output wire[31:0] addr_remain
);




assign addr_remain =        (selector_enabled==1'b1)? {4'b0,addr_src[31:4]}:32'b0;
assign addr_positional =    (selector_enabled==1'b1)? addr_src[3:0] : 4'b0;

endmodule



module Selector_16
(

    input wire[15:0] addr,

    output wire[65535:0] addr_positional
);





 

   wire[31:0] addr_src;

   address_decode_16 sel_1 (addr, addr_src);wire[3:0] wires_0_0;

wire[31:0] addr_0_0;

Selector_2 s0_0(1'b1, addr_src, wires_0_0, addr_0_0);

wire[3:0] wires_0_1;

wire[31:0] addr_0_1;

Selector_2 s0_1(wires_0_0[0], addr_0_0, wires_0_1,addr_0_1);

wire[3:0] wires_1_1;

wire[31:0] addr_1_1;

Selector_2 s1_1(wires_0_0[1], addr_0_0, wires_1_1,addr_1_1);

wire[3:0] wires_2_1;

wire[31:0] addr_2_1;

Selector_2 s2_1(wires_0_0[2], addr_0_0, wires_2_1,addr_2_1);

wire[3:0] wires_3_1;

wire[31:0] addr_3_1;

Selector_2 s3_1(wires_0_0[3], addr_0_0, wires_3_1,addr_3_1);

wire[3:0] wires_0_2;

wire[31:0] addr_0_2;

Selector_2 s0_2(wires_0_1[0], addr_0_1, wires_0_2,addr_0_2);

wire[3:0] wires_1_2;

wire[31:0] addr_1_2;

Selector_2 s1_2(wires_0_1[1], addr_0_1, wires_1_2,addr_1_2);

wire[3:0] wires_2_2;

wire[31:0] addr_2_2;

Selector_2 s2_2(wires_0_1[2], addr_0_1, wires_2_2,addr_2_2);

wire[3:0] wires_3_2;

wire[31:0] addr_3_2;

Selector_2 s3_2(wires_0_1[3], addr_0_1, wires_3_2,addr_3_2);

wire[3:0] wires_4_2;

wire[31:0] addr_4_2;

Selector_2 s4_2(wires_1_1[0], addr_1_1, wires_4_2,addr_4_2);

wire[3:0] wires_5_2;

wire[31:0] addr_5_2;

Selector_2 s5_2(wires_1_1[1], addr_1_1, wires_5_2,addr_5_2);

wire[3:0] wires_6_2;

wire[31:0] addr_6_2;

Selector_2 s6_2(wires_1_1[2], addr_1_1, wires_6_2,addr_6_2);

wire[3:0] wires_7_2;

wire[31:0] addr_7_2;

Selector_2 s7_2(wires_1_1[3], addr_1_1, wires_7_2,addr_7_2);

wire[3:0] wires_8_2;

wire[31:0] addr_8_2;

Selector_2 s8_2(wires_2_1[0], addr_2_1, wires_8_2,addr_8_2);

wire[3:0] wires_9_2;

wire[31:0] addr_9_2;

Selector_2 s9_2(wires_2_1[1], addr_2_1, wires_9_2,addr_9_2);

wire[3:0] wires_10_2;

wire[31:0] addr_10_2;

Selector_2 s10_2(wires_2_1[2], addr_2_1, wires_10_2,addr_10_2);

wire[3:0] wires_11_2;

wire[31:0] addr_11_2;

Selector_2 s11_2(wires_2_1[3], addr_2_1, wires_11_2,addr_11_2);

wire[3:0] wires_12_2;

wire[31:0] addr_12_2;

Selector_2 s12_2(wires_3_1[0], addr_3_1, wires_12_2,addr_12_2);

wire[3:0] wires_13_2;

wire[31:0] addr_13_2;

Selector_2 s13_2(wires_3_1[1], addr_3_1, wires_13_2,addr_13_2);

wire[3:0] wires_14_2;

wire[31:0] addr_14_2;

Selector_2 s14_2(wires_3_1[2], addr_3_1, wires_14_2,addr_14_2);

wire[3:0] wires_15_2;

wire[31:0] addr_15_2;

Selector_2 s15_2(wires_3_1[3], addr_3_1, wires_15_2,addr_15_2);

wire[3:0] wires_0_3;

wire[31:0] addr_0_3;

Selector_2 s0_3(wires_0_2[0], addr_0_2, wires_0_3,addr_0_3);

wire[3:0] wires_1_3;

wire[31:0] addr_1_3;

Selector_2 s1_3(wires_0_2[1], addr_0_2, wires_1_3,addr_1_3);

wire[3:0] wires_2_3;

wire[31:0] addr_2_3;

Selector_2 s2_3(wires_0_2[2], addr_0_2, wires_2_3,addr_2_3);

wire[3:0] wires_3_3;

wire[31:0] addr_3_3;

Selector_2 s3_3(wires_0_2[3], addr_0_2, wires_3_3,addr_3_3);

wire[3:0] wires_4_3;

wire[31:0] addr_4_3;

Selector_2 s4_3(wires_1_2[0], addr_1_2, wires_4_3,addr_4_3);

wire[3:0] wires_5_3;

wire[31:0] addr_5_3;

Selector_2 s5_3(wires_1_2[1], addr_1_2, wires_5_3,addr_5_3);

wire[3:0] wires_6_3;

wire[31:0] addr_6_3;

Selector_2 s6_3(wires_1_2[2], addr_1_2, wires_6_3,addr_6_3);

wire[3:0] wires_7_3;

wire[31:0] addr_7_3;

Selector_2 s7_3(wires_1_2[3], addr_1_2, wires_7_3,addr_7_3);

wire[3:0] wires_8_3;

wire[31:0] addr_8_3;

Selector_2 s8_3(wires_2_2[0], addr_2_2, wires_8_3,addr_8_3);

wire[3:0] wires_9_3;

wire[31:0] addr_9_3;

Selector_2 s9_3(wires_2_2[1], addr_2_2, wires_9_3,addr_9_3);

wire[3:0] wires_10_3;

wire[31:0] addr_10_3;

Selector_2 s10_3(wires_2_2[2], addr_2_2, wires_10_3,addr_10_3);

wire[3:0] wires_11_3;

wire[31:0] addr_11_3;

Selector_2 s11_3(wires_2_2[3], addr_2_2, wires_11_3,addr_11_3);

wire[3:0] wires_12_3;

wire[31:0] addr_12_3;

Selector_2 s12_3(wires_3_2[0], addr_3_2, wires_12_3,addr_12_3);

wire[3:0] wires_13_3;

wire[31:0] addr_13_3;

Selector_2 s13_3(wires_3_2[1], addr_3_2, wires_13_3,addr_13_3);

wire[3:0] wires_14_3;

wire[31:0] addr_14_3;

Selector_2 s14_3(wires_3_2[2], addr_3_2, wires_14_3,addr_14_3);

wire[3:0] wires_15_3;

wire[31:0] addr_15_3;

Selector_2 s15_3(wires_3_2[3], addr_3_2, wires_15_3,addr_15_3);

wire[3:0] wires_16_3;

wire[31:0] addr_16_3;

Selector_2 s16_3(wires_4_2[0], addr_4_2, wires_16_3,addr_16_3);

wire[3:0] wires_17_3;

wire[31:0] addr_17_3;

Selector_2 s17_3(wires_4_2[1], addr_4_2, wires_17_3,addr_17_3);

wire[3:0] wires_18_3;

wire[31:0] addr_18_3;

Selector_2 s18_3(wires_4_2[2], addr_4_2, wires_18_3,addr_18_3);

wire[3:0] wires_19_3;

wire[31:0] addr_19_3;

Selector_2 s19_3(wires_4_2[3], addr_4_2, wires_19_3,addr_19_3);

wire[3:0] wires_20_3;

wire[31:0] addr_20_3;

Selector_2 s20_3(wires_5_2[0], addr_5_2, wires_20_3,addr_20_3);

wire[3:0] wires_21_3;

wire[31:0] addr_21_3;

Selector_2 s21_3(wires_5_2[1], addr_5_2, wires_21_3,addr_21_3);

wire[3:0] wires_22_3;

wire[31:0] addr_22_3;

Selector_2 s22_3(wires_5_2[2], addr_5_2, wires_22_3,addr_22_3);

wire[3:0] wires_23_3;

wire[31:0] addr_23_3;

Selector_2 s23_3(wires_5_2[3], addr_5_2, wires_23_3,addr_23_3);

wire[3:0] wires_24_3;

wire[31:0] addr_24_3;

Selector_2 s24_3(wires_6_2[0], addr_6_2, wires_24_3,addr_24_3);

wire[3:0] wires_25_3;

wire[31:0] addr_25_3;

Selector_2 s25_3(wires_6_2[1], addr_6_2, wires_25_3,addr_25_3);

wire[3:0] wires_26_3;

wire[31:0] addr_26_3;

Selector_2 s26_3(wires_6_2[2], addr_6_2, wires_26_3,addr_26_3);

wire[3:0] wires_27_3;

wire[31:0] addr_27_3;

Selector_2 s27_3(wires_6_2[3], addr_6_2, wires_27_3,addr_27_3);

wire[3:0] wires_28_3;

wire[31:0] addr_28_3;

Selector_2 s28_3(wires_7_2[0], addr_7_2, wires_28_3,addr_28_3);

wire[3:0] wires_29_3;

wire[31:0] addr_29_3;

Selector_2 s29_3(wires_7_2[1], addr_7_2, wires_29_3,addr_29_3);

wire[3:0] wires_30_3;

wire[31:0] addr_30_3;

Selector_2 s30_3(wires_7_2[2], addr_7_2, wires_30_3,addr_30_3);

wire[3:0] wires_31_3;

wire[31:0] addr_31_3;

Selector_2 s31_3(wires_7_2[3], addr_7_2, wires_31_3,addr_31_3);

wire[3:0] wires_32_3;

wire[31:0] addr_32_3;

Selector_2 s32_3(wires_8_2[0], addr_8_2, wires_32_3,addr_32_3);

wire[3:0] wires_33_3;

wire[31:0] addr_33_3;

Selector_2 s33_3(wires_8_2[1], addr_8_2, wires_33_3,addr_33_3);

wire[3:0] wires_34_3;

wire[31:0] addr_34_3;

Selector_2 s34_3(wires_8_2[2], addr_8_2, wires_34_3,addr_34_3);

wire[3:0] wires_35_3;

wire[31:0] addr_35_3;

Selector_2 s35_3(wires_8_2[3], addr_8_2, wires_35_3,addr_35_3);

wire[3:0] wires_36_3;

wire[31:0] addr_36_3;

Selector_2 s36_3(wires_9_2[0], addr_9_2, wires_36_3,addr_36_3);

wire[3:0] wires_37_3;

wire[31:0] addr_37_3;

Selector_2 s37_3(wires_9_2[1], addr_9_2, wires_37_3,addr_37_3);

wire[3:0] wires_38_3;

wire[31:0] addr_38_3;

Selector_2 s38_3(wires_9_2[2], addr_9_2, wires_38_3,addr_38_3);

wire[3:0] wires_39_3;

wire[31:0] addr_39_3;

Selector_2 s39_3(wires_9_2[3], addr_9_2, wires_39_3,addr_39_3);

wire[3:0] wires_40_3;

wire[31:0] addr_40_3;

Selector_2 s40_3(wires_10_2[0], addr_10_2, wires_40_3,addr_40_3);

wire[3:0] wires_41_3;

wire[31:0] addr_41_3;

Selector_2 s41_3(wires_10_2[1], addr_10_2, wires_41_3,addr_41_3);

wire[3:0] wires_42_3;

wire[31:0] addr_42_3;

Selector_2 s42_3(wires_10_2[2], addr_10_2, wires_42_3,addr_42_3);

wire[3:0] wires_43_3;

wire[31:0] addr_43_3;

Selector_2 s43_3(wires_10_2[3], addr_10_2, wires_43_3,addr_43_3);

wire[3:0] wires_44_3;

wire[31:0] addr_44_3;

Selector_2 s44_3(wires_11_2[0], addr_11_2, wires_44_3,addr_44_3);

wire[3:0] wires_45_3;

wire[31:0] addr_45_3;

Selector_2 s45_3(wires_11_2[1], addr_11_2, wires_45_3,addr_45_3);

wire[3:0] wires_46_3;

wire[31:0] addr_46_3;

Selector_2 s46_3(wires_11_2[2], addr_11_2, wires_46_3,addr_46_3);

wire[3:0] wires_47_3;

wire[31:0] addr_47_3;

Selector_2 s47_3(wires_11_2[3], addr_11_2, wires_47_3,addr_47_3);

wire[3:0] wires_48_3;

wire[31:0] addr_48_3;

Selector_2 s48_3(wires_12_2[0], addr_12_2, wires_48_3,addr_48_3);

wire[3:0] wires_49_3;

wire[31:0] addr_49_3;

Selector_2 s49_3(wires_12_2[1], addr_12_2, wires_49_3,addr_49_3);

wire[3:0] wires_50_3;

wire[31:0] addr_50_3;

Selector_2 s50_3(wires_12_2[2], addr_12_2, wires_50_3,addr_50_3);

wire[3:0] wires_51_3;

wire[31:0] addr_51_3;

Selector_2 s51_3(wires_12_2[3], addr_12_2, wires_51_3,addr_51_3);

wire[3:0] wires_52_3;

wire[31:0] addr_52_3;

Selector_2 s52_3(wires_13_2[0], addr_13_2, wires_52_3,addr_52_3);

wire[3:0] wires_53_3;

wire[31:0] addr_53_3;

Selector_2 s53_3(wires_13_2[1], addr_13_2, wires_53_3,addr_53_3);

wire[3:0] wires_54_3;

wire[31:0] addr_54_3;

Selector_2 s54_3(wires_13_2[2], addr_13_2, wires_54_3,addr_54_3);

wire[3:0] wires_55_3;

wire[31:0] addr_55_3;

Selector_2 s55_3(wires_13_2[3], addr_13_2, wires_55_3,addr_55_3);

wire[3:0] wires_56_3;

wire[31:0] addr_56_3;

Selector_2 s56_3(wires_14_2[0], addr_14_2, wires_56_3,addr_56_3);

wire[3:0] wires_57_3;

wire[31:0] addr_57_3;

Selector_2 s57_3(wires_14_2[1], addr_14_2, wires_57_3,addr_57_3);

wire[3:0] wires_58_3;

wire[31:0] addr_58_3;

Selector_2 s58_3(wires_14_2[2], addr_14_2, wires_58_3,addr_58_3);

wire[3:0] wires_59_3;

wire[31:0] addr_59_3;

Selector_2 s59_3(wires_14_2[3], addr_14_2, wires_59_3,addr_59_3);

wire[3:0] wires_60_3;

wire[31:0] addr_60_3;

Selector_2 s60_3(wires_15_2[0], addr_15_2, wires_60_3,addr_60_3);

wire[3:0] wires_61_3;

wire[31:0] addr_61_3;

Selector_2 s61_3(wires_15_2[1], addr_15_2, wires_61_3,addr_61_3);

wire[3:0] wires_62_3;

wire[31:0] addr_62_3;

Selector_2 s62_3(wires_15_2[2], addr_15_2, wires_62_3,addr_62_3);

wire[3:0] wires_63_3;

wire[31:0] addr_63_3;

Selector_2 s63_3(wires_15_2[3], addr_15_2, wires_63_3,addr_63_3);

wire[3:0] wires_0_4;

wire[31:0] addr_0_4;

Selector_2 s0_4(wires_0_3[0], addr_0_3, wires_0_4,addr_0_4);

wire[3:0] wires_1_4;

wire[31:0] addr_1_4;

Selector_2 s1_4(wires_0_3[1], addr_0_3, wires_1_4,addr_1_4);

wire[3:0] wires_2_4;

wire[31:0] addr_2_4;

Selector_2 s2_4(wires_0_3[2], addr_0_3, wires_2_4,addr_2_4);

wire[3:0] wires_3_4;

wire[31:0] addr_3_4;

Selector_2 s3_4(wires_0_3[3], addr_0_3, wires_3_4,addr_3_4);

wire[3:0] wires_4_4;

wire[31:0] addr_4_4;

Selector_2 s4_4(wires_1_3[0], addr_1_3, wires_4_4,addr_4_4);

wire[3:0] wires_5_4;

wire[31:0] addr_5_4;

Selector_2 s5_4(wires_1_3[1], addr_1_3, wires_5_4,addr_5_4);

wire[3:0] wires_6_4;

wire[31:0] addr_6_4;

Selector_2 s6_4(wires_1_3[2], addr_1_3, wires_6_4,addr_6_4);

wire[3:0] wires_7_4;

wire[31:0] addr_7_4;

Selector_2 s7_4(wires_1_3[3], addr_1_3, wires_7_4,addr_7_4);

wire[3:0] wires_8_4;

wire[31:0] addr_8_4;

Selector_2 s8_4(wires_2_3[0], addr_2_3, wires_8_4,addr_8_4);

wire[3:0] wires_9_4;

wire[31:0] addr_9_4;

Selector_2 s9_4(wires_2_3[1], addr_2_3, wires_9_4,addr_9_4);

wire[3:0] wires_10_4;

wire[31:0] addr_10_4;

Selector_2 s10_4(wires_2_3[2], addr_2_3, wires_10_4,addr_10_4);

wire[3:0] wires_11_4;

wire[31:0] addr_11_4;

Selector_2 s11_4(wires_2_3[3], addr_2_3, wires_11_4,addr_11_4);

wire[3:0] wires_12_4;

wire[31:0] addr_12_4;

Selector_2 s12_4(wires_3_3[0], addr_3_3, wires_12_4,addr_12_4);

wire[3:0] wires_13_4;

wire[31:0] addr_13_4;

Selector_2 s13_4(wires_3_3[1], addr_3_3, wires_13_4,addr_13_4);

wire[3:0] wires_14_4;

wire[31:0] addr_14_4;

Selector_2 s14_4(wires_3_3[2], addr_3_3, wires_14_4,addr_14_4);

wire[3:0] wires_15_4;

wire[31:0] addr_15_4;

Selector_2 s15_4(wires_3_3[3], addr_3_3, wires_15_4,addr_15_4);

wire[3:0] wires_16_4;

wire[31:0] addr_16_4;

Selector_2 s16_4(wires_4_3[0], addr_4_3, wires_16_4,addr_16_4);

wire[3:0] wires_17_4;

wire[31:0] addr_17_4;

Selector_2 s17_4(wires_4_3[1], addr_4_3, wires_17_4,addr_17_4);

wire[3:0] wires_18_4;

wire[31:0] addr_18_4;

Selector_2 s18_4(wires_4_3[2], addr_4_3, wires_18_4,addr_18_4);

wire[3:0] wires_19_4;

wire[31:0] addr_19_4;

Selector_2 s19_4(wires_4_3[3], addr_4_3, wires_19_4,addr_19_4);

wire[3:0] wires_20_4;

wire[31:0] addr_20_4;

Selector_2 s20_4(wires_5_3[0], addr_5_3, wires_20_4,addr_20_4);

wire[3:0] wires_21_4;

wire[31:0] addr_21_4;

Selector_2 s21_4(wires_5_3[1], addr_5_3, wires_21_4,addr_21_4);

wire[3:0] wires_22_4;

wire[31:0] addr_22_4;

Selector_2 s22_4(wires_5_3[2], addr_5_3, wires_22_4,addr_22_4);

wire[3:0] wires_23_4;

wire[31:0] addr_23_4;

Selector_2 s23_4(wires_5_3[3], addr_5_3, wires_23_4,addr_23_4);

wire[3:0] wires_24_4;

wire[31:0] addr_24_4;

Selector_2 s24_4(wires_6_3[0], addr_6_3, wires_24_4,addr_24_4);

wire[3:0] wires_25_4;

wire[31:0] addr_25_4;

Selector_2 s25_4(wires_6_3[1], addr_6_3, wires_25_4,addr_25_4);

wire[3:0] wires_26_4;

wire[31:0] addr_26_4;

Selector_2 s26_4(wires_6_3[2], addr_6_3, wires_26_4,addr_26_4);

wire[3:0] wires_27_4;

wire[31:0] addr_27_4;

Selector_2 s27_4(wires_6_3[3], addr_6_3, wires_27_4,addr_27_4);

wire[3:0] wires_28_4;

wire[31:0] addr_28_4;

Selector_2 s28_4(wires_7_3[0], addr_7_3, wires_28_4,addr_28_4);

wire[3:0] wires_29_4;

wire[31:0] addr_29_4;

Selector_2 s29_4(wires_7_3[1], addr_7_3, wires_29_4,addr_29_4);

wire[3:0] wires_30_4;

wire[31:0] addr_30_4;

Selector_2 s30_4(wires_7_3[2], addr_7_3, wires_30_4,addr_30_4);

wire[3:0] wires_31_4;

wire[31:0] addr_31_4;

Selector_2 s31_4(wires_7_3[3], addr_7_3, wires_31_4,addr_31_4);

wire[3:0] wires_32_4;

wire[31:0] addr_32_4;

Selector_2 s32_4(wires_8_3[0], addr_8_3, wires_32_4,addr_32_4);

wire[3:0] wires_33_4;

wire[31:0] addr_33_4;

Selector_2 s33_4(wires_8_3[1], addr_8_3, wires_33_4,addr_33_4);

wire[3:0] wires_34_4;

wire[31:0] addr_34_4;

Selector_2 s34_4(wires_8_3[2], addr_8_3, wires_34_4,addr_34_4);

wire[3:0] wires_35_4;

wire[31:0] addr_35_4;

Selector_2 s35_4(wires_8_3[3], addr_8_3, wires_35_4,addr_35_4);

wire[3:0] wires_36_4;

wire[31:0] addr_36_4;

Selector_2 s36_4(wires_9_3[0], addr_9_3, wires_36_4,addr_36_4);

wire[3:0] wires_37_4;

wire[31:0] addr_37_4;

Selector_2 s37_4(wires_9_3[1], addr_9_3, wires_37_4,addr_37_4);

wire[3:0] wires_38_4;

wire[31:0] addr_38_4;

Selector_2 s38_4(wires_9_3[2], addr_9_3, wires_38_4,addr_38_4);

wire[3:0] wires_39_4;

wire[31:0] addr_39_4;

Selector_2 s39_4(wires_9_3[3], addr_9_3, wires_39_4,addr_39_4);

wire[3:0] wires_40_4;

wire[31:0] addr_40_4;

Selector_2 s40_4(wires_10_3[0], addr_10_3, wires_40_4,addr_40_4);

wire[3:0] wires_41_4;

wire[31:0] addr_41_4;

Selector_2 s41_4(wires_10_3[1], addr_10_3, wires_41_4,addr_41_4);

wire[3:0] wires_42_4;

wire[31:0] addr_42_4;

Selector_2 s42_4(wires_10_3[2], addr_10_3, wires_42_4,addr_42_4);

wire[3:0] wires_43_4;

wire[31:0] addr_43_4;

Selector_2 s43_4(wires_10_3[3], addr_10_3, wires_43_4,addr_43_4);

wire[3:0] wires_44_4;

wire[31:0] addr_44_4;

Selector_2 s44_4(wires_11_3[0], addr_11_3, wires_44_4,addr_44_4);

wire[3:0] wires_45_4;

wire[31:0] addr_45_4;

Selector_2 s45_4(wires_11_3[1], addr_11_3, wires_45_4,addr_45_4);

wire[3:0] wires_46_4;

wire[31:0] addr_46_4;

Selector_2 s46_4(wires_11_3[2], addr_11_3, wires_46_4,addr_46_4);

wire[3:0] wires_47_4;

wire[31:0] addr_47_4;

Selector_2 s47_4(wires_11_3[3], addr_11_3, wires_47_4,addr_47_4);

wire[3:0] wires_48_4;

wire[31:0] addr_48_4;

Selector_2 s48_4(wires_12_3[0], addr_12_3, wires_48_4,addr_48_4);

wire[3:0] wires_49_4;

wire[31:0] addr_49_4;

Selector_2 s49_4(wires_12_3[1], addr_12_3, wires_49_4,addr_49_4);

wire[3:0] wires_50_4;

wire[31:0] addr_50_4;

Selector_2 s50_4(wires_12_3[2], addr_12_3, wires_50_4,addr_50_4);

wire[3:0] wires_51_4;

wire[31:0] addr_51_4;

Selector_2 s51_4(wires_12_3[3], addr_12_3, wires_51_4,addr_51_4);

wire[3:0] wires_52_4;

wire[31:0] addr_52_4;

Selector_2 s52_4(wires_13_3[0], addr_13_3, wires_52_4,addr_52_4);

wire[3:0] wires_53_4;

wire[31:0] addr_53_4;

Selector_2 s53_4(wires_13_3[1], addr_13_3, wires_53_4,addr_53_4);

wire[3:0] wires_54_4;

wire[31:0] addr_54_4;

Selector_2 s54_4(wires_13_3[2], addr_13_3, wires_54_4,addr_54_4);

wire[3:0] wires_55_4;

wire[31:0] addr_55_4;

Selector_2 s55_4(wires_13_3[3], addr_13_3, wires_55_4,addr_55_4);

wire[3:0] wires_56_4;

wire[31:0] addr_56_4;

Selector_2 s56_4(wires_14_3[0], addr_14_3, wires_56_4,addr_56_4);

wire[3:0] wires_57_4;

wire[31:0] addr_57_4;

Selector_2 s57_4(wires_14_3[1], addr_14_3, wires_57_4,addr_57_4);

wire[3:0] wires_58_4;

wire[31:0] addr_58_4;

Selector_2 s58_4(wires_14_3[2], addr_14_3, wires_58_4,addr_58_4);

wire[3:0] wires_59_4;

wire[31:0] addr_59_4;

Selector_2 s59_4(wires_14_3[3], addr_14_3, wires_59_4,addr_59_4);

wire[3:0] wires_60_4;

wire[31:0] addr_60_4;

Selector_2 s60_4(wires_15_3[0], addr_15_3, wires_60_4,addr_60_4);

wire[3:0] wires_61_4;

wire[31:0] addr_61_4;

Selector_2 s61_4(wires_15_3[1], addr_15_3, wires_61_4,addr_61_4);

wire[3:0] wires_62_4;

wire[31:0] addr_62_4;

Selector_2 s62_4(wires_15_3[2], addr_15_3, wires_62_4,addr_62_4);

wire[3:0] wires_63_4;

wire[31:0] addr_63_4;

Selector_2 s63_4(wires_15_3[3], addr_15_3, wires_63_4,addr_63_4);

wire[3:0] wires_64_4;

wire[31:0] addr_64_4;

Selector_2 s64_4(wires_16_3[0], addr_16_3, wires_64_4,addr_64_4);

wire[3:0] wires_65_4;

wire[31:0] addr_65_4;

Selector_2 s65_4(wires_16_3[1], addr_16_3, wires_65_4,addr_65_4);

wire[3:0] wires_66_4;

wire[31:0] addr_66_4;

Selector_2 s66_4(wires_16_3[2], addr_16_3, wires_66_4,addr_66_4);

wire[3:0] wires_67_4;

wire[31:0] addr_67_4;

Selector_2 s67_4(wires_16_3[3], addr_16_3, wires_67_4,addr_67_4);

wire[3:0] wires_68_4;

wire[31:0] addr_68_4;

Selector_2 s68_4(wires_17_3[0], addr_17_3, wires_68_4,addr_68_4);

wire[3:0] wires_69_4;

wire[31:0] addr_69_4;

Selector_2 s69_4(wires_17_3[1], addr_17_3, wires_69_4,addr_69_4);

wire[3:0] wires_70_4;

wire[31:0] addr_70_4;

Selector_2 s70_4(wires_17_3[2], addr_17_3, wires_70_4,addr_70_4);

wire[3:0] wires_71_4;

wire[31:0] addr_71_4;

Selector_2 s71_4(wires_17_3[3], addr_17_3, wires_71_4,addr_71_4);

wire[3:0] wires_72_4;

wire[31:0] addr_72_4;

Selector_2 s72_4(wires_18_3[0], addr_18_3, wires_72_4,addr_72_4);

wire[3:0] wires_73_4;

wire[31:0] addr_73_4;

Selector_2 s73_4(wires_18_3[1], addr_18_3, wires_73_4,addr_73_4);

wire[3:0] wires_74_4;

wire[31:0] addr_74_4;

Selector_2 s74_4(wires_18_3[2], addr_18_3, wires_74_4,addr_74_4);

wire[3:0] wires_75_4;

wire[31:0] addr_75_4;

Selector_2 s75_4(wires_18_3[3], addr_18_3, wires_75_4,addr_75_4);

wire[3:0] wires_76_4;

wire[31:0] addr_76_4;

Selector_2 s76_4(wires_19_3[0], addr_19_3, wires_76_4,addr_76_4);

wire[3:0] wires_77_4;

wire[31:0] addr_77_4;

Selector_2 s77_4(wires_19_3[1], addr_19_3, wires_77_4,addr_77_4);

wire[3:0] wires_78_4;

wire[31:0] addr_78_4;

Selector_2 s78_4(wires_19_3[2], addr_19_3, wires_78_4,addr_78_4);

wire[3:0] wires_79_4;

wire[31:0] addr_79_4;

Selector_2 s79_4(wires_19_3[3], addr_19_3, wires_79_4,addr_79_4);

wire[3:0] wires_80_4;

wire[31:0] addr_80_4;

Selector_2 s80_4(wires_20_3[0], addr_20_3, wires_80_4,addr_80_4);

wire[3:0] wires_81_4;

wire[31:0] addr_81_4;

Selector_2 s81_4(wires_20_3[1], addr_20_3, wires_81_4,addr_81_4);

wire[3:0] wires_82_4;

wire[31:0] addr_82_4;

Selector_2 s82_4(wires_20_3[2], addr_20_3, wires_82_4,addr_82_4);

wire[3:0] wires_83_4;

wire[31:0] addr_83_4;

Selector_2 s83_4(wires_20_3[3], addr_20_3, wires_83_4,addr_83_4);

wire[3:0] wires_84_4;

wire[31:0] addr_84_4;

Selector_2 s84_4(wires_21_3[0], addr_21_3, wires_84_4,addr_84_4);

wire[3:0] wires_85_4;

wire[31:0] addr_85_4;

Selector_2 s85_4(wires_21_3[1], addr_21_3, wires_85_4,addr_85_4);

wire[3:0] wires_86_4;

wire[31:0] addr_86_4;

Selector_2 s86_4(wires_21_3[2], addr_21_3, wires_86_4,addr_86_4);

wire[3:0] wires_87_4;

wire[31:0] addr_87_4;

Selector_2 s87_4(wires_21_3[3], addr_21_3, wires_87_4,addr_87_4);

wire[3:0] wires_88_4;

wire[31:0] addr_88_4;

Selector_2 s88_4(wires_22_3[0], addr_22_3, wires_88_4,addr_88_4);

wire[3:0] wires_89_4;

wire[31:0] addr_89_4;

Selector_2 s89_4(wires_22_3[1], addr_22_3, wires_89_4,addr_89_4);

wire[3:0] wires_90_4;

wire[31:0] addr_90_4;

Selector_2 s90_4(wires_22_3[2], addr_22_3, wires_90_4,addr_90_4);

wire[3:0] wires_91_4;

wire[31:0] addr_91_4;

Selector_2 s91_4(wires_22_3[3], addr_22_3, wires_91_4,addr_91_4);

wire[3:0] wires_92_4;

wire[31:0] addr_92_4;

Selector_2 s92_4(wires_23_3[0], addr_23_3, wires_92_4,addr_92_4);

wire[3:0] wires_93_4;

wire[31:0] addr_93_4;

Selector_2 s93_4(wires_23_3[1], addr_23_3, wires_93_4,addr_93_4);

wire[3:0] wires_94_4;

wire[31:0] addr_94_4;

Selector_2 s94_4(wires_23_3[2], addr_23_3, wires_94_4,addr_94_4);

wire[3:0] wires_95_4;

wire[31:0] addr_95_4;

Selector_2 s95_4(wires_23_3[3], addr_23_3, wires_95_4,addr_95_4);

wire[3:0] wires_96_4;

wire[31:0] addr_96_4;

Selector_2 s96_4(wires_24_3[0], addr_24_3, wires_96_4,addr_96_4);

wire[3:0] wires_97_4;

wire[31:0] addr_97_4;

Selector_2 s97_4(wires_24_3[1], addr_24_3, wires_97_4,addr_97_4);

wire[3:0] wires_98_4;

wire[31:0] addr_98_4;

Selector_2 s98_4(wires_24_3[2], addr_24_3, wires_98_4,addr_98_4);

wire[3:0] wires_99_4;

wire[31:0] addr_99_4;

Selector_2 s99_4(wires_24_3[3], addr_24_3, wires_99_4,addr_99_4);

wire[3:0] wires_100_4;

wire[31:0] addr_100_4;

Selector_2 s100_4(wires_25_3[0], addr_25_3, wires_100_4,addr_100_4);

wire[3:0] wires_101_4;

wire[31:0] addr_101_4;

Selector_2 s101_4(wires_25_3[1], addr_25_3, wires_101_4,addr_101_4);

wire[3:0] wires_102_4;

wire[31:0] addr_102_4;

Selector_2 s102_4(wires_25_3[2], addr_25_3, wires_102_4,addr_102_4);

wire[3:0] wires_103_4;

wire[31:0] addr_103_4;

Selector_2 s103_4(wires_25_3[3], addr_25_3, wires_103_4,addr_103_4);

wire[3:0] wires_104_4;

wire[31:0] addr_104_4;

Selector_2 s104_4(wires_26_3[0], addr_26_3, wires_104_4,addr_104_4);

wire[3:0] wires_105_4;

wire[31:0] addr_105_4;

Selector_2 s105_4(wires_26_3[1], addr_26_3, wires_105_4,addr_105_4);

wire[3:0] wires_106_4;

wire[31:0] addr_106_4;

Selector_2 s106_4(wires_26_3[2], addr_26_3, wires_106_4,addr_106_4);

wire[3:0] wires_107_4;

wire[31:0] addr_107_4;

Selector_2 s107_4(wires_26_3[3], addr_26_3, wires_107_4,addr_107_4);

wire[3:0] wires_108_4;

wire[31:0] addr_108_4;

Selector_2 s108_4(wires_27_3[0], addr_27_3, wires_108_4,addr_108_4);

wire[3:0] wires_109_4;

wire[31:0] addr_109_4;

Selector_2 s109_4(wires_27_3[1], addr_27_3, wires_109_4,addr_109_4);

wire[3:0] wires_110_4;

wire[31:0] addr_110_4;

Selector_2 s110_4(wires_27_3[2], addr_27_3, wires_110_4,addr_110_4);

wire[3:0] wires_111_4;

wire[31:0] addr_111_4;

Selector_2 s111_4(wires_27_3[3], addr_27_3, wires_111_4,addr_111_4);

wire[3:0] wires_112_4;

wire[31:0] addr_112_4;

Selector_2 s112_4(wires_28_3[0], addr_28_3, wires_112_4,addr_112_4);

wire[3:0] wires_113_4;

wire[31:0] addr_113_4;

Selector_2 s113_4(wires_28_3[1], addr_28_3, wires_113_4,addr_113_4);

wire[3:0] wires_114_4;

wire[31:0] addr_114_4;

Selector_2 s114_4(wires_28_3[2], addr_28_3, wires_114_4,addr_114_4);

wire[3:0] wires_115_4;

wire[31:0] addr_115_4;

Selector_2 s115_4(wires_28_3[3], addr_28_3, wires_115_4,addr_115_4);

wire[3:0] wires_116_4;

wire[31:0] addr_116_4;

Selector_2 s116_4(wires_29_3[0], addr_29_3, wires_116_4,addr_116_4);

wire[3:0] wires_117_4;

wire[31:0] addr_117_4;

Selector_2 s117_4(wires_29_3[1], addr_29_3, wires_117_4,addr_117_4);

wire[3:0] wires_118_4;

wire[31:0] addr_118_4;

Selector_2 s118_4(wires_29_3[2], addr_29_3, wires_118_4,addr_118_4);

wire[3:0] wires_119_4;

wire[31:0] addr_119_4;

Selector_2 s119_4(wires_29_3[3], addr_29_3, wires_119_4,addr_119_4);

wire[3:0] wires_120_4;

wire[31:0] addr_120_4;

Selector_2 s120_4(wires_30_3[0], addr_30_3, wires_120_4,addr_120_4);

wire[3:0] wires_121_4;

wire[31:0] addr_121_4;

Selector_2 s121_4(wires_30_3[1], addr_30_3, wires_121_4,addr_121_4);

wire[3:0] wires_122_4;

wire[31:0] addr_122_4;

Selector_2 s122_4(wires_30_3[2], addr_30_3, wires_122_4,addr_122_4);

wire[3:0] wires_123_4;

wire[31:0] addr_123_4;

Selector_2 s123_4(wires_30_3[3], addr_30_3, wires_123_4,addr_123_4);

wire[3:0] wires_124_4;

wire[31:0] addr_124_4;

Selector_2 s124_4(wires_31_3[0], addr_31_3, wires_124_4,addr_124_4);

wire[3:0] wires_125_4;

wire[31:0] addr_125_4;

Selector_2 s125_4(wires_31_3[1], addr_31_3, wires_125_4,addr_125_4);

wire[3:0] wires_126_4;

wire[31:0] addr_126_4;

Selector_2 s126_4(wires_31_3[2], addr_31_3, wires_126_4,addr_126_4);

wire[3:0] wires_127_4;

wire[31:0] addr_127_4;

Selector_2 s127_4(wires_31_3[3], addr_31_3, wires_127_4,addr_127_4);

wire[3:0] wires_128_4;

wire[31:0] addr_128_4;

Selector_2 s128_4(wires_32_3[0], addr_32_3, wires_128_4,addr_128_4);

wire[3:0] wires_129_4;

wire[31:0] addr_129_4;

Selector_2 s129_4(wires_32_3[1], addr_32_3, wires_129_4,addr_129_4);

wire[3:0] wires_130_4;

wire[31:0] addr_130_4;

Selector_2 s130_4(wires_32_3[2], addr_32_3, wires_130_4,addr_130_4);

wire[3:0] wires_131_4;

wire[31:0] addr_131_4;

Selector_2 s131_4(wires_32_3[3], addr_32_3, wires_131_4,addr_131_4);

wire[3:0] wires_132_4;

wire[31:0] addr_132_4;

Selector_2 s132_4(wires_33_3[0], addr_33_3, wires_132_4,addr_132_4);

wire[3:0] wires_133_4;

wire[31:0] addr_133_4;

Selector_2 s133_4(wires_33_3[1], addr_33_3, wires_133_4,addr_133_4);

wire[3:0] wires_134_4;

wire[31:0] addr_134_4;

Selector_2 s134_4(wires_33_3[2], addr_33_3, wires_134_4,addr_134_4);

wire[3:0] wires_135_4;

wire[31:0] addr_135_4;

Selector_2 s135_4(wires_33_3[3], addr_33_3, wires_135_4,addr_135_4);

wire[3:0] wires_136_4;

wire[31:0] addr_136_4;

Selector_2 s136_4(wires_34_3[0], addr_34_3, wires_136_4,addr_136_4);

wire[3:0] wires_137_4;

wire[31:0] addr_137_4;

Selector_2 s137_4(wires_34_3[1], addr_34_3, wires_137_4,addr_137_4);

wire[3:0] wires_138_4;

wire[31:0] addr_138_4;

Selector_2 s138_4(wires_34_3[2], addr_34_3, wires_138_4,addr_138_4);

wire[3:0] wires_139_4;

wire[31:0] addr_139_4;

Selector_2 s139_4(wires_34_3[3], addr_34_3, wires_139_4,addr_139_4);

wire[3:0] wires_140_4;

wire[31:0] addr_140_4;

Selector_2 s140_4(wires_35_3[0], addr_35_3, wires_140_4,addr_140_4);

wire[3:0] wires_141_4;

wire[31:0] addr_141_4;

Selector_2 s141_4(wires_35_3[1], addr_35_3, wires_141_4,addr_141_4);

wire[3:0] wires_142_4;

wire[31:0] addr_142_4;

Selector_2 s142_4(wires_35_3[2], addr_35_3, wires_142_4,addr_142_4);

wire[3:0] wires_143_4;

wire[31:0] addr_143_4;

Selector_2 s143_4(wires_35_3[3], addr_35_3, wires_143_4,addr_143_4);

wire[3:0] wires_144_4;

wire[31:0] addr_144_4;

Selector_2 s144_4(wires_36_3[0], addr_36_3, wires_144_4,addr_144_4);

wire[3:0] wires_145_4;

wire[31:0] addr_145_4;

Selector_2 s145_4(wires_36_3[1], addr_36_3, wires_145_4,addr_145_4);

wire[3:0] wires_146_4;

wire[31:0] addr_146_4;

Selector_2 s146_4(wires_36_3[2], addr_36_3, wires_146_4,addr_146_4);

wire[3:0] wires_147_4;

wire[31:0] addr_147_4;

Selector_2 s147_4(wires_36_3[3], addr_36_3, wires_147_4,addr_147_4);

wire[3:0] wires_148_4;

wire[31:0] addr_148_4;

Selector_2 s148_4(wires_37_3[0], addr_37_3, wires_148_4,addr_148_4);

wire[3:0] wires_149_4;

wire[31:0] addr_149_4;

Selector_2 s149_4(wires_37_3[1], addr_37_3, wires_149_4,addr_149_4);

wire[3:0] wires_150_4;

wire[31:0] addr_150_4;

Selector_2 s150_4(wires_37_3[2], addr_37_3, wires_150_4,addr_150_4);

wire[3:0] wires_151_4;

wire[31:0] addr_151_4;

Selector_2 s151_4(wires_37_3[3], addr_37_3, wires_151_4,addr_151_4);

wire[3:0] wires_152_4;

wire[31:0] addr_152_4;

Selector_2 s152_4(wires_38_3[0], addr_38_3, wires_152_4,addr_152_4);

wire[3:0] wires_153_4;

wire[31:0] addr_153_4;

Selector_2 s153_4(wires_38_3[1], addr_38_3, wires_153_4,addr_153_4);

wire[3:0] wires_154_4;

wire[31:0] addr_154_4;

Selector_2 s154_4(wires_38_3[2], addr_38_3, wires_154_4,addr_154_4);

wire[3:0] wires_155_4;

wire[31:0] addr_155_4;

Selector_2 s155_4(wires_38_3[3], addr_38_3, wires_155_4,addr_155_4);

wire[3:0] wires_156_4;

wire[31:0] addr_156_4;

Selector_2 s156_4(wires_39_3[0], addr_39_3, wires_156_4,addr_156_4);

wire[3:0] wires_157_4;

wire[31:0] addr_157_4;

Selector_2 s157_4(wires_39_3[1], addr_39_3, wires_157_4,addr_157_4);

wire[3:0] wires_158_4;

wire[31:0] addr_158_4;

Selector_2 s158_4(wires_39_3[2], addr_39_3, wires_158_4,addr_158_4);

wire[3:0] wires_159_4;

wire[31:0] addr_159_4;

Selector_2 s159_4(wires_39_3[3], addr_39_3, wires_159_4,addr_159_4);

wire[3:0] wires_160_4;

wire[31:0] addr_160_4;

Selector_2 s160_4(wires_40_3[0], addr_40_3, wires_160_4,addr_160_4);

wire[3:0] wires_161_4;

wire[31:0] addr_161_4;

Selector_2 s161_4(wires_40_3[1], addr_40_3, wires_161_4,addr_161_4);

wire[3:0] wires_162_4;

wire[31:0] addr_162_4;

Selector_2 s162_4(wires_40_3[2], addr_40_3, wires_162_4,addr_162_4);

wire[3:0] wires_163_4;

wire[31:0] addr_163_4;

Selector_2 s163_4(wires_40_3[3], addr_40_3, wires_163_4,addr_163_4);

wire[3:0] wires_164_4;

wire[31:0] addr_164_4;

Selector_2 s164_4(wires_41_3[0], addr_41_3, wires_164_4,addr_164_4);

wire[3:0] wires_165_4;

wire[31:0] addr_165_4;

Selector_2 s165_4(wires_41_3[1], addr_41_3, wires_165_4,addr_165_4);

wire[3:0] wires_166_4;

wire[31:0] addr_166_4;

Selector_2 s166_4(wires_41_3[2], addr_41_3, wires_166_4,addr_166_4);

wire[3:0] wires_167_4;

wire[31:0] addr_167_4;

Selector_2 s167_4(wires_41_3[3], addr_41_3, wires_167_4,addr_167_4);

wire[3:0] wires_168_4;

wire[31:0] addr_168_4;

Selector_2 s168_4(wires_42_3[0], addr_42_3, wires_168_4,addr_168_4);

wire[3:0] wires_169_4;

wire[31:0] addr_169_4;

Selector_2 s169_4(wires_42_3[1], addr_42_3, wires_169_4,addr_169_4);

wire[3:0] wires_170_4;

wire[31:0] addr_170_4;

Selector_2 s170_4(wires_42_3[2], addr_42_3, wires_170_4,addr_170_4);

wire[3:0] wires_171_4;

wire[31:0] addr_171_4;

Selector_2 s171_4(wires_42_3[3], addr_42_3, wires_171_4,addr_171_4);

wire[3:0] wires_172_4;

wire[31:0] addr_172_4;

Selector_2 s172_4(wires_43_3[0], addr_43_3, wires_172_4,addr_172_4);

wire[3:0] wires_173_4;

wire[31:0] addr_173_4;

Selector_2 s173_4(wires_43_3[1], addr_43_3, wires_173_4,addr_173_4);

wire[3:0] wires_174_4;

wire[31:0] addr_174_4;

Selector_2 s174_4(wires_43_3[2], addr_43_3, wires_174_4,addr_174_4);

wire[3:0] wires_175_4;

wire[31:0] addr_175_4;

Selector_2 s175_4(wires_43_3[3], addr_43_3, wires_175_4,addr_175_4);

wire[3:0] wires_176_4;

wire[31:0] addr_176_4;

Selector_2 s176_4(wires_44_3[0], addr_44_3, wires_176_4,addr_176_4);

wire[3:0] wires_177_4;

wire[31:0] addr_177_4;

Selector_2 s177_4(wires_44_3[1], addr_44_3, wires_177_4,addr_177_4);

wire[3:0] wires_178_4;

wire[31:0] addr_178_4;

Selector_2 s178_4(wires_44_3[2], addr_44_3, wires_178_4,addr_178_4);

wire[3:0] wires_179_4;

wire[31:0] addr_179_4;

Selector_2 s179_4(wires_44_3[3], addr_44_3, wires_179_4,addr_179_4);

wire[3:0] wires_180_4;

wire[31:0] addr_180_4;

Selector_2 s180_4(wires_45_3[0], addr_45_3, wires_180_4,addr_180_4);

wire[3:0] wires_181_4;

wire[31:0] addr_181_4;

Selector_2 s181_4(wires_45_3[1], addr_45_3, wires_181_4,addr_181_4);

wire[3:0] wires_182_4;

wire[31:0] addr_182_4;

Selector_2 s182_4(wires_45_3[2], addr_45_3, wires_182_4,addr_182_4);

wire[3:0] wires_183_4;

wire[31:0] addr_183_4;

Selector_2 s183_4(wires_45_3[3], addr_45_3, wires_183_4,addr_183_4);

wire[3:0] wires_184_4;

wire[31:0] addr_184_4;

Selector_2 s184_4(wires_46_3[0], addr_46_3, wires_184_4,addr_184_4);

wire[3:0] wires_185_4;

wire[31:0] addr_185_4;

Selector_2 s185_4(wires_46_3[1], addr_46_3, wires_185_4,addr_185_4);

wire[3:0] wires_186_4;

wire[31:0] addr_186_4;

Selector_2 s186_4(wires_46_3[2], addr_46_3, wires_186_4,addr_186_4);

wire[3:0] wires_187_4;

wire[31:0] addr_187_4;

Selector_2 s187_4(wires_46_3[3], addr_46_3, wires_187_4,addr_187_4);

wire[3:0] wires_188_4;

wire[31:0] addr_188_4;

Selector_2 s188_4(wires_47_3[0], addr_47_3, wires_188_4,addr_188_4);

wire[3:0] wires_189_4;

wire[31:0] addr_189_4;

Selector_2 s189_4(wires_47_3[1], addr_47_3, wires_189_4,addr_189_4);

wire[3:0] wires_190_4;

wire[31:0] addr_190_4;

Selector_2 s190_4(wires_47_3[2], addr_47_3, wires_190_4,addr_190_4);

wire[3:0] wires_191_4;

wire[31:0] addr_191_4;

Selector_2 s191_4(wires_47_3[3], addr_47_3, wires_191_4,addr_191_4);

wire[3:0] wires_192_4;

wire[31:0] addr_192_4;

Selector_2 s192_4(wires_48_3[0], addr_48_3, wires_192_4,addr_192_4);

wire[3:0] wires_193_4;

wire[31:0] addr_193_4;

Selector_2 s193_4(wires_48_3[1], addr_48_3, wires_193_4,addr_193_4);

wire[3:0] wires_194_4;

wire[31:0] addr_194_4;

Selector_2 s194_4(wires_48_3[2], addr_48_3, wires_194_4,addr_194_4);

wire[3:0] wires_195_4;

wire[31:0] addr_195_4;

Selector_2 s195_4(wires_48_3[3], addr_48_3, wires_195_4,addr_195_4);

wire[3:0] wires_196_4;

wire[31:0] addr_196_4;

Selector_2 s196_4(wires_49_3[0], addr_49_3, wires_196_4,addr_196_4);

wire[3:0] wires_197_4;

wire[31:0] addr_197_4;

Selector_2 s197_4(wires_49_3[1], addr_49_3, wires_197_4,addr_197_4);

wire[3:0] wires_198_4;

wire[31:0] addr_198_4;

Selector_2 s198_4(wires_49_3[2], addr_49_3, wires_198_4,addr_198_4);

wire[3:0] wires_199_4;

wire[31:0] addr_199_4;

Selector_2 s199_4(wires_49_3[3], addr_49_3, wires_199_4,addr_199_4);

wire[3:0] wires_200_4;

wire[31:0] addr_200_4;

Selector_2 s200_4(wires_50_3[0], addr_50_3, wires_200_4,addr_200_4);

wire[3:0] wires_201_4;

wire[31:0] addr_201_4;

Selector_2 s201_4(wires_50_3[1], addr_50_3, wires_201_4,addr_201_4);

wire[3:0] wires_202_4;

wire[31:0] addr_202_4;

Selector_2 s202_4(wires_50_3[2], addr_50_3, wires_202_4,addr_202_4);

wire[3:0] wires_203_4;

wire[31:0] addr_203_4;

Selector_2 s203_4(wires_50_3[3], addr_50_3, wires_203_4,addr_203_4);

wire[3:0] wires_204_4;

wire[31:0] addr_204_4;

Selector_2 s204_4(wires_51_3[0], addr_51_3, wires_204_4,addr_204_4);

wire[3:0] wires_205_4;

wire[31:0] addr_205_4;

Selector_2 s205_4(wires_51_3[1], addr_51_3, wires_205_4,addr_205_4);

wire[3:0] wires_206_4;

wire[31:0] addr_206_4;

Selector_2 s206_4(wires_51_3[2], addr_51_3, wires_206_4,addr_206_4);

wire[3:0] wires_207_4;

wire[31:0] addr_207_4;

Selector_2 s207_4(wires_51_3[3], addr_51_3, wires_207_4,addr_207_4);

wire[3:0] wires_208_4;

wire[31:0] addr_208_4;

Selector_2 s208_4(wires_52_3[0], addr_52_3, wires_208_4,addr_208_4);

wire[3:0] wires_209_4;

wire[31:0] addr_209_4;

Selector_2 s209_4(wires_52_3[1], addr_52_3, wires_209_4,addr_209_4);

wire[3:0] wires_210_4;

wire[31:0] addr_210_4;

Selector_2 s210_4(wires_52_3[2], addr_52_3, wires_210_4,addr_210_4);

wire[3:0] wires_211_4;

wire[31:0] addr_211_4;

Selector_2 s211_4(wires_52_3[3], addr_52_3, wires_211_4,addr_211_4);

wire[3:0] wires_212_4;

wire[31:0] addr_212_4;

Selector_2 s212_4(wires_53_3[0], addr_53_3, wires_212_4,addr_212_4);

wire[3:0] wires_213_4;

wire[31:0] addr_213_4;

Selector_2 s213_4(wires_53_3[1], addr_53_3, wires_213_4,addr_213_4);

wire[3:0] wires_214_4;

wire[31:0] addr_214_4;

Selector_2 s214_4(wires_53_3[2], addr_53_3, wires_214_4,addr_214_4);

wire[3:0] wires_215_4;

wire[31:0] addr_215_4;

Selector_2 s215_4(wires_53_3[3], addr_53_3, wires_215_4,addr_215_4);

wire[3:0] wires_216_4;

wire[31:0] addr_216_4;

Selector_2 s216_4(wires_54_3[0], addr_54_3, wires_216_4,addr_216_4);

wire[3:0] wires_217_4;

wire[31:0] addr_217_4;

Selector_2 s217_4(wires_54_3[1], addr_54_3, wires_217_4,addr_217_4);

wire[3:0] wires_218_4;

wire[31:0] addr_218_4;

Selector_2 s218_4(wires_54_3[2], addr_54_3, wires_218_4,addr_218_4);

wire[3:0] wires_219_4;

wire[31:0] addr_219_4;

Selector_2 s219_4(wires_54_3[3], addr_54_3, wires_219_4,addr_219_4);

wire[3:0] wires_220_4;

wire[31:0] addr_220_4;

Selector_2 s220_4(wires_55_3[0], addr_55_3, wires_220_4,addr_220_4);

wire[3:0] wires_221_4;

wire[31:0] addr_221_4;

Selector_2 s221_4(wires_55_3[1], addr_55_3, wires_221_4,addr_221_4);

wire[3:0] wires_222_4;

wire[31:0] addr_222_4;

Selector_2 s222_4(wires_55_3[2], addr_55_3, wires_222_4,addr_222_4);

wire[3:0] wires_223_4;

wire[31:0] addr_223_4;

Selector_2 s223_4(wires_55_3[3], addr_55_3, wires_223_4,addr_223_4);

wire[3:0] wires_224_4;

wire[31:0] addr_224_4;

Selector_2 s224_4(wires_56_3[0], addr_56_3, wires_224_4,addr_224_4);

wire[3:0] wires_225_4;

wire[31:0] addr_225_4;

Selector_2 s225_4(wires_56_3[1], addr_56_3, wires_225_4,addr_225_4);

wire[3:0] wires_226_4;

wire[31:0] addr_226_4;

Selector_2 s226_4(wires_56_3[2], addr_56_3, wires_226_4,addr_226_4);

wire[3:0] wires_227_4;

wire[31:0] addr_227_4;

Selector_2 s227_4(wires_56_3[3], addr_56_3, wires_227_4,addr_227_4);

wire[3:0] wires_228_4;

wire[31:0] addr_228_4;

Selector_2 s228_4(wires_57_3[0], addr_57_3, wires_228_4,addr_228_4);

wire[3:0] wires_229_4;

wire[31:0] addr_229_4;

Selector_2 s229_4(wires_57_3[1], addr_57_3, wires_229_4,addr_229_4);

wire[3:0] wires_230_4;

wire[31:0] addr_230_4;

Selector_2 s230_4(wires_57_3[2], addr_57_3, wires_230_4,addr_230_4);

wire[3:0] wires_231_4;

wire[31:0] addr_231_4;

Selector_2 s231_4(wires_57_3[3], addr_57_3, wires_231_4,addr_231_4);

wire[3:0] wires_232_4;

wire[31:0] addr_232_4;

Selector_2 s232_4(wires_58_3[0], addr_58_3, wires_232_4,addr_232_4);

wire[3:0] wires_233_4;

wire[31:0] addr_233_4;

Selector_2 s233_4(wires_58_3[1], addr_58_3, wires_233_4,addr_233_4);

wire[3:0] wires_234_4;

wire[31:0] addr_234_4;

Selector_2 s234_4(wires_58_3[2], addr_58_3, wires_234_4,addr_234_4);

wire[3:0] wires_235_4;

wire[31:0] addr_235_4;

Selector_2 s235_4(wires_58_3[3], addr_58_3, wires_235_4,addr_235_4);

wire[3:0] wires_236_4;

wire[31:0] addr_236_4;

Selector_2 s236_4(wires_59_3[0], addr_59_3, wires_236_4,addr_236_4);

wire[3:0] wires_237_4;

wire[31:0] addr_237_4;

Selector_2 s237_4(wires_59_3[1], addr_59_3, wires_237_4,addr_237_4);

wire[3:0] wires_238_4;

wire[31:0] addr_238_4;

Selector_2 s238_4(wires_59_3[2], addr_59_3, wires_238_4,addr_238_4);

wire[3:0] wires_239_4;

wire[31:0] addr_239_4;

Selector_2 s239_4(wires_59_3[3], addr_59_3, wires_239_4,addr_239_4);

wire[3:0] wires_240_4;

wire[31:0] addr_240_4;

Selector_2 s240_4(wires_60_3[0], addr_60_3, wires_240_4,addr_240_4);

wire[3:0] wires_241_4;

wire[31:0] addr_241_4;

Selector_2 s241_4(wires_60_3[1], addr_60_3, wires_241_4,addr_241_4);

wire[3:0] wires_242_4;

wire[31:0] addr_242_4;

Selector_2 s242_4(wires_60_3[2], addr_60_3, wires_242_4,addr_242_4);

wire[3:0] wires_243_4;

wire[31:0] addr_243_4;

Selector_2 s243_4(wires_60_3[3], addr_60_3, wires_243_4,addr_243_4);

wire[3:0] wires_244_4;

wire[31:0] addr_244_4;

Selector_2 s244_4(wires_61_3[0], addr_61_3, wires_244_4,addr_244_4);

wire[3:0] wires_245_4;

wire[31:0] addr_245_4;

Selector_2 s245_4(wires_61_3[1], addr_61_3, wires_245_4,addr_245_4);

wire[3:0] wires_246_4;

wire[31:0] addr_246_4;

Selector_2 s246_4(wires_61_3[2], addr_61_3, wires_246_4,addr_246_4);

wire[3:0] wires_247_4;

wire[31:0] addr_247_4;

Selector_2 s247_4(wires_61_3[3], addr_61_3, wires_247_4,addr_247_4);

wire[3:0] wires_248_4;

wire[31:0] addr_248_4;

Selector_2 s248_4(wires_62_3[0], addr_62_3, wires_248_4,addr_248_4);

wire[3:0] wires_249_4;

wire[31:0] addr_249_4;

Selector_2 s249_4(wires_62_3[1], addr_62_3, wires_249_4,addr_249_4);

wire[3:0] wires_250_4;

wire[31:0] addr_250_4;

Selector_2 s250_4(wires_62_3[2], addr_62_3, wires_250_4,addr_250_4);

wire[3:0] wires_251_4;

wire[31:0] addr_251_4;

Selector_2 s251_4(wires_62_3[3], addr_62_3, wires_251_4,addr_251_4);

wire[3:0] wires_252_4;

wire[31:0] addr_252_4;

Selector_2 s252_4(wires_63_3[0], addr_63_3, wires_252_4,addr_252_4);

wire[3:0] wires_253_4;

wire[31:0] addr_253_4;

Selector_2 s253_4(wires_63_3[1], addr_63_3, wires_253_4,addr_253_4);

wire[3:0] wires_254_4;

wire[31:0] addr_254_4;

Selector_2 s254_4(wires_63_3[2], addr_63_3, wires_254_4,addr_254_4);

wire[3:0] wires_255_4;

wire[31:0] addr_255_4;

Selector_2 s255_4(wires_63_3[3], addr_63_3, wires_255_4,addr_255_4);

wire[3:0] wires_0_5;

wire[31:0] addr_0_5;

Selector_2 s0_5(wires_0_4[0], addr_0_4, wires_0_5,addr_0_5);

wire[3:0] wires_1_5;

wire[31:0] addr_1_5;

Selector_2 s1_5(wires_0_4[1], addr_0_4, wires_1_5,addr_1_5);

wire[3:0] wires_2_5;

wire[31:0] addr_2_5;

Selector_2 s2_5(wires_0_4[2], addr_0_4, wires_2_5,addr_2_5);

wire[3:0] wires_3_5;

wire[31:0] addr_3_5;

Selector_2 s3_5(wires_0_4[3], addr_0_4, wires_3_5,addr_3_5);

wire[3:0] wires_4_5;

wire[31:0] addr_4_5;

Selector_2 s4_5(wires_1_4[0], addr_1_4, wires_4_5,addr_4_5);

wire[3:0] wires_5_5;

wire[31:0] addr_5_5;

Selector_2 s5_5(wires_1_4[1], addr_1_4, wires_5_5,addr_5_5);

wire[3:0] wires_6_5;

wire[31:0] addr_6_5;

Selector_2 s6_5(wires_1_4[2], addr_1_4, wires_6_5,addr_6_5);

wire[3:0] wires_7_5;

wire[31:0] addr_7_5;

Selector_2 s7_5(wires_1_4[3], addr_1_4, wires_7_5,addr_7_5);

wire[3:0] wires_8_5;

wire[31:0] addr_8_5;

Selector_2 s8_5(wires_2_4[0], addr_2_4, wires_8_5,addr_8_5);

wire[3:0] wires_9_5;

wire[31:0] addr_9_5;

Selector_2 s9_5(wires_2_4[1], addr_2_4, wires_9_5,addr_9_5);

wire[3:0] wires_10_5;

wire[31:0] addr_10_5;

Selector_2 s10_5(wires_2_4[2], addr_2_4, wires_10_5,addr_10_5);

wire[3:0] wires_11_5;

wire[31:0] addr_11_5;

Selector_2 s11_5(wires_2_4[3], addr_2_4, wires_11_5,addr_11_5);

wire[3:0] wires_12_5;

wire[31:0] addr_12_5;

Selector_2 s12_5(wires_3_4[0], addr_3_4, wires_12_5,addr_12_5);

wire[3:0] wires_13_5;

wire[31:0] addr_13_5;

Selector_2 s13_5(wires_3_4[1], addr_3_4, wires_13_5,addr_13_5);

wire[3:0] wires_14_5;

wire[31:0] addr_14_5;

Selector_2 s14_5(wires_3_4[2], addr_3_4, wires_14_5,addr_14_5);

wire[3:0] wires_15_5;

wire[31:0] addr_15_5;

Selector_2 s15_5(wires_3_4[3], addr_3_4, wires_15_5,addr_15_5);

wire[3:0] wires_16_5;

wire[31:0] addr_16_5;

Selector_2 s16_5(wires_4_4[0], addr_4_4, wires_16_5,addr_16_5);

wire[3:0] wires_17_5;

wire[31:0] addr_17_5;

Selector_2 s17_5(wires_4_4[1], addr_4_4, wires_17_5,addr_17_5);

wire[3:0] wires_18_5;

wire[31:0] addr_18_5;

Selector_2 s18_5(wires_4_4[2], addr_4_4, wires_18_5,addr_18_5);

wire[3:0] wires_19_5;

wire[31:0] addr_19_5;

Selector_2 s19_5(wires_4_4[3], addr_4_4, wires_19_5,addr_19_5);

wire[3:0] wires_20_5;

wire[31:0] addr_20_5;

Selector_2 s20_5(wires_5_4[0], addr_5_4, wires_20_5,addr_20_5);

wire[3:0] wires_21_5;

wire[31:0] addr_21_5;

Selector_2 s21_5(wires_5_4[1], addr_5_4, wires_21_5,addr_21_5);

wire[3:0] wires_22_5;

wire[31:0] addr_22_5;

Selector_2 s22_5(wires_5_4[2], addr_5_4, wires_22_5,addr_22_5);

wire[3:0] wires_23_5;

wire[31:0] addr_23_5;

Selector_2 s23_5(wires_5_4[3], addr_5_4, wires_23_5,addr_23_5);

wire[3:0] wires_24_5;

wire[31:0] addr_24_5;

Selector_2 s24_5(wires_6_4[0], addr_6_4, wires_24_5,addr_24_5);

wire[3:0] wires_25_5;

wire[31:0] addr_25_5;

Selector_2 s25_5(wires_6_4[1], addr_6_4, wires_25_5,addr_25_5);

wire[3:0] wires_26_5;

wire[31:0] addr_26_5;

Selector_2 s26_5(wires_6_4[2], addr_6_4, wires_26_5,addr_26_5);

wire[3:0] wires_27_5;

wire[31:0] addr_27_5;

Selector_2 s27_5(wires_6_4[3], addr_6_4, wires_27_5,addr_27_5);

wire[3:0] wires_28_5;

wire[31:0] addr_28_5;

Selector_2 s28_5(wires_7_4[0], addr_7_4, wires_28_5,addr_28_5);

wire[3:0] wires_29_5;

wire[31:0] addr_29_5;

Selector_2 s29_5(wires_7_4[1], addr_7_4, wires_29_5,addr_29_5);

wire[3:0] wires_30_5;

wire[31:0] addr_30_5;

Selector_2 s30_5(wires_7_4[2], addr_7_4, wires_30_5,addr_30_5);

wire[3:0] wires_31_5;

wire[31:0] addr_31_5;

Selector_2 s31_5(wires_7_4[3], addr_7_4, wires_31_5,addr_31_5);

wire[3:0] wires_32_5;

wire[31:0] addr_32_5;

Selector_2 s32_5(wires_8_4[0], addr_8_4, wires_32_5,addr_32_5);

wire[3:0] wires_33_5;

wire[31:0] addr_33_5;

Selector_2 s33_5(wires_8_4[1], addr_8_4, wires_33_5,addr_33_5);

wire[3:0] wires_34_5;

wire[31:0] addr_34_5;

Selector_2 s34_5(wires_8_4[2], addr_8_4, wires_34_5,addr_34_5);

wire[3:0] wires_35_5;

wire[31:0] addr_35_5;

Selector_2 s35_5(wires_8_4[3], addr_8_4, wires_35_5,addr_35_5);

wire[3:0] wires_36_5;

wire[31:0] addr_36_5;

Selector_2 s36_5(wires_9_4[0], addr_9_4, wires_36_5,addr_36_5);

wire[3:0] wires_37_5;

wire[31:0] addr_37_5;

Selector_2 s37_5(wires_9_4[1], addr_9_4, wires_37_5,addr_37_5);

wire[3:0] wires_38_5;

wire[31:0] addr_38_5;

Selector_2 s38_5(wires_9_4[2], addr_9_4, wires_38_5,addr_38_5);

wire[3:0] wires_39_5;

wire[31:0] addr_39_5;

Selector_2 s39_5(wires_9_4[3], addr_9_4, wires_39_5,addr_39_5);

wire[3:0] wires_40_5;

wire[31:0] addr_40_5;

Selector_2 s40_5(wires_10_4[0], addr_10_4, wires_40_5,addr_40_5);

wire[3:0] wires_41_5;

wire[31:0] addr_41_5;

Selector_2 s41_5(wires_10_4[1], addr_10_4, wires_41_5,addr_41_5);

wire[3:0] wires_42_5;

wire[31:0] addr_42_5;

Selector_2 s42_5(wires_10_4[2], addr_10_4, wires_42_5,addr_42_5);

wire[3:0] wires_43_5;

wire[31:0] addr_43_5;

Selector_2 s43_5(wires_10_4[3], addr_10_4, wires_43_5,addr_43_5);

wire[3:0] wires_44_5;

wire[31:0] addr_44_5;

Selector_2 s44_5(wires_11_4[0], addr_11_4, wires_44_5,addr_44_5);

wire[3:0] wires_45_5;

wire[31:0] addr_45_5;

Selector_2 s45_5(wires_11_4[1], addr_11_4, wires_45_5,addr_45_5);

wire[3:0] wires_46_5;

wire[31:0] addr_46_5;

Selector_2 s46_5(wires_11_4[2], addr_11_4, wires_46_5,addr_46_5);

wire[3:0] wires_47_5;

wire[31:0] addr_47_5;

Selector_2 s47_5(wires_11_4[3], addr_11_4, wires_47_5,addr_47_5);

wire[3:0] wires_48_5;

wire[31:0] addr_48_5;

Selector_2 s48_5(wires_12_4[0], addr_12_4, wires_48_5,addr_48_5);

wire[3:0] wires_49_5;

wire[31:0] addr_49_5;

Selector_2 s49_5(wires_12_4[1], addr_12_4, wires_49_5,addr_49_5);

wire[3:0] wires_50_5;

wire[31:0] addr_50_5;

Selector_2 s50_5(wires_12_4[2], addr_12_4, wires_50_5,addr_50_5);

wire[3:0] wires_51_5;

wire[31:0] addr_51_5;

Selector_2 s51_5(wires_12_4[3], addr_12_4, wires_51_5,addr_51_5);

wire[3:0] wires_52_5;

wire[31:0] addr_52_5;

Selector_2 s52_5(wires_13_4[0], addr_13_4, wires_52_5,addr_52_5);

wire[3:0] wires_53_5;

wire[31:0] addr_53_5;

Selector_2 s53_5(wires_13_4[1], addr_13_4, wires_53_5,addr_53_5);

wire[3:0] wires_54_5;

wire[31:0] addr_54_5;

Selector_2 s54_5(wires_13_4[2], addr_13_4, wires_54_5,addr_54_5);

wire[3:0] wires_55_5;

wire[31:0] addr_55_5;

Selector_2 s55_5(wires_13_4[3], addr_13_4, wires_55_5,addr_55_5);

wire[3:0] wires_56_5;

wire[31:0] addr_56_5;

Selector_2 s56_5(wires_14_4[0], addr_14_4, wires_56_5,addr_56_5);

wire[3:0] wires_57_5;

wire[31:0] addr_57_5;

Selector_2 s57_5(wires_14_4[1], addr_14_4, wires_57_5,addr_57_5);

wire[3:0] wires_58_5;

wire[31:0] addr_58_5;

Selector_2 s58_5(wires_14_4[2], addr_14_4, wires_58_5,addr_58_5);

wire[3:0] wires_59_5;

wire[31:0] addr_59_5;

Selector_2 s59_5(wires_14_4[3], addr_14_4, wires_59_5,addr_59_5);

wire[3:0] wires_60_5;

wire[31:0] addr_60_5;

Selector_2 s60_5(wires_15_4[0], addr_15_4, wires_60_5,addr_60_5);

wire[3:0] wires_61_5;

wire[31:0] addr_61_5;

Selector_2 s61_5(wires_15_4[1], addr_15_4, wires_61_5,addr_61_5);

wire[3:0] wires_62_5;

wire[31:0] addr_62_5;

Selector_2 s62_5(wires_15_4[2], addr_15_4, wires_62_5,addr_62_5);

wire[3:0] wires_63_5;

wire[31:0] addr_63_5;

Selector_2 s63_5(wires_15_4[3], addr_15_4, wires_63_5,addr_63_5);

wire[3:0] wires_64_5;

wire[31:0] addr_64_5;

Selector_2 s64_5(wires_16_4[0], addr_16_4, wires_64_5,addr_64_5);

wire[3:0] wires_65_5;

wire[31:0] addr_65_5;

Selector_2 s65_5(wires_16_4[1], addr_16_4, wires_65_5,addr_65_5);

wire[3:0] wires_66_5;

wire[31:0] addr_66_5;

Selector_2 s66_5(wires_16_4[2], addr_16_4, wires_66_5,addr_66_5);

wire[3:0] wires_67_5;

wire[31:0] addr_67_5;

Selector_2 s67_5(wires_16_4[3], addr_16_4, wires_67_5,addr_67_5);

wire[3:0] wires_68_5;

wire[31:0] addr_68_5;

Selector_2 s68_5(wires_17_4[0], addr_17_4, wires_68_5,addr_68_5);

wire[3:0] wires_69_5;

wire[31:0] addr_69_5;

Selector_2 s69_5(wires_17_4[1], addr_17_4, wires_69_5,addr_69_5);

wire[3:0] wires_70_5;

wire[31:0] addr_70_5;

Selector_2 s70_5(wires_17_4[2], addr_17_4, wires_70_5,addr_70_5);

wire[3:0] wires_71_5;

wire[31:0] addr_71_5;

Selector_2 s71_5(wires_17_4[3], addr_17_4, wires_71_5,addr_71_5);

wire[3:0] wires_72_5;

wire[31:0] addr_72_5;

Selector_2 s72_5(wires_18_4[0], addr_18_4, wires_72_5,addr_72_5);

wire[3:0] wires_73_5;

wire[31:0] addr_73_5;

Selector_2 s73_5(wires_18_4[1], addr_18_4, wires_73_5,addr_73_5);

wire[3:0] wires_74_5;

wire[31:0] addr_74_5;

Selector_2 s74_5(wires_18_4[2], addr_18_4, wires_74_5,addr_74_5);

wire[3:0] wires_75_5;

wire[31:0] addr_75_5;

Selector_2 s75_5(wires_18_4[3], addr_18_4, wires_75_5,addr_75_5);

wire[3:0] wires_76_5;

wire[31:0] addr_76_5;

Selector_2 s76_5(wires_19_4[0], addr_19_4, wires_76_5,addr_76_5);

wire[3:0] wires_77_5;

wire[31:0] addr_77_5;

Selector_2 s77_5(wires_19_4[1], addr_19_4, wires_77_5,addr_77_5);

wire[3:0] wires_78_5;

wire[31:0] addr_78_5;

Selector_2 s78_5(wires_19_4[2], addr_19_4, wires_78_5,addr_78_5);

wire[3:0] wires_79_5;

wire[31:0] addr_79_5;

Selector_2 s79_5(wires_19_4[3], addr_19_4, wires_79_5,addr_79_5);

wire[3:0] wires_80_5;

wire[31:0] addr_80_5;

Selector_2 s80_5(wires_20_4[0], addr_20_4, wires_80_5,addr_80_5);

wire[3:0] wires_81_5;

wire[31:0] addr_81_5;

Selector_2 s81_5(wires_20_4[1], addr_20_4, wires_81_5,addr_81_5);

wire[3:0] wires_82_5;

wire[31:0] addr_82_5;

Selector_2 s82_5(wires_20_4[2], addr_20_4, wires_82_5,addr_82_5);

wire[3:0] wires_83_5;

wire[31:0] addr_83_5;

Selector_2 s83_5(wires_20_4[3], addr_20_4, wires_83_5,addr_83_5);

wire[3:0] wires_84_5;

wire[31:0] addr_84_5;

Selector_2 s84_5(wires_21_4[0], addr_21_4, wires_84_5,addr_84_5);

wire[3:0] wires_85_5;

wire[31:0] addr_85_5;

Selector_2 s85_5(wires_21_4[1], addr_21_4, wires_85_5,addr_85_5);

wire[3:0] wires_86_5;

wire[31:0] addr_86_5;

Selector_2 s86_5(wires_21_4[2], addr_21_4, wires_86_5,addr_86_5);

wire[3:0] wires_87_5;

wire[31:0] addr_87_5;

Selector_2 s87_5(wires_21_4[3], addr_21_4, wires_87_5,addr_87_5);

wire[3:0] wires_88_5;

wire[31:0] addr_88_5;

Selector_2 s88_5(wires_22_4[0], addr_22_4, wires_88_5,addr_88_5);

wire[3:0] wires_89_5;

wire[31:0] addr_89_5;

Selector_2 s89_5(wires_22_4[1], addr_22_4, wires_89_5,addr_89_5);

wire[3:0] wires_90_5;

wire[31:0] addr_90_5;

Selector_2 s90_5(wires_22_4[2], addr_22_4, wires_90_5,addr_90_5);

wire[3:0] wires_91_5;

wire[31:0] addr_91_5;

Selector_2 s91_5(wires_22_4[3], addr_22_4, wires_91_5,addr_91_5);

wire[3:0] wires_92_5;

wire[31:0] addr_92_5;

Selector_2 s92_5(wires_23_4[0], addr_23_4, wires_92_5,addr_92_5);

wire[3:0] wires_93_5;

wire[31:0] addr_93_5;

Selector_2 s93_5(wires_23_4[1], addr_23_4, wires_93_5,addr_93_5);

wire[3:0] wires_94_5;

wire[31:0] addr_94_5;

Selector_2 s94_5(wires_23_4[2], addr_23_4, wires_94_5,addr_94_5);

wire[3:0] wires_95_5;

wire[31:0] addr_95_5;

Selector_2 s95_5(wires_23_4[3], addr_23_4, wires_95_5,addr_95_5);

wire[3:0] wires_96_5;

wire[31:0] addr_96_5;

Selector_2 s96_5(wires_24_4[0], addr_24_4, wires_96_5,addr_96_5);

wire[3:0] wires_97_5;

wire[31:0] addr_97_5;

Selector_2 s97_5(wires_24_4[1], addr_24_4, wires_97_5,addr_97_5);

wire[3:0] wires_98_5;

wire[31:0] addr_98_5;

Selector_2 s98_5(wires_24_4[2], addr_24_4, wires_98_5,addr_98_5);

wire[3:0] wires_99_5;

wire[31:0] addr_99_5;

Selector_2 s99_5(wires_24_4[3], addr_24_4, wires_99_5,addr_99_5);

wire[3:0] wires_100_5;

wire[31:0] addr_100_5;

Selector_2 s100_5(wires_25_4[0], addr_25_4, wires_100_5,addr_100_5);

wire[3:0] wires_101_5;

wire[31:0] addr_101_5;

Selector_2 s101_5(wires_25_4[1], addr_25_4, wires_101_5,addr_101_5);

wire[3:0] wires_102_5;

wire[31:0] addr_102_5;

Selector_2 s102_5(wires_25_4[2], addr_25_4, wires_102_5,addr_102_5);

wire[3:0] wires_103_5;

wire[31:0] addr_103_5;

Selector_2 s103_5(wires_25_4[3], addr_25_4, wires_103_5,addr_103_5);

wire[3:0] wires_104_5;

wire[31:0] addr_104_5;

Selector_2 s104_5(wires_26_4[0], addr_26_4, wires_104_5,addr_104_5);

wire[3:0] wires_105_5;

wire[31:0] addr_105_5;

Selector_2 s105_5(wires_26_4[1], addr_26_4, wires_105_5,addr_105_5);

wire[3:0] wires_106_5;

wire[31:0] addr_106_5;

Selector_2 s106_5(wires_26_4[2], addr_26_4, wires_106_5,addr_106_5);

wire[3:0] wires_107_5;

wire[31:0] addr_107_5;

Selector_2 s107_5(wires_26_4[3], addr_26_4, wires_107_5,addr_107_5);

wire[3:0] wires_108_5;

wire[31:0] addr_108_5;

Selector_2 s108_5(wires_27_4[0], addr_27_4, wires_108_5,addr_108_5);

wire[3:0] wires_109_5;

wire[31:0] addr_109_5;

Selector_2 s109_5(wires_27_4[1], addr_27_4, wires_109_5,addr_109_5);

wire[3:0] wires_110_5;

wire[31:0] addr_110_5;

Selector_2 s110_5(wires_27_4[2], addr_27_4, wires_110_5,addr_110_5);

wire[3:0] wires_111_5;

wire[31:0] addr_111_5;

Selector_2 s111_5(wires_27_4[3], addr_27_4, wires_111_5,addr_111_5);

wire[3:0] wires_112_5;

wire[31:0] addr_112_5;

Selector_2 s112_5(wires_28_4[0], addr_28_4, wires_112_5,addr_112_5);

wire[3:0] wires_113_5;

wire[31:0] addr_113_5;

Selector_2 s113_5(wires_28_4[1], addr_28_4, wires_113_5,addr_113_5);

wire[3:0] wires_114_5;

wire[31:0] addr_114_5;

Selector_2 s114_5(wires_28_4[2], addr_28_4, wires_114_5,addr_114_5);

wire[3:0] wires_115_5;

wire[31:0] addr_115_5;

Selector_2 s115_5(wires_28_4[3], addr_28_4, wires_115_5,addr_115_5);

wire[3:0] wires_116_5;

wire[31:0] addr_116_5;

Selector_2 s116_5(wires_29_4[0], addr_29_4, wires_116_5,addr_116_5);

wire[3:0] wires_117_5;

wire[31:0] addr_117_5;

Selector_2 s117_5(wires_29_4[1], addr_29_4, wires_117_5,addr_117_5);

wire[3:0] wires_118_5;

wire[31:0] addr_118_5;

Selector_2 s118_5(wires_29_4[2], addr_29_4, wires_118_5,addr_118_5);

wire[3:0] wires_119_5;

wire[31:0] addr_119_5;

Selector_2 s119_5(wires_29_4[3], addr_29_4, wires_119_5,addr_119_5);

wire[3:0] wires_120_5;

wire[31:0] addr_120_5;

Selector_2 s120_5(wires_30_4[0], addr_30_4, wires_120_5,addr_120_5);

wire[3:0] wires_121_5;

wire[31:0] addr_121_5;

Selector_2 s121_5(wires_30_4[1], addr_30_4, wires_121_5,addr_121_5);

wire[3:0] wires_122_5;

wire[31:0] addr_122_5;

Selector_2 s122_5(wires_30_4[2], addr_30_4, wires_122_5,addr_122_5);

wire[3:0] wires_123_5;

wire[31:0] addr_123_5;

Selector_2 s123_5(wires_30_4[3], addr_30_4, wires_123_5,addr_123_5);

wire[3:0] wires_124_5;

wire[31:0] addr_124_5;

Selector_2 s124_5(wires_31_4[0], addr_31_4, wires_124_5,addr_124_5);

wire[3:0] wires_125_5;

wire[31:0] addr_125_5;

Selector_2 s125_5(wires_31_4[1], addr_31_4, wires_125_5,addr_125_5);

wire[3:0] wires_126_5;

wire[31:0] addr_126_5;

Selector_2 s126_5(wires_31_4[2], addr_31_4, wires_126_5,addr_126_5);

wire[3:0] wires_127_5;

wire[31:0] addr_127_5;

Selector_2 s127_5(wires_31_4[3], addr_31_4, wires_127_5,addr_127_5);

wire[3:0] wires_128_5;

wire[31:0] addr_128_5;

Selector_2 s128_5(wires_32_4[0], addr_32_4, wires_128_5,addr_128_5);

wire[3:0] wires_129_5;

wire[31:0] addr_129_5;

Selector_2 s129_5(wires_32_4[1], addr_32_4, wires_129_5,addr_129_5);

wire[3:0] wires_130_5;

wire[31:0] addr_130_5;

Selector_2 s130_5(wires_32_4[2], addr_32_4, wires_130_5,addr_130_5);

wire[3:0] wires_131_5;

wire[31:0] addr_131_5;

Selector_2 s131_5(wires_32_4[3], addr_32_4, wires_131_5,addr_131_5);

wire[3:0] wires_132_5;

wire[31:0] addr_132_5;

Selector_2 s132_5(wires_33_4[0], addr_33_4, wires_132_5,addr_132_5);

wire[3:0] wires_133_5;

wire[31:0] addr_133_5;

Selector_2 s133_5(wires_33_4[1], addr_33_4, wires_133_5,addr_133_5);

wire[3:0] wires_134_5;

wire[31:0] addr_134_5;

Selector_2 s134_5(wires_33_4[2], addr_33_4, wires_134_5,addr_134_5);

wire[3:0] wires_135_5;

wire[31:0] addr_135_5;

Selector_2 s135_5(wires_33_4[3], addr_33_4, wires_135_5,addr_135_5);

wire[3:0] wires_136_5;

wire[31:0] addr_136_5;

Selector_2 s136_5(wires_34_4[0], addr_34_4, wires_136_5,addr_136_5);

wire[3:0] wires_137_5;

wire[31:0] addr_137_5;

Selector_2 s137_5(wires_34_4[1], addr_34_4, wires_137_5,addr_137_5);

wire[3:0] wires_138_5;

wire[31:0] addr_138_5;

Selector_2 s138_5(wires_34_4[2], addr_34_4, wires_138_5,addr_138_5);

wire[3:0] wires_139_5;

wire[31:0] addr_139_5;

Selector_2 s139_5(wires_34_4[3], addr_34_4, wires_139_5,addr_139_5);

wire[3:0] wires_140_5;

wire[31:0] addr_140_5;

Selector_2 s140_5(wires_35_4[0], addr_35_4, wires_140_5,addr_140_5);

wire[3:0] wires_141_5;

wire[31:0] addr_141_5;

Selector_2 s141_5(wires_35_4[1], addr_35_4, wires_141_5,addr_141_5);

wire[3:0] wires_142_5;

wire[31:0] addr_142_5;

Selector_2 s142_5(wires_35_4[2], addr_35_4, wires_142_5,addr_142_5);

wire[3:0] wires_143_5;

wire[31:0] addr_143_5;

Selector_2 s143_5(wires_35_4[3], addr_35_4, wires_143_5,addr_143_5);

wire[3:0] wires_144_5;

wire[31:0] addr_144_5;

Selector_2 s144_5(wires_36_4[0], addr_36_4, wires_144_5,addr_144_5);

wire[3:0] wires_145_5;

wire[31:0] addr_145_5;

Selector_2 s145_5(wires_36_4[1], addr_36_4, wires_145_5,addr_145_5);

wire[3:0] wires_146_5;

wire[31:0] addr_146_5;

Selector_2 s146_5(wires_36_4[2], addr_36_4, wires_146_5,addr_146_5);

wire[3:0] wires_147_5;

wire[31:0] addr_147_5;

Selector_2 s147_5(wires_36_4[3], addr_36_4, wires_147_5,addr_147_5);

wire[3:0] wires_148_5;

wire[31:0] addr_148_5;

Selector_2 s148_5(wires_37_4[0], addr_37_4, wires_148_5,addr_148_5);

wire[3:0] wires_149_5;

wire[31:0] addr_149_5;

Selector_2 s149_5(wires_37_4[1], addr_37_4, wires_149_5,addr_149_5);

wire[3:0] wires_150_5;

wire[31:0] addr_150_5;

Selector_2 s150_5(wires_37_4[2], addr_37_4, wires_150_5,addr_150_5);

wire[3:0] wires_151_5;

wire[31:0] addr_151_5;

Selector_2 s151_5(wires_37_4[3], addr_37_4, wires_151_5,addr_151_5);

wire[3:0] wires_152_5;

wire[31:0] addr_152_5;

Selector_2 s152_5(wires_38_4[0], addr_38_4, wires_152_5,addr_152_5);

wire[3:0] wires_153_5;

wire[31:0] addr_153_5;

Selector_2 s153_5(wires_38_4[1], addr_38_4, wires_153_5,addr_153_5);

wire[3:0] wires_154_5;

wire[31:0] addr_154_5;

Selector_2 s154_5(wires_38_4[2], addr_38_4, wires_154_5,addr_154_5);

wire[3:0] wires_155_5;

wire[31:0] addr_155_5;

Selector_2 s155_5(wires_38_4[3], addr_38_4, wires_155_5,addr_155_5);

wire[3:0] wires_156_5;

wire[31:0] addr_156_5;

Selector_2 s156_5(wires_39_4[0], addr_39_4, wires_156_5,addr_156_5);

wire[3:0] wires_157_5;

wire[31:0] addr_157_5;

Selector_2 s157_5(wires_39_4[1], addr_39_4, wires_157_5,addr_157_5);

wire[3:0] wires_158_5;

wire[31:0] addr_158_5;

Selector_2 s158_5(wires_39_4[2], addr_39_4, wires_158_5,addr_158_5);

wire[3:0] wires_159_5;

wire[31:0] addr_159_5;

Selector_2 s159_5(wires_39_4[3], addr_39_4, wires_159_5,addr_159_5);

wire[3:0] wires_160_5;

wire[31:0] addr_160_5;

Selector_2 s160_5(wires_40_4[0], addr_40_4, wires_160_5,addr_160_5);

wire[3:0] wires_161_5;

wire[31:0] addr_161_5;

Selector_2 s161_5(wires_40_4[1], addr_40_4, wires_161_5,addr_161_5);

wire[3:0] wires_162_5;

wire[31:0] addr_162_5;

Selector_2 s162_5(wires_40_4[2], addr_40_4, wires_162_5,addr_162_5);

wire[3:0] wires_163_5;

wire[31:0] addr_163_5;

Selector_2 s163_5(wires_40_4[3], addr_40_4, wires_163_5,addr_163_5);

wire[3:0] wires_164_5;

wire[31:0] addr_164_5;

Selector_2 s164_5(wires_41_4[0], addr_41_4, wires_164_5,addr_164_5);

wire[3:0] wires_165_5;

wire[31:0] addr_165_5;

Selector_2 s165_5(wires_41_4[1], addr_41_4, wires_165_5,addr_165_5);

wire[3:0] wires_166_5;

wire[31:0] addr_166_5;

Selector_2 s166_5(wires_41_4[2], addr_41_4, wires_166_5,addr_166_5);

wire[3:0] wires_167_5;

wire[31:0] addr_167_5;

Selector_2 s167_5(wires_41_4[3], addr_41_4, wires_167_5,addr_167_5);

wire[3:0] wires_168_5;

wire[31:0] addr_168_5;

Selector_2 s168_5(wires_42_4[0], addr_42_4, wires_168_5,addr_168_5);

wire[3:0] wires_169_5;

wire[31:0] addr_169_5;

Selector_2 s169_5(wires_42_4[1], addr_42_4, wires_169_5,addr_169_5);

wire[3:0] wires_170_5;

wire[31:0] addr_170_5;

Selector_2 s170_5(wires_42_4[2], addr_42_4, wires_170_5,addr_170_5);

wire[3:0] wires_171_5;

wire[31:0] addr_171_5;

Selector_2 s171_5(wires_42_4[3], addr_42_4, wires_171_5,addr_171_5);

wire[3:0] wires_172_5;

wire[31:0] addr_172_5;

Selector_2 s172_5(wires_43_4[0], addr_43_4, wires_172_5,addr_172_5);

wire[3:0] wires_173_5;

wire[31:0] addr_173_5;

Selector_2 s173_5(wires_43_4[1], addr_43_4, wires_173_5,addr_173_5);

wire[3:0] wires_174_5;

wire[31:0] addr_174_5;

Selector_2 s174_5(wires_43_4[2], addr_43_4, wires_174_5,addr_174_5);

wire[3:0] wires_175_5;

wire[31:0] addr_175_5;

Selector_2 s175_5(wires_43_4[3], addr_43_4, wires_175_5,addr_175_5);

wire[3:0] wires_176_5;

wire[31:0] addr_176_5;

Selector_2 s176_5(wires_44_4[0], addr_44_4, wires_176_5,addr_176_5);

wire[3:0] wires_177_5;

wire[31:0] addr_177_5;

Selector_2 s177_5(wires_44_4[1], addr_44_4, wires_177_5,addr_177_5);

wire[3:0] wires_178_5;

wire[31:0] addr_178_5;

Selector_2 s178_5(wires_44_4[2], addr_44_4, wires_178_5,addr_178_5);

wire[3:0] wires_179_5;

wire[31:0] addr_179_5;

Selector_2 s179_5(wires_44_4[3], addr_44_4, wires_179_5,addr_179_5);

wire[3:0] wires_180_5;

wire[31:0] addr_180_5;

Selector_2 s180_5(wires_45_4[0], addr_45_4, wires_180_5,addr_180_5);

wire[3:0] wires_181_5;

wire[31:0] addr_181_5;

Selector_2 s181_5(wires_45_4[1], addr_45_4, wires_181_5,addr_181_5);

wire[3:0] wires_182_5;

wire[31:0] addr_182_5;

Selector_2 s182_5(wires_45_4[2], addr_45_4, wires_182_5,addr_182_5);

wire[3:0] wires_183_5;

wire[31:0] addr_183_5;

Selector_2 s183_5(wires_45_4[3], addr_45_4, wires_183_5,addr_183_5);

wire[3:0] wires_184_5;

wire[31:0] addr_184_5;

Selector_2 s184_5(wires_46_4[0], addr_46_4, wires_184_5,addr_184_5);

wire[3:0] wires_185_5;

wire[31:0] addr_185_5;

Selector_2 s185_5(wires_46_4[1], addr_46_4, wires_185_5,addr_185_5);

wire[3:0] wires_186_5;

wire[31:0] addr_186_5;

Selector_2 s186_5(wires_46_4[2], addr_46_4, wires_186_5,addr_186_5);

wire[3:0] wires_187_5;

wire[31:0] addr_187_5;

Selector_2 s187_5(wires_46_4[3], addr_46_4, wires_187_5,addr_187_5);

wire[3:0] wires_188_5;

wire[31:0] addr_188_5;

Selector_2 s188_5(wires_47_4[0], addr_47_4, wires_188_5,addr_188_5);

wire[3:0] wires_189_5;

wire[31:0] addr_189_5;

Selector_2 s189_5(wires_47_4[1], addr_47_4, wires_189_5,addr_189_5);

wire[3:0] wires_190_5;

wire[31:0] addr_190_5;

Selector_2 s190_5(wires_47_4[2], addr_47_4, wires_190_5,addr_190_5);

wire[3:0] wires_191_5;

wire[31:0] addr_191_5;

Selector_2 s191_5(wires_47_4[3], addr_47_4, wires_191_5,addr_191_5);

wire[3:0] wires_192_5;

wire[31:0] addr_192_5;

Selector_2 s192_5(wires_48_4[0], addr_48_4, wires_192_5,addr_192_5);

wire[3:0] wires_193_5;

wire[31:0] addr_193_5;

Selector_2 s193_5(wires_48_4[1], addr_48_4, wires_193_5,addr_193_5);

wire[3:0] wires_194_5;

wire[31:0] addr_194_5;

Selector_2 s194_5(wires_48_4[2], addr_48_4, wires_194_5,addr_194_5);

wire[3:0] wires_195_5;

wire[31:0] addr_195_5;

Selector_2 s195_5(wires_48_4[3], addr_48_4, wires_195_5,addr_195_5);

wire[3:0] wires_196_5;

wire[31:0] addr_196_5;

Selector_2 s196_5(wires_49_4[0], addr_49_4, wires_196_5,addr_196_5);

wire[3:0] wires_197_5;

wire[31:0] addr_197_5;

Selector_2 s197_5(wires_49_4[1], addr_49_4, wires_197_5,addr_197_5);

wire[3:0] wires_198_5;

wire[31:0] addr_198_5;

Selector_2 s198_5(wires_49_4[2], addr_49_4, wires_198_5,addr_198_5);

wire[3:0] wires_199_5;

wire[31:0] addr_199_5;

Selector_2 s199_5(wires_49_4[3], addr_49_4, wires_199_5,addr_199_5);

wire[3:0] wires_200_5;

wire[31:0] addr_200_5;

Selector_2 s200_5(wires_50_4[0], addr_50_4, wires_200_5,addr_200_5);

wire[3:0] wires_201_5;

wire[31:0] addr_201_5;

Selector_2 s201_5(wires_50_4[1], addr_50_4, wires_201_5,addr_201_5);

wire[3:0] wires_202_5;

wire[31:0] addr_202_5;

Selector_2 s202_5(wires_50_4[2], addr_50_4, wires_202_5,addr_202_5);

wire[3:0] wires_203_5;

wire[31:0] addr_203_5;

Selector_2 s203_5(wires_50_4[3], addr_50_4, wires_203_5,addr_203_5);

wire[3:0] wires_204_5;

wire[31:0] addr_204_5;

Selector_2 s204_5(wires_51_4[0], addr_51_4, wires_204_5,addr_204_5);

wire[3:0] wires_205_5;

wire[31:0] addr_205_5;

Selector_2 s205_5(wires_51_4[1], addr_51_4, wires_205_5,addr_205_5);

wire[3:0] wires_206_5;

wire[31:0] addr_206_5;

Selector_2 s206_5(wires_51_4[2], addr_51_4, wires_206_5,addr_206_5);

wire[3:0] wires_207_5;

wire[31:0] addr_207_5;

Selector_2 s207_5(wires_51_4[3], addr_51_4, wires_207_5,addr_207_5);

wire[3:0] wires_208_5;

wire[31:0] addr_208_5;

Selector_2 s208_5(wires_52_4[0], addr_52_4, wires_208_5,addr_208_5);

wire[3:0] wires_209_5;

wire[31:0] addr_209_5;

Selector_2 s209_5(wires_52_4[1], addr_52_4, wires_209_5,addr_209_5);

wire[3:0] wires_210_5;

wire[31:0] addr_210_5;

Selector_2 s210_5(wires_52_4[2], addr_52_4, wires_210_5,addr_210_5);

wire[3:0] wires_211_5;

wire[31:0] addr_211_5;

Selector_2 s211_5(wires_52_4[3], addr_52_4, wires_211_5,addr_211_5);

wire[3:0] wires_212_5;

wire[31:0] addr_212_5;

Selector_2 s212_5(wires_53_4[0], addr_53_4, wires_212_5,addr_212_5);

wire[3:0] wires_213_5;

wire[31:0] addr_213_5;

Selector_2 s213_5(wires_53_4[1], addr_53_4, wires_213_5,addr_213_5);

wire[3:0] wires_214_5;

wire[31:0] addr_214_5;

Selector_2 s214_5(wires_53_4[2], addr_53_4, wires_214_5,addr_214_5);

wire[3:0] wires_215_5;

wire[31:0] addr_215_5;

Selector_2 s215_5(wires_53_4[3], addr_53_4, wires_215_5,addr_215_5);

wire[3:0] wires_216_5;

wire[31:0] addr_216_5;

Selector_2 s216_5(wires_54_4[0], addr_54_4, wires_216_5,addr_216_5);

wire[3:0] wires_217_5;

wire[31:0] addr_217_5;

Selector_2 s217_5(wires_54_4[1], addr_54_4, wires_217_5,addr_217_5);

wire[3:0] wires_218_5;

wire[31:0] addr_218_5;

Selector_2 s218_5(wires_54_4[2], addr_54_4, wires_218_5,addr_218_5);

wire[3:0] wires_219_5;

wire[31:0] addr_219_5;

Selector_2 s219_5(wires_54_4[3], addr_54_4, wires_219_5,addr_219_5);

wire[3:0] wires_220_5;

wire[31:0] addr_220_5;

Selector_2 s220_5(wires_55_4[0], addr_55_4, wires_220_5,addr_220_5);

wire[3:0] wires_221_5;

wire[31:0] addr_221_5;

Selector_2 s221_5(wires_55_4[1], addr_55_4, wires_221_5,addr_221_5);

wire[3:0] wires_222_5;

wire[31:0] addr_222_5;

Selector_2 s222_5(wires_55_4[2], addr_55_4, wires_222_5,addr_222_5);

wire[3:0] wires_223_5;

wire[31:0] addr_223_5;

Selector_2 s223_5(wires_55_4[3], addr_55_4, wires_223_5,addr_223_5);

wire[3:0] wires_224_5;

wire[31:0] addr_224_5;

Selector_2 s224_5(wires_56_4[0], addr_56_4, wires_224_5,addr_224_5);

wire[3:0] wires_225_5;

wire[31:0] addr_225_5;

Selector_2 s225_5(wires_56_4[1], addr_56_4, wires_225_5,addr_225_5);

wire[3:0] wires_226_5;

wire[31:0] addr_226_5;

Selector_2 s226_5(wires_56_4[2], addr_56_4, wires_226_5,addr_226_5);

wire[3:0] wires_227_5;

wire[31:0] addr_227_5;

Selector_2 s227_5(wires_56_4[3], addr_56_4, wires_227_5,addr_227_5);

wire[3:0] wires_228_5;

wire[31:0] addr_228_5;

Selector_2 s228_5(wires_57_4[0], addr_57_4, wires_228_5,addr_228_5);

wire[3:0] wires_229_5;

wire[31:0] addr_229_5;

Selector_2 s229_5(wires_57_4[1], addr_57_4, wires_229_5,addr_229_5);

wire[3:0] wires_230_5;

wire[31:0] addr_230_5;

Selector_2 s230_5(wires_57_4[2], addr_57_4, wires_230_5,addr_230_5);

wire[3:0] wires_231_5;

wire[31:0] addr_231_5;

Selector_2 s231_5(wires_57_4[3], addr_57_4, wires_231_5,addr_231_5);

wire[3:0] wires_232_5;

wire[31:0] addr_232_5;

Selector_2 s232_5(wires_58_4[0], addr_58_4, wires_232_5,addr_232_5);

wire[3:0] wires_233_5;

wire[31:0] addr_233_5;

Selector_2 s233_5(wires_58_4[1], addr_58_4, wires_233_5,addr_233_5);

wire[3:0] wires_234_5;

wire[31:0] addr_234_5;

Selector_2 s234_5(wires_58_4[2], addr_58_4, wires_234_5,addr_234_5);

wire[3:0] wires_235_5;

wire[31:0] addr_235_5;

Selector_2 s235_5(wires_58_4[3], addr_58_4, wires_235_5,addr_235_5);

wire[3:0] wires_236_5;

wire[31:0] addr_236_5;

Selector_2 s236_5(wires_59_4[0], addr_59_4, wires_236_5,addr_236_5);

wire[3:0] wires_237_5;

wire[31:0] addr_237_5;

Selector_2 s237_5(wires_59_4[1], addr_59_4, wires_237_5,addr_237_5);

wire[3:0] wires_238_5;

wire[31:0] addr_238_5;

Selector_2 s238_5(wires_59_4[2], addr_59_4, wires_238_5,addr_238_5);

wire[3:0] wires_239_5;

wire[31:0] addr_239_5;

Selector_2 s239_5(wires_59_4[3], addr_59_4, wires_239_5,addr_239_5);

wire[3:0] wires_240_5;

wire[31:0] addr_240_5;

Selector_2 s240_5(wires_60_4[0], addr_60_4, wires_240_5,addr_240_5);

wire[3:0] wires_241_5;

wire[31:0] addr_241_5;

Selector_2 s241_5(wires_60_4[1], addr_60_4, wires_241_5,addr_241_5);

wire[3:0] wires_242_5;

wire[31:0] addr_242_5;

Selector_2 s242_5(wires_60_4[2], addr_60_4, wires_242_5,addr_242_5);

wire[3:0] wires_243_5;

wire[31:0] addr_243_5;

Selector_2 s243_5(wires_60_4[3], addr_60_4, wires_243_5,addr_243_5);

wire[3:0] wires_244_5;

wire[31:0] addr_244_5;

Selector_2 s244_5(wires_61_4[0], addr_61_4, wires_244_5,addr_244_5);

wire[3:0] wires_245_5;

wire[31:0] addr_245_5;

Selector_2 s245_5(wires_61_4[1], addr_61_4, wires_245_5,addr_245_5);

wire[3:0] wires_246_5;

wire[31:0] addr_246_5;

Selector_2 s246_5(wires_61_4[2], addr_61_4, wires_246_5,addr_246_5);

wire[3:0] wires_247_5;

wire[31:0] addr_247_5;

Selector_2 s247_5(wires_61_4[3], addr_61_4, wires_247_5,addr_247_5);

wire[3:0] wires_248_5;

wire[31:0] addr_248_5;

Selector_2 s248_5(wires_62_4[0], addr_62_4, wires_248_5,addr_248_5);

wire[3:0] wires_249_5;

wire[31:0] addr_249_5;

Selector_2 s249_5(wires_62_4[1], addr_62_4, wires_249_5,addr_249_5);

wire[3:0] wires_250_5;

wire[31:0] addr_250_5;

Selector_2 s250_5(wires_62_4[2], addr_62_4, wires_250_5,addr_250_5);

wire[3:0] wires_251_5;

wire[31:0] addr_251_5;

Selector_2 s251_5(wires_62_4[3], addr_62_4, wires_251_5,addr_251_5);

wire[3:0] wires_252_5;

wire[31:0] addr_252_5;

Selector_2 s252_5(wires_63_4[0], addr_63_4, wires_252_5,addr_252_5);

wire[3:0] wires_253_5;

wire[31:0] addr_253_5;

Selector_2 s253_5(wires_63_4[1], addr_63_4, wires_253_5,addr_253_5);

wire[3:0] wires_254_5;

wire[31:0] addr_254_5;

Selector_2 s254_5(wires_63_4[2], addr_63_4, wires_254_5,addr_254_5);

wire[3:0] wires_255_5;

wire[31:0] addr_255_5;

Selector_2 s255_5(wires_63_4[3], addr_63_4, wires_255_5,addr_255_5);

wire[3:0] wires_256_5;

wire[31:0] addr_256_5;

Selector_2 s256_5(wires_64_4[0], addr_64_4, wires_256_5,addr_256_5);

wire[3:0] wires_257_5;

wire[31:0] addr_257_5;

Selector_2 s257_5(wires_64_4[1], addr_64_4, wires_257_5,addr_257_5);

wire[3:0] wires_258_5;

wire[31:0] addr_258_5;

Selector_2 s258_5(wires_64_4[2], addr_64_4, wires_258_5,addr_258_5);

wire[3:0] wires_259_5;

wire[31:0] addr_259_5;

Selector_2 s259_5(wires_64_4[3], addr_64_4, wires_259_5,addr_259_5);

wire[3:0] wires_260_5;

wire[31:0] addr_260_5;

Selector_2 s260_5(wires_65_4[0], addr_65_4, wires_260_5,addr_260_5);

wire[3:0] wires_261_5;

wire[31:0] addr_261_5;

Selector_2 s261_5(wires_65_4[1], addr_65_4, wires_261_5,addr_261_5);

wire[3:0] wires_262_5;

wire[31:0] addr_262_5;

Selector_2 s262_5(wires_65_4[2], addr_65_4, wires_262_5,addr_262_5);

wire[3:0] wires_263_5;

wire[31:0] addr_263_5;

Selector_2 s263_5(wires_65_4[3], addr_65_4, wires_263_5,addr_263_5);

wire[3:0] wires_264_5;

wire[31:0] addr_264_5;

Selector_2 s264_5(wires_66_4[0], addr_66_4, wires_264_5,addr_264_5);

wire[3:0] wires_265_5;

wire[31:0] addr_265_5;

Selector_2 s265_5(wires_66_4[1], addr_66_4, wires_265_5,addr_265_5);

wire[3:0] wires_266_5;

wire[31:0] addr_266_5;

Selector_2 s266_5(wires_66_4[2], addr_66_4, wires_266_5,addr_266_5);

wire[3:0] wires_267_5;

wire[31:0] addr_267_5;

Selector_2 s267_5(wires_66_4[3], addr_66_4, wires_267_5,addr_267_5);

wire[3:0] wires_268_5;

wire[31:0] addr_268_5;

Selector_2 s268_5(wires_67_4[0], addr_67_4, wires_268_5,addr_268_5);

wire[3:0] wires_269_5;

wire[31:0] addr_269_5;

Selector_2 s269_5(wires_67_4[1], addr_67_4, wires_269_5,addr_269_5);

wire[3:0] wires_270_5;

wire[31:0] addr_270_5;

Selector_2 s270_5(wires_67_4[2], addr_67_4, wires_270_5,addr_270_5);

wire[3:0] wires_271_5;

wire[31:0] addr_271_5;

Selector_2 s271_5(wires_67_4[3], addr_67_4, wires_271_5,addr_271_5);

wire[3:0] wires_272_5;

wire[31:0] addr_272_5;

Selector_2 s272_5(wires_68_4[0], addr_68_4, wires_272_5,addr_272_5);

wire[3:0] wires_273_5;

wire[31:0] addr_273_5;

Selector_2 s273_5(wires_68_4[1], addr_68_4, wires_273_5,addr_273_5);

wire[3:0] wires_274_5;

wire[31:0] addr_274_5;

Selector_2 s274_5(wires_68_4[2], addr_68_4, wires_274_5,addr_274_5);

wire[3:0] wires_275_5;

wire[31:0] addr_275_5;

Selector_2 s275_5(wires_68_4[3], addr_68_4, wires_275_5,addr_275_5);

wire[3:0] wires_276_5;

wire[31:0] addr_276_5;

Selector_2 s276_5(wires_69_4[0], addr_69_4, wires_276_5,addr_276_5);

wire[3:0] wires_277_5;

wire[31:0] addr_277_5;

Selector_2 s277_5(wires_69_4[1], addr_69_4, wires_277_5,addr_277_5);

wire[3:0] wires_278_5;

wire[31:0] addr_278_5;

Selector_2 s278_5(wires_69_4[2], addr_69_4, wires_278_5,addr_278_5);

wire[3:0] wires_279_5;

wire[31:0] addr_279_5;

Selector_2 s279_5(wires_69_4[3], addr_69_4, wires_279_5,addr_279_5);

wire[3:0] wires_280_5;

wire[31:0] addr_280_5;

Selector_2 s280_5(wires_70_4[0], addr_70_4, wires_280_5,addr_280_5);

wire[3:0] wires_281_5;

wire[31:0] addr_281_5;

Selector_2 s281_5(wires_70_4[1], addr_70_4, wires_281_5,addr_281_5);

wire[3:0] wires_282_5;

wire[31:0] addr_282_5;

Selector_2 s282_5(wires_70_4[2], addr_70_4, wires_282_5,addr_282_5);

wire[3:0] wires_283_5;

wire[31:0] addr_283_5;

Selector_2 s283_5(wires_70_4[3], addr_70_4, wires_283_5,addr_283_5);

wire[3:0] wires_284_5;

wire[31:0] addr_284_5;

Selector_2 s284_5(wires_71_4[0], addr_71_4, wires_284_5,addr_284_5);

wire[3:0] wires_285_5;

wire[31:0] addr_285_5;

Selector_2 s285_5(wires_71_4[1], addr_71_4, wires_285_5,addr_285_5);

wire[3:0] wires_286_5;

wire[31:0] addr_286_5;

Selector_2 s286_5(wires_71_4[2], addr_71_4, wires_286_5,addr_286_5);

wire[3:0] wires_287_5;

wire[31:0] addr_287_5;

Selector_2 s287_5(wires_71_4[3], addr_71_4, wires_287_5,addr_287_5);

wire[3:0] wires_288_5;

wire[31:0] addr_288_5;

Selector_2 s288_5(wires_72_4[0], addr_72_4, wires_288_5,addr_288_5);

wire[3:0] wires_289_5;

wire[31:0] addr_289_5;

Selector_2 s289_5(wires_72_4[1], addr_72_4, wires_289_5,addr_289_5);

wire[3:0] wires_290_5;

wire[31:0] addr_290_5;

Selector_2 s290_5(wires_72_4[2], addr_72_4, wires_290_5,addr_290_5);

wire[3:0] wires_291_5;

wire[31:0] addr_291_5;

Selector_2 s291_5(wires_72_4[3], addr_72_4, wires_291_5,addr_291_5);

wire[3:0] wires_292_5;

wire[31:0] addr_292_5;

Selector_2 s292_5(wires_73_4[0], addr_73_4, wires_292_5,addr_292_5);

wire[3:0] wires_293_5;

wire[31:0] addr_293_5;

Selector_2 s293_5(wires_73_4[1], addr_73_4, wires_293_5,addr_293_5);

wire[3:0] wires_294_5;

wire[31:0] addr_294_5;

Selector_2 s294_5(wires_73_4[2], addr_73_4, wires_294_5,addr_294_5);

wire[3:0] wires_295_5;

wire[31:0] addr_295_5;

Selector_2 s295_5(wires_73_4[3], addr_73_4, wires_295_5,addr_295_5);

wire[3:0] wires_296_5;

wire[31:0] addr_296_5;

Selector_2 s296_5(wires_74_4[0], addr_74_4, wires_296_5,addr_296_5);

wire[3:0] wires_297_5;

wire[31:0] addr_297_5;

Selector_2 s297_5(wires_74_4[1], addr_74_4, wires_297_5,addr_297_5);

wire[3:0] wires_298_5;

wire[31:0] addr_298_5;

Selector_2 s298_5(wires_74_4[2], addr_74_4, wires_298_5,addr_298_5);

wire[3:0] wires_299_5;

wire[31:0] addr_299_5;

Selector_2 s299_5(wires_74_4[3], addr_74_4, wires_299_5,addr_299_5);

wire[3:0] wires_300_5;

wire[31:0] addr_300_5;

Selector_2 s300_5(wires_75_4[0], addr_75_4, wires_300_5,addr_300_5);

wire[3:0] wires_301_5;

wire[31:0] addr_301_5;

Selector_2 s301_5(wires_75_4[1], addr_75_4, wires_301_5,addr_301_5);

wire[3:0] wires_302_5;

wire[31:0] addr_302_5;

Selector_2 s302_5(wires_75_4[2], addr_75_4, wires_302_5,addr_302_5);

wire[3:0] wires_303_5;

wire[31:0] addr_303_5;

Selector_2 s303_5(wires_75_4[3], addr_75_4, wires_303_5,addr_303_5);

wire[3:0] wires_304_5;

wire[31:0] addr_304_5;

Selector_2 s304_5(wires_76_4[0], addr_76_4, wires_304_5,addr_304_5);

wire[3:0] wires_305_5;

wire[31:0] addr_305_5;

Selector_2 s305_5(wires_76_4[1], addr_76_4, wires_305_5,addr_305_5);

wire[3:0] wires_306_5;

wire[31:0] addr_306_5;

Selector_2 s306_5(wires_76_4[2], addr_76_4, wires_306_5,addr_306_5);

wire[3:0] wires_307_5;

wire[31:0] addr_307_5;

Selector_2 s307_5(wires_76_4[3], addr_76_4, wires_307_5,addr_307_5);

wire[3:0] wires_308_5;

wire[31:0] addr_308_5;

Selector_2 s308_5(wires_77_4[0], addr_77_4, wires_308_5,addr_308_5);

wire[3:0] wires_309_5;

wire[31:0] addr_309_5;

Selector_2 s309_5(wires_77_4[1], addr_77_4, wires_309_5,addr_309_5);

wire[3:0] wires_310_5;

wire[31:0] addr_310_5;

Selector_2 s310_5(wires_77_4[2], addr_77_4, wires_310_5,addr_310_5);

wire[3:0] wires_311_5;

wire[31:0] addr_311_5;

Selector_2 s311_5(wires_77_4[3], addr_77_4, wires_311_5,addr_311_5);

wire[3:0] wires_312_5;

wire[31:0] addr_312_5;

Selector_2 s312_5(wires_78_4[0], addr_78_4, wires_312_5,addr_312_5);

wire[3:0] wires_313_5;

wire[31:0] addr_313_5;

Selector_2 s313_5(wires_78_4[1], addr_78_4, wires_313_5,addr_313_5);

wire[3:0] wires_314_5;

wire[31:0] addr_314_5;

Selector_2 s314_5(wires_78_4[2], addr_78_4, wires_314_5,addr_314_5);

wire[3:0] wires_315_5;

wire[31:0] addr_315_5;

Selector_2 s315_5(wires_78_4[3], addr_78_4, wires_315_5,addr_315_5);

wire[3:0] wires_316_5;

wire[31:0] addr_316_5;

Selector_2 s316_5(wires_79_4[0], addr_79_4, wires_316_5,addr_316_5);

wire[3:0] wires_317_5;

wire[31:0] addr_317_5;

Selector_2 s317_5(wires_79_4[1], addr_79_4, wires_317_5,addr_317_5);

wire[3:0] wires_318_5;

wire[31:0] addr_318_5;

Selector_2 s318_5(wires_79_4[2], addr_79_4, wires_318_5,addr_318_5);

wire[3:0] wires_319_5;

wire[31:0] addr_319_5;

Selector_2 s319_5(wires_79_4[3], addr_79_4, wires_319_5,addr_319_5);

wire[3:0] wires_320_5;

wire[31:0] addr_320_5;

Selector_2 s320_5(wires_80_4[0], addr_80_4, wires_320_5,addr_320_5);

wire[3:0] wires_321_5;

wire[31:0] addr_321_5;

Selector_2 s321_5(wires_80_4[1], addr_80_4, wires_321_5,addr_321_5);

wire[3:0] wires_322_5;

wire[31:0] addr_322_5;

Selector_2 s322_5(wires_80_4[2], addr_80_4, wires_322_5,addr_322_5);

wire[3:0] wires_323_5;

wire[31:0] addr_323_5;

Selector_2 s323_5(wires_80_4[3], addr_80_4, wires_323_5,addr_323_5);

wire[3:0] wires_324_5;

wire[31:0] addr_324_5;

Selector_2 s324_5(wires_81_4[0], addr_81_4, wires_324_5,addr_324_5);

wire[3:0] wires_325_5;

wire[31:0] addr_325_5;

Selector_2 s325_5(wires_81_4[1], addr_81_4, wires_325_5,addr_325_5);

wire[3:0] wires_326_5;

wire[31:0] addr_326_5;

Selector_2 s326_5(wires_81_4[2], addr_81_4, wires_326_5,addr_326_5);

wire[3:0] wires_327_5;

wire[31:0] addr_327_5;

Selector_2 s327_5(wires_81_4[3], addr_81_4, wires_327_5,addr_327_5);

wire[3:0] wires_328_5;

wire[31:0] addr_328_5;

Selector_2 s328_5(wires_82_4[0], addr_82_4, wires_328_5,addr_328_5);

wire[3:0] wires_329_5;

wire[31:0] addr_329_5;

Selector_2 s329_5(wires_82_4[1], addr_82_4, wires_329_5,addr_329_5);

wire[3:0] wires_330_5;

wire[31:0] addr_330_5;

Selector_2 s330_5(wires_82_4[2], addr_82_4, wires_330_5,addr_330_5);

wire[3:0] wires_331_5;

wire[31:0] addr_331_5;

Selector_2 s331_5(wires_82_4[3], addr_82_4, wires_331_5,addr_331_5);

wire[3:0] wires_332_5;

wire[31:0] addr_332_5;

Selector_2 s332_5(wires_83_4[0], addr_83_4, wires_332_5,addr_332_5);

wire[3:0] wires_333_5;

wire[31:0] addr_333_5;

Selector_2 s333_5(wires_83_4[1], addr_83_4, wires_333_5,addr_333_5);

wire[3:0] wires_334_5;

wire[31:0] addr_334_5;

Selector_2 s334_5(wires_83_4[2], addr_83_4, wires_334_5,addr_334_5);

wire[3:0] wires_335_5;

wire[31:0] addr_335_5;

Selector_2 s335_5(wires_83_4[3], addr_83_4, wires_335_5,addr_335_5);

wire[3:0] wires_336_5;

wire[31:0] addr_336_5;

Selector_2 s336_5(wires_84_4[0], addr_84_4, wires_336_5,addr_336_5);

wire[3:0] wires_337_5;

wire[31:0] addr_337_5;

Selector_2 s337_5(wires_84_4[1], addr_84_4, wires_337_5,addr_337_5);

wire[3:0] wires_338_5;

wire[31:0] addr_338_5;

Selector_2 s338_5(wires_84_4[2], addr_84_4, wires_338_5,addr_338_5);

wire[3:0] wires_339_5;

wire[31:0] addr_339_5;

Selector_2 s339_5(wires_84_4[3], addr_84_4, wires_339_5,addr_339_5);

wire[3:0] wires_340_5;

wire[31:0] addr_340_5;

Selector_2 s340_5(wires_85_4[0], addr_85_4, wires_340_5,addr_340_5);

wire[3:0] wires_341_5;

wire[31:0] addr_341_5;

Selector_2 s341_5(wires_85_4[1], addr_85_4, wires_341_5,addr_341_5);

wire[3:0] wires_342_5;

wire[31:0] addr_342_5;

Selector_2 s342_5(wires_85_4[2], addr_85_4, wires_342_5,addr_342_5);

wire[3:0] wires_343_5;

wire[31:0] addr_343_5;

Selector_2 s343_5(wires_85_4[3], addr_85_4, wires_343_5,addr_343_5);

wire[3:0] wires_344_5;

wire[31:0] addr_344_5;

Selector_2 s344_5(wires_86_4[0], addr_86_4, wires_344_5,addr_344_5);

wire[3:0] wires_345_5;

wire[31:0] addr_345_5;

Selector_2 s345_5(wires_86_4[1], addr_86_4, wires_345_5,addr_345_5);

wire[3:0] wires_346_5;

wire[31:0] addr_346_5;

Selector_2 s346_5(wires_86_4[2], addr_86_4, wires_346_5,addr_346_5);

wire[3:0] wires_347_5;

wire[31:0] addr_347_5;

Selector_2 s347_5(wires_86_4[3], addr_86_4, wires_347_5,addr_347_5);

wire[3:0] wires_348_5;

wire[31:0] addr_348_5;

Selector_2 s348_5(wires_87_4[0], addr_87_4, wires_348_5,addr_348_5);

wire[3:0] wires_349_5;

wire[31:0] addr_349_5;

Selector_2 s349_5(wires_87_4[1], addr_87_4, wires_349_5,addr_349_5);

wire[3:0] wires_350_5;

wire[31:0] addr_350_5;

Selector_2 s350_5(wires_87_4[2], addr_87_4, wires_350_5,addr_350_5);

wire[3:0] wires_351_5;

wire[31:0] addr_351_5;

Selector_2 s351_5(wires_87_4[3], addr_87_4, wires_351_5,addr_351_5);

wire[3:0] wires_352_5;

wire[31:0] addr_352_5;

Selector_2 s352_5(wires_88_4[0], addr_88_4, wires_352_5,addr_352_5);

wire[3:0] wires_353_5;

wire[31:0] addr_353_5;

Selector_2 s353_5(wires_88_4[1], addr_88_4, wires_353_5,addr_353_5);

wire[3:0] wires_354_5;

wire[31:0] addr_354_5;

Selector_2 s354_5(wires_88_4[2], addr_88_4, wires_354_5,addr_354_5);

wire[3:0] wires_355_5;

wire[31:0] addr_355_5;

Selector_2 s355_5(wires_88_4[3], addr_88_4, wires_355_5,addr_355_5);

wire[3:0] wires_356_5;

wire[31:0] addr_356_5;

Selector_2 s356_5(wires_89_4[0], addr_89_4, wires_356_5,addr_356_5);

wire[3:0] wires_357_5;

wire[31:0] addr_357_5;

Selector_2 s357_5(wires_89_4[1], addr_89_4, wires_357_5,addr_357_5);

wire[3:0] wires_358_5;

wire[31:0] addr_358_5;

Selector_2 s358_5(wires_89_4[2], addr_89_4, wires_358_5,addr_358_5);

wire[3:0] wires_359_5;

wire[31:0] addr_359_5;

Selector_2 s359_5(wires_89_4[3], addr_89_4, wires_359_5,addr_359_5);

wire[3:0] wires_360_5;

wire[31:0] addr_360_5;

Selector_2 s360_5(wires_90_4[0], addr_90_4, wires_360_5,addr_360_5);

wire[3:0] wires_361_5;

wire[31:0] addr_361_5;

Selector_2 s361_5(wires_90_4[1], addr_90_4, wires_361_5,addr_361_5);

wire[3:0] wires_362_5;

wire[31:0] addr_362_5;

Selector_2 s362_5(wires_90_4[2], addr_90_4, wires_362_5,addr_362_5);

wire[3:0] wires_363_5;

wire[31:0] addr_363_5;

Selector_2 s363_5(wires_90_4[3], addr_90_4, wires_363_5,addr_363_5);

wire[3:0] wires_364_5;

wire[31:0] addr_364_5;

Selector_2 s364_5(wires_91_4[0], addr_91_4, wires_364_5,addr_364_5);

wire[3:0] wires_365_5;

wire[31:0] addr_365_5;

Selector_2 s365_5(wires_91_4[1], addr_91_4, wires_365_5,addr_365_5);

wire[3:0] wires_366_5;

wire[31:0] addr_366_5;

Selector_2 s366_5(wires_91_4[2], addr_91_4, wires_366_5,addr_366_5);

wire[3:0] wires_367_5;

wire[31:0] addr_367_5;

Selector_2 s367_5(wires_91_4[3], addr_91_4, wires_367_5,addr_367_5);

wire[3:0] wires_368_5;

wire[31:0] addr_368_5;

Selector_2 s368_5(wires_92_4[0], addr_92_4, wires_368_5,addr_368_5);

wire[3:0] wires_369_5;

wire[31:0] addr_369_5;

Selector_2 s369_5(wires_92_4[1], addr_92_4, wires_369_5,addr_369_5);

wire[3:0] wires_370_5;

wire[31:0] addr_370_5;

Selector_2 s370_5(wires_92_4[2], addr_92_4, wires_370_5,addr_370_5);

wire[3:0] wires_371_5;

wire[31:0] addr_371_5;

Selector_2 s371_5(wires_92_4[3], addr_92_4, wires_371_5,addr_371_5);

wire[3:0] wires_372_5;

wire[31:0] addr_372_5;

Selector_2 s372_5(wires_93_4[0], addr_93_4, wires_372_5,addr_372_5);

wire[3:0] wires_373_5;

wire[31:0] addr_373_5;

Selector_2 s373_5(wires_93_4[1], addr_93_4, wires_373_5,addr_373_5);

wire[3:0] wires_374_5;

wire[31:0] addr_374_5;

Selector_2 s374_5(wires_93_4[2], addr_93_4, wires_374_5,addr_374_5);

wire[3:0] wires_375_5;

wire[31:0] addr_375_5;

Selector_2 s375_5(wires_93_4[3], addr_93_4, wires_375_5,addr_375_5);

wire[3:0] wires_376_5;

wire[31:0] addr_376_5;

Selector_2 s376_5(wires_94_4[0], addr_94_4, wires_376_5,addr_376_5);

wire[3:0] wires_377_5;

wire[31:0] addr_377_5;

Selector_2 s377_5(wires_94_4[1], addr_94_4, wires_377_5,addr_377_5);

wire[3:0] wires_378_5;

wire[31:0] addr_378_5;

Selector_2 s378_5(wires_94_4[2], addr_94_4, wires_378_5,addr_378_5);

wire[3:0] wires_379_5;

wire[31:0] addr_379_5;

Selector_2 s379_5(wires_94_4[3], addr_94_4, wires_379_5,addr_379_5);

wire[3:0] wires_380_5;

wire[31:0] addr_380_5;

Selector_2 s380_5(wires_95_4[0], addr_95_4, wires_380_5,addr_380_5);

wire[3:0] wires_381_5;

wire[31:0] addr_381_5;

Selector_2 s381_5(wires_95_4[1], addr_95_4, wires_381_5,addr_381_5);

wire[3:0] wires_382_5;

wire[31:0] addr_382_5;

Selector_2 s382_5(wires_95_4[2], addr_95_4, wires_382_5,addr_382_5);

wire[3:0] wires_383_5;

wire[31:0] addr_383_5;

Selector_2 s383_5(wires_95_4[3], addr_95_4, wires_383_5,addr_383_5);

wire[3:0] wires_384_5;

wire[31:0] addr_384_5;

Selector_2 s384_5(wires_96_4[0], addr_96_4, wires_384_5,addr_384_5);

wire[3:0] wires_385_5;

wire[31:0] addr_385_5;

Selector_2 s385_5(wires_96_4[1], addr_96_4, wires_385_5,addr_385_5);

wire[3:0] wires_386_5;

wire[31:0] addr_386_5;

Selector_2 s386_5(wires_96_4[2], addr_96_4, wires_386_5,addr_386_5);

wire[3:0] wires_387_5;

wire[31:0] addr_387_5;

Selector_2 s387_5(wires_96_4[3], addr_96_4, wires_387_5,addr_387_5);

wire[3:0] wires_388_5;

wire[31:0] addr_388_5;

Selector_2 s388_5(wires_97_4[0], addr_97_4, wires_388_5,addr_388_5);

wire[3:0] wires_389_5;

wire[31:0] addr_389_5;

Selector_2 s389_5(wires_97_4[1], addr_97_4, wires_389_5,addr_389_5);

wire[3:0] wires_390_5;

wire[31:0] addr_390_5;

Selector_2 s390_5(wires_97_4[2], addr_97_4, wires_390_5,addr_390_5);

wire[3:0] wires_391_5;

wire[31:0] addr_391_5;

Selector_2 s391_5(wires_97_4[3], addr_97_4, wires_391_5,addr_391_5);

wire[3:0] wires_392_5;

wire[31:0] addr_392_5;

Selector_2 s392_5(wires_98_4[0], addr_98_4, wires_392_5,addr_392_5);

wire[3:0] wires_393_5;

wire[31:0] addr_393_5;

Selector_2 s393_5(wires_98_4[1], addr_98_4, wires_393_5,addr_393_5);

wire[3:0] wires_394_5;

wire[31:0] addr_394_5;

Selector_2 s394_5(wires_98_4[2], addr_98_4, wires_394_5,addr_394_5);

wire[3:0] wires_395_5;

wire[31:0] addr_395_5;

Selector_2 s395_5(wires_98_4[3], addr_98_4, wires_395_5,addr_395_5);

wire[3:0] wires_396_5;

wire[31:0] addr_396_5;

Selector_2 s396_5(wires_99_4[0], addr_99_4, wires_396_5,addr_396_5);

wire[3:0] wires_397_5;

wire[31:0] addr_397_5;

Selector_2 s397_5(wires_99_4[1], addr_99_4, wires_397_5,addr_397_5);

wire[3:0] wires_398_5;

wire[31:0] addr_398_5;

Selector_2 s398_5(wires_99_4[2], addr_99_4, wires_398_5,addr_398_5);

wire[3:0] wires_399_5;

wire[31:0] addr_399_5;

Selector_2 s399_5(wires_99_4[3], addr_99_4, wires_399_5,addr_399_5);

wire[3:0] wires_400_5;

wire[31:0] addr_400_5;

Selector_2 s400_5(wires_100_4[0], addr_100_4, wires_400_5,addr_400_5);

wire[3:0] wires_401_5;

wire[31:0] addr_401_5;

Selector_2 s401_5(wires_100_4[1], addr_100_4, wires_401_5,addr_401_5);

wire[3:0] wires_402_5;

wire[31:0] addr_402_5;

Selector_2 s402_5(wires_100_4[2], addr_100_4, wires_402_5,addr_402_5);

wire[3:0] wires_403_5;

wire[31:0] addr_403_5;

Selector_2 s403_5(wires_100_4[3], addr_100_4, wires_403_5,addr_403_5);

wire[3:0] wires_404_5;

wire[31:0] addr_404_5;

Selector_2 s404_5(wires_101_4[0], addr_101_4, wires_404_5,addr_404_5);

wire[3:0] wires_405_5;

wire[31:0] addr_405_5;

Selector_2 s405_5(wires_101_4[1], addr_101_4, wires_405_5,addr_405_5);

wire[3:0] wires_406_5;

wire[31:0] addr_406_5;

Selector_2 s406_5(wires_101_4[2], addr_101_4, wires_406_5,addr_406_5);

wire[3:0] wires_407_5;

wire[31:0] addr_407_5;

Selector_2 s407_5(wires_101_4[3], addr_101_4, wires_407_5,addr_407_5);

wire[3:0] wires_408_5;

wire[31:0] addr_408_5;

Selector_2 s408_5(wires_102_4[0], addr_102_4, wires_408_5,addr_408_5);

wire[3:0] wires_409_5;

wire[31:0] addr_409_5;

Selector_2 s409_5(wires_102_4[1], addr_102_4, wires_409_5,addr_409_5);

wire[3:0] wires_410_5;

wire[31:0] addr_410_5;

Selector_2 s410_5(wires_102_4[2], addr_102_4, wires_410_5,addr_410_5);

wire[3:0] wires_411_5;

wire[31:0] addr_411_5;

Selector_2 s411_5(wires_102_4[3], addr_102_4, wires_411_5,addr_411_5);

wire[3:0] wires_412_5;

wire[31:0] addr_412_5;

Selector_2 s412_5(wires_103_4[0], addr_103_4, wires_412_5,addr_412_5);

wire[3:0] wires_413_5;

wire[31:0] addr_413_5;

Selector_2 s413_5(wires_103_4[1], addr_103_4, wires_413_5,addr_413_5);

wire[3:0] wires_414_5;

wire[31:0] addr_414_5;

Selector_2 s414_5(wires_103_4[2], addr_103_4, wires_414_5,addr_414_5);

wire[3:0] wires_415_5;

wire[31:0] addr_415_5;

Selector_2 s415_5(wires_103_4[3], addr_103_4, wires_415_5,addr_415_5);

wire[3:0] wires_416_5;

wire[31:0] addr_416_5;

Selector_2 s416_5(wires_104_4[0], addr_104_4, wires_416_5,addr_416_5);

wire[3:0] wires_417_5;

wire[31:0] addr_417_5;

Selector_2 s417_5(wires_104_4[1], addr_104_4, wires_417_5,addr_417_5);

wire[3:0] wires_418_5;

wire[31:0] addr_418_5;

Selector_2 s418_5(wires_104_4[2], addr_104_4, wires_418_5,addr_418_5);

wire[3:0] wires_419_5;

wire[31:0] addr_419_5;

Selector_2 s419_5(wires_104_4[3], addr_104_4, wires_419_5,addr_419_5);

wire[3:0] wires_420_5;

wire[31:0] addr_420_5;

Selector_2 s420_5(wires_105_4[0], addr_105_4, wires_420_5,addr_420_5);

wire[3:0] wires_421_5;

wire[31:0] addr_421_5;

Selector_2 s421_5(wires_105_4[1], addr_105_4, wires_421_5,addr_421_5);

wire[3:0] wires_422_5;

wire[31:0] addr_422_5;

Selector_2 s422_5(wires_105_4[2], addr_105_4, wires_422_5,addr_422_5);

wire[3:0] wires_423_5;

wire[31:0] addr_423_5;

Selector_2 s423_5(wires_105_4[3], addr_105_4, wires_423_5,addr_423_5);

wire[3:0] wires_424_5;

wire[31:0] addr_424_5;

Selector_2 s424_5(wires_106_4[0], addr_106_4, wires_424_5,addr_424_5);

wire[3:0] wires_425_5;

wire[31:0] addr_425_5;

Selector_2 s425_5(wires_106_4[1], addr_106_4, wires_425_5,addr_425_5);

wire[3:0] wires_426_5;

wire[31:0] addr_426_5;

Selector_2 s426_5(wires_106_4[2], addr_106_4, wires_426_5,addr_426_5);

wire[3:0] wires_427_5;

wire[31:0] addr_427_5;

Selector_2 s427_5(wires_106_4[3], addr_106_4, wires_427_5,addr_427_5);

wire[3:0] wires_428_5;

wire[31:0] addr_428_5;

Selector_2 s428_5(wires_107_4[0], addr_107_4, wires_428_5,addr_428_5);

wire[3:0] wires_429_5;

wire[31:0] addr_429_5;

Selector_2 s429_5(wires_107_4[1], addr_107_4, wires_429_5,addr_429_5);

wire[3:0] wires_430_5;

wire[31:0] addr_430_5;

Selector_2 s430_5(wires_107_4[2], addr_107_4, wires_430_5,addr_430_5);

wire[3:0] wires_431_5;

wire[31:0] addr_431_5;

Selector_2 s431_5(wires_107_4[3], addr_107_4, wires_431_5,addr_431_5);

wire[3:0] wires_432_5;

wire[31:0] addr_432_5;

Selector_2 s432_5(wires_108_4[0], addr_108_4, wires_432_5,addr_432_5);

wire[3:0] wires_433_5;

wire[31:0] addr_433_5;

Selector_2 s433_5(wires_108_4[1], addr_108_4, wires_433_5,addr_433_5);

wire[3:0] wires_434_5;

wire[31:0] addr_434_5;

Selector_2 s434_5(wires_108_4[2], addr_108_4, wires_434_5,addr_434_5);

wire[3:0] wires_435_5;

wire[31:0] addr_435_5;

Selector_2 s435_5(wires_108_4[3], addr_108_4, wires_435_5,addr_435_5);

wire[3:0] wires_436_5;

wire[31:0] addr_436_5;

Selector_2 s436_5(wires_109_4[0], addr_109_4, wires_436_5,addr_436_5);

wire[3:0] wires_437_5;

wire[31:0] addr_437_5;

Selector_2 s437_5(wires_109_4[1], addr_109_4, wires_437_5,addr_437_5);

wire[3:0] wires_438_5;

wire[31:0] addr_438_5;

Selector_2 s438_5(wires_109_4[2], addr_109_4, wires_438_5,addr_438_5);

wire[3:0] wires_439_5;

wire[31:0] addr_439_5;

Selector_2 s439_5(wires_109_4[3], addr_109_4, wires_439_5,addr_439_5);

wire[3:0] wires_440_5;

wire[31:0] addr_440_5;

Selector_2 s440_5(wires_110_4[0], addr_110_4, wires_440_5,addr_440_5);

wire[3:0] wires_441_5;

wire[31:0] addr_441_5;

Selector_2 s441_5(wires_110_4[1], addr_110_4, wires_441_5,addr_441_5);

wire[3:0] wires_442_5;

wire[31:0] addr_442_5;

Selector_2 s442_5(wires_110_4[2], addr_110_4, wires_442_5,addr_442_5);

wire[3:0] wires_443_5;

wire[31:0] addr_443_5;

Selector_2 s443_5(wires_110_4[3], addr_110_4, wires_443_5,addr_443_5);

wire[3:0] wires_444_5;

wire[31:0] addr_444_5;

Selector_2 s444_5(wires_111_4[0], addr_111_4, wires_444_5,addr_444_5);

wire[3:0] wires_445_5;

wire[31:0] addr_445_5;

Selector_2 s445_5(wires_111_4[1], addr_111_4, wires_445_5,addr_445_5);

wire[3:0] wires_446_5;

wire[31:0] addr_446_5;

Selector_2 s446_5(wires_111_4[2], addr_111_4, wires_446_5,addr_446_5);

wire[3:0] wires_447_5;

wire[31:0] addr_447_5;

Selector_2 s447_5(wires_111_4[3], addr_111_4, wires_447_5,addr_447_5);

wire[3:0] wires_448_5;

wire[31:0] addr_448_5;

Selector_2 s448_5(wires_112_4[0], addr_112_4, wires_448_5,addr_448_5);

wire[3:0] wires_449_5;

wire[31:0] addr_449_5;

Selector_2 s449_5(wires_112_4[1], addr_112_4, wires_449_5,addr_449_5);

wire[3:0] wires_450_5;

wire[31:0] addr_450_5;

Selector_2 s450_5(wires_112_4[2], addr_112_4, wires_450_5,addr_450_5);

wire[3:0] wires_451_5;

wire[31:0] addr_451_5;

Selector_2 s451_5(wires_112_4[3], addr_112_4, wires_451_5,addr_451_5);

wire[3:0] wires_452_5;

wire[31:0] addr_452_5;

Selector_2 s452_5(wires_113_4[0], addr_113_4, wires_452_5,addr_452_5);

wire[3:0] wires_453_5;

wire[31:0] addr_453_5;

Selector_2 s453_5(wires_113_4[1], addr_113_4, wires_453_5,addr_453_5);

wire[3:0] wires_454_5;

wire[31:0] addr_454_5;

Selector_2 s454_5(wires_113_4[2], addr_113_4, wires_454_5,addr_454_5);

wire[3:0] wires_455_5;

wire[31:0] addr_455_5;

Selector_2 s455_5(wires_113_4[3], addr_113_4, wires_455_5,addr_455_5);

wire[3:0] wires_456_5;

wire[31:0] addr_456_5;

Selector_2 s456_5(wires_114_4[0], addr_114_4, wires_456_5,addr_456_5);

wire[3:0] wires_457_5;

wire[31:0] addr_457_5;

Selector_2 s457_5(wires_114_4[1], addr_114_4, wires_457_5,addr_457_5);

wire[3:0] wires_458_5;

wire[31:0] addr_458_5;

Selector_2 s458_5(wires_114_4[2], addr_114_4, wires_458_5,addr_458_5);

wire[3:0] wires_459_5;

wire[31:0] addr_459_5;

Selector_2 s459_5(wires_114_4[3], addr_114_4, wires_459_5,addr_459_5);

wire[3:0] wires_460_5;

wire[31:0] addr_460_5;

Selector_2 s460_5(wires_115_4[0], addr_115_4, wires_460_5,addr_460_5);

wire[3:0] wires_461_5;

wire[31:0] addr_461_5;

Selector_2 s461_5(wires_115_4[1], addr_115_4, wires_461_5,addr_461_5);

wire[3:0] wires_462_5;

wire[31:0] addr_462_5;

Selector_2 s462_5(wires_115_4[2], addr_115_4, wires_462_5,addr_462_5);

wire[3:0] wires_463_5;

wire[31:0] addr_463_5;

Selector_2 s463_5(wires_115_4[3], addr_115_4, wires_463_5,addr_463_5);

wire[3:0] wires_464_5;

wire[31:0] addr_464_5;

Selector_2 s464_5(wires_116_4[0], addr_116_4, wires_464_5,addr_464_5);

wire[3:0] wires_465_5;

wire[31:0] addr_465_5;

Selector_2 s465_5(wires_116_4[1], addr_116_4, wires_465_5,addr_465_5);

wire[3:0] wires_466_5;

wire[31:0] addr_466_5;

Selector_2 s466_5(wires_116_4[2], addr_116_4, wires_466_5,addr_466_5);

wire[3:0] wires_467_5;

wire[31:0] addr_467_5;

Selector_2 s467_5(wires_116_4[3], addr_116_4, wires_467_5,addr_467_5);

wire[3:0] wires_468_5;

wire[31:0] addr_468_5;

Selector_2 s468_5(wires_117_4[0], addr_117_4, wires_468_5,addr_468_5);

wire[3:0] wires_469_5;

wire[31:0] addr_469_5;

Selector_2 s469_5(wires_117_4[1], addr_117_4, wires_469_5,addr_469_5);

wire[3:0] wires_470_5;

wire[31:0] addr_470_5;

Selector_2 s470_5(wires_117_4[2], addr_117_4, wires_470_5,addr_470_5);

wire[3:0] wires_471_5;

wire[31:0] addr_471_5;

Selector_2 s471_5(wires_117_4[3], addr_117_4, wires_471_5,addr_471_5);

wire[3:0] wires_472_5;

wire[31:0] addr_472_5;

Selector_2 s472_5(wires_118_4[0], addr_118_4, wires_472_5,addr_472_5);

wire[3:0] wires_473_5;

wire[31:0] addr_473_5;

Selector_2 s473_5(wires_118_4[1], addr_118_4, wires_473_5,addr_473_5);

wire[3:0] wires_474_5;

wire[31:0] addr_474_5;

Selector_2 s474_5(wires_118_4[2], addr_118_4, wires_474_5,addr_474_5);

wire[3:0] wires_475_5;

wire[31:0] addr_475_5;

Selector_2 s475_5(wires_118_4[3], addr_118_4, wires_475_5,addr_475_5);

wire[3:0] wires_476_5;

wire[31:0] addr_476_5;

Selector_2 s476_5(wires_119_4[0], addr_119_4, wires_476_5,addr_476_5);

wire[3:0] wires_477_5;

wire[31:0] addr_477_5;

Selector_2 s477_5(wires_119_4[1], addr_119_4, wires_477_5,addr_477_5);

wire[3:0] wires_478_5;

wire[31:0] addr_478_5;

Selector_2 s478_5(wires_119_4[2], addr_119_4, wires_478_5,addr_478_5);

wire[3:0] wires_479_5;

wire[31:0] addr_479_5;

Selector_2 s479_5(wires_119_4[3], addr_119_4, wires_479_5,addr_479_5);

wire[3:0] wires_480_5;

wire[31:0] addr_480_5;

Selector_2 s480_5(wires_120_4[0], addr_120_4, wires_480_5,addr_480_5);

wire[3:0] wires_481_5;

wire[31:0] addr_481_5;

Selector_2 s481_5(wires_120_4[1], addr_120_4, wires_481_5,addr_481_5);

wire[3:0] wires_482_5;

wire[31:0] addr_482_5;

Selector_2 s482_5(wires_120_4[2], addr_120_4, wires_482_5,addr_482_5);

wire[3:0] wires_483_5;

wire[31:0] addr_483_5;

Selector_2 s483_5(wires_120_4[3], addr_120_4, wires_483_5,addr_483_5);

wire[3:0] wires_484_5;

wire[31:0] addr_484_5;

Selector_2 s484_5(wires_121_4[0], addr_121_4, wires_484_5,addr_484_5);

wire[3:0] wires_485_5;

wire[31:0] addr_485_5;

Selector_2 s485_5(wires_121_4[1], addr_121_4, wires_485_5,addr_485_5);

wire[3:0] wires_486_5;

wire[31:0] addr_486_5;

Selector_2 s486_5(wires_121_4[2], addr_121_4, wires_486_5,addr_486_5);

wire[3:0] wires_487_5;

wire[31:0] addr_487_5;

Selector_2 s487_5(wires_121_4[3], addr_121_4, wires_487_5,addr_487_5);

wire[3:0] wires_488_5;

wire[31:0] addr_488_5;

Selector_2 s488_5(wires_122_4[0], addr_122_4, wires_488_5,addr_488_5);

wire[3:0] wires_489_5;

wire[31:0] addr_489_5;

Selector_2 s489_5(wires_122_4[1], addr_122_4, wires_489_5,addr_489_5);

wire[3:0] wires_490_5;

wire[31:0] addr_490_5;

Selector_2 s490_5(wires_122_4[2], addr_122_4, wires_490_5,addr_490_5);

wire[3:0] wires_491_5;

wire[31:0] addr_491_5;

Selector_2 s491_5(wires_122_4[3], addr_122_4, wires_491_5,addr_491_5);

wire[3:0] wires_492_5;

wire[31:0] addr_492_5;

Selector_2 s492_5(wires_123_4[0], addr_123_4, wires_492_5,addr_492_5);

wire[3:0] wires_493_5;

wire[31:0] addr_493_5;

Selector_2 s493_5(wires_123_4[1], addr_123_4, wires_493_5,addr_493_5);

wire[3:0] wires_494_5;

wire[31:0] addr_494_5;

Selector_2 s494_5(wires_123_4[2], addr_123_4, wires_494_5,addr_494_5);

wire[3:0] wires_495_5;

wire[31:0] addr_495_5;

Selector_2 s495_5(wires_123_4[3], addr_123_4, wires_495_5,addr_495_5);

wire[3:0] wires_496_5;

wire[31:0] addr_496_5;

Selector_2 s496_5(wires_124_4[0], addr_124_4, wires_496_5,addr_496_5);

wire[3:0] wires_497_5;

wire[31:0] addr_497_5;

Selector_2 s497_5(wires_124_4[1], addr_124_4, wires_497_5,addr_497_5);

wire[3:0] wires_498_5;

wire[31:0] addr_498_5;

Selector_2 s498_5(wires_124_4[2], addr_124_4, wires_498_5,addr_498_5);

wire[3:0] wires_499_5;

wire[31:0] addr_499_5;

Selector_2 s499_5(wires_124_4[3], addr_124_4, wires_499_5,addr_499_5);

wire[3:0] wires_500_5;

wire[31:0] addr_500_5;

Selector_2 s500_5(wires_125_4[0], addr_125_4, wires_500_5,addr_500_5);

wire[3:0] wires_501_5;

wire[31:0] addr_501_5;

Selector_2 s501_5(wires_125_4[1], addr_125_4, wires_501_5,addr_501_5);

wire[3:0] wires_502_5;

wire[31:0] addr_502_5;

Selector_2 s502_5(wires_125_4[2], addr_125_4, wires_502_5,addr_502_5);

wire[3:0] wires_503_5;

wire[31:0] addr_503_5;

Selector_2 s503_5(wires_125_4[3], addr_125_4, wires_503_5,addr_503_5);

wire[3:0] wires_504_5;

wire[31:0] addr_504_5;

Selector_2 s504_5(wires_126_4[0], addr_126_4, wires_504_5,addr_504_5);

wire[3:0] wires_505_5;

wire[31:0] addr_505_5;

Selector_2 s505_5(wires_126_4[1], addr_126_4, wires_505_5,addr_505_5);

wire[3:0] wires_506_5;

wire[31:0] addr_506_5;

Selector_2 s506_5(wires_126_4[2], addr_126_4, wires_506_5,addr_506_5);

wire[3:0] wires_507_5;

wire[31:0] addr_507_5;

Selector_2 s507_5(wires_126_4[3], addr_126_4, wires_507_5,addr_507_5);

wire[3:0] wires_508_5;

wire[31:0] addr_508_5;

Selector_2 s508_5(wires_127_4[0], addr_127_4, wires_508_5,addr_508_5);

wire[3:0] wires_509_5;

wire[31:0] addr_509_5;

Selector_2 s509_5(wires_127_4[1], addr_127_4, wires_509_5,addr_509_5);

wire[3:0] wires_510_5;

wire[31:0] addr_510_5;

Selector_2 s510_5(wires_127_4[2], addr_127_4, wires_510_5,addr_510_5);

wire[3:0] wires_511_5;

wire[31:0] addr_511_5;

Selector_2 s511_5(wires_127_4[3], addr_127_4, wires_511_5,addr_511_5);

wire[3:0] wires_512_5;

wire[31:0] addr_512_5;

Selector_2 s512_5(wires_128_4[0], addr_128_4, wires_512_5,addr_512_5);

wire[3:0] wires_513_5;

wire[31:0] addr_513_5;

Selector_2 s513_5(wires_128_4[1], addr_128_4, wires_513_5,addr_513_5);

wire[3:0] wires_514_5;

wire[31:0] addr_514_5;

Selector_2 s514_5(wires_128_4[2], addr_128_4, wires_514_5,addr_514_5);

wire[3:0] wires_515_5;

wire[31:0] addr_515_5;

Selector_2 s515_5(wires_128_4[3], addr_128_4, wires_515_5,addr_515_5);

wire[3:0] wires_516_5;

wire[31:0] addr_516_5;

Selector_2 s516_5(wires_129_4[0], addr_129_4, wires_516_5,addr_516_5);

wire[3:0] wires_517_5;

wire[31:0] addr_517_5;

Selector_2 s517_5(wires_129_4[1], addr_129_4, wires_517_5,addr_517_5);

wire[3:0] wires_518_5;

wire[31:0] addr_518_5;

Selector_2 s518_5(wires_129_4[2], addr_129_4, wires_518_5,addr_518_5);

wire[3:0] wires_519_5;

wire[31:0] addr_519_5;

Selector_2 s519_5(wires_129_4[3], addr_129_4, wires_519_5,addr_519_5);

wire[3:0] wires_520_5;

wire[31:0] addr_520_5;

Selector_2 s520_5(wires_130_4[0], addr_130_4, wires_520_5,addr_520_5);

wire[3:0] wires_521_5;

wire[31:0] addr_521_5;

Selector_2 s521_5(wires_130_4[1], addr_130_4, wires_521_5,addr_521_5);

wire[3:0] wires_522_5;

wire[31:0] addr_522_5;

Selector_2 s522_5(wires_130_4[2], addr_130_4, wires_522_5,addr_522_5);

wire[3:0] wires_523_5;

wire[31:0] addr_523_5;

Selector_2 s523_5(wires_130_4[3], addr_130_4, wires_523_5,addr_523_5);

wire[3:0] wires_524_5;

wire[31:0] addr_524_5;

Selector_2 s524_5(wires_131_4[0], addr_131_4, wires_524_5,addr_524_5);

wire[3:0] wires_525_5;

wire[31:0] addr_525_5;

Selector_2 s525_5(wires_131_4[1], addr_131_4, wires_525_5,addr_525_5);

wire[3:0] wires_526_5;

wire[31:0] addr_526_5;

Selector_2 s526_5(wires_131_4[2], addr_131_4, wires_526_5,addr_526_5);

wire[3:0] wires_527_5;

wire[31:0] addr_527_5;

Selector_2 s527_5(wires_131_4[3], addr_131_4, wires_527_5,addr_527_5);

wire[3:0] wires_528_5;

wire[31:0] addr_528_5;

Selector_2 s528_5(wires_132_4[0], addr_132_4, wires_528_5,addr_528_5);

wire[3:0] wires_529_5;

wire[31:0] addr_529_5;

Selector_2 s529_5(wires_132_4[1], addr_132_4, wires_529_5,addr_529_5);

wire[3:0] wires_530_5;

wire[31:0] addr_530_5;

Selector_2 s530_5(wires_132_4[2], addr_132_4, wires_530_5,addr_530_5);

wire[3:0] wires_531_5;

wire[31:0] addr_531_5;

Selector_2 s531_5(wires_132_4[3], addr_132_4, wires_531_5,addr_531_5);

wire[3:0] wires_532_5;

wire[31:0] addr_532_5;

Selector_2 s532_5(wires_133_4[0], addr_133_4, wires_532_5,addr_532_5);

wire[3:0] wires_533_5;

wire[31:0] addr_533_5;

Selector_2 s533_5(wires_133_4[1], addr_133_4, wires_533_5,addr_533_5);

wire[3:0] wires_534_5;

wire[31:0] addr_534_5;

Selector_2 s534_5(wires_133_4[2], addr_133_4, wires_534_5,addr_534_5);

wire[3:0] wires_535_5;

wire[31:0] addr_535_5;

Selector_2 s535_5(wires_133_4[3], addr_133_4, wires_535_5,addr_535_5);

wire[3:0] wires_536_5;

wire[31:0] addr_536_5;

Selector_2 s536_5(wires_134_4[0], addr_134_4, wires_536_5,addr_536_5);

wire[3:0] wires_537_5;

wire[31:0] addr_537_5;

Selector_2 s537_5(wires_134_4[1], addr_134_4, wires_537_5,addr_537_5);

wire[3:0] wires_538_5;

wire[31:0] addr_538_5;

Selector_2 s538_5(wires_134_4[2], addr_134_4, wires_538_5,addr_538_5);

wire[3:0] wires_539_5;

wire[31:0] addr_539_5;

Selector_2 s539_5(wires_134_4[3], addr_134_4, wires_539_5,addr_539_5);

wire[3:0] wires_540_5;

wire[31:0] addr_540_5;

Selector_2 s540_5(wires_135_4[0], addr_135_4, wires_540_5,addr_540_5);

wire[3:0] wires_541_5;

wire[31:0] addr_541_5;

Selector_2 s541_5(wires_135_4[1], addr_135_4, wires_541_5,addr_541_5);

wire[3:0] wires_542_5;

wire[31:0] addr_542_5;

Selector_2 s542_5(wires_135_4[2], addr_135_4, wires_542_5,addr_542_5);

wire[3:0] wires_543_5;

wire[31:0] addr_543_5;

Selector_2 s543_5(wires_135_4[3], addr_135_4, wires_543_5,addr_543_5);

wire[3:0] wires_544_5;

wire[31:0] addr_544_5;

Selector_2 s544_5(wires_136_4[0], addr_136_4, wires_544_5,addr_544_5);

wire[3:0] wires_545_5;

wire[31:0] addr_545_5;

Selector_2 s545_5(wires_136_4[1], addr_136_4, wires_545_5,addr_545_5);

wire[3:0] wires_546_5;

wire[31:0] addr_546_5;

Selector_2 s546_5(wires_136_4[2], addr_136_4, wires_546_5,addr_546_5);

wire[3:0] wires_547_5;

wire[31:0] addr_547_5;

Selector_2 s547_5(wires_136_4[3], addr_136_4, wires_547_5,addr_547_5);

wire[3:0] wires_548_5;

wire[31:0] addr_548_5;

Selector_2 s548_5(wires_137_4[0], addr_137_4, wires_548_5,addr_548_5);

wire[3:0] wires_549_5;

wire[31:0] addr_549_5;

Selector_2 s549_5(wires_137_4[1], addr_137_4, wires_549_5,addr_549_5);

wire[3:0] wires_550_5;

wire[31:0] addr_550_5;

Selector_2 s550_5(wires_137_4[2], addr_137_4, wires_550_5,addr_550_5);

wire[3:0] wires_551_5;

wire[31:0] addr_551_5;

Selector_2 s551_5(wires_137_4[3], addr_137_4, wires_551_5,addr_551_5);

wire[3:0] wires_552_5;

wire[31:0] addr_552_5;

Selector_2 s552_5(wires_138_4[0], addr_138_4, wires_552_5,addr_552_5);

wire[3:0] wires_553_5;

wire[31:0] addr_553_5;

Selector_2 s553_5(wires_138_4[1], addr_138_4, wires_553_5,addr_553_5);

wire[3:0] wires_554_5;

wire[31:0] addr_554_5;

Selector_2 s554_5(wires_138_4[2], addr_138_4, wires_554_5,addr_554_5);

wire[3:0] wires_555_5;

wire[31:0] addr_555_5;

Selector_2 s555_5(wires_138_4[3], addr_138_4, wires_555_5,addr_555_5);

wire[3:0] wires_556_5;

wire[31:0] addr_556_5;

Selector_2 s556_5(wires_139_4[0], addr_139_4, wires_556_5,addr_556_5);

wire[3:0] wires_557_5;

wire[31:0] addr_557_5;

Selector_2 s557_5(wires_139_4[1], addr_139_4, wires_557_5,addr_557_5);

wire[3:0] wires_558_5;

wire[31:0] addr_558_5;

Selector_2 s558_5(wires_139_4[2], addr_139_4, wires_558_5,addr_558_5);

wire[3:0] wires_559_5;

wire[31:0] addr_559_5;

Selector_2 s559_5(wires_139_4[3], addr_139_4, wires_559_5,addr_559_5);

wire[3:0] wires_560_5;

wire[31:0] addr_560_5;

Selector_2 s560_5(wires_140_4[0], addr_140_4, wires_560_5,addr_560_5);

wire[3:0] wires_561_5;

wire[31:0] addr_561_5;

Selector_2 s561_5(wires_140_4[1], addr_140_4, wires_561_5,addr_561_5);

wire[3:0] wires_562_5;

wire[31:0] addr_562_5;

Selector_2 s562_5(wires_140_4[2], addr_140_4, wires_562_5,addr_562_5);

wire[3:0] wires_563_5;

wire[31:0] addr_563_5;

Selector_2 s563_5(wires_140_4[3], addr_140_4, wires_563_5,addr_563_5);

wire[3:0] wires_564_5;

wire[31:0] addr_564_5;

Selector_2 s564_5(wires_141_4[0], addr_141_4, wires_564_5,addr_564_5);

wire[3:0] wires_565_5;

wire[31:0] addr_565_5;

Selector_2 s565_5(wires_141_4[1], addr_141_4, wires_565_5,addr_565_5);

wire[3:0] wires_566_5;

wire[31:0] addr_566_5;

Selector_2 s566_5(wires_141_4[2], addr_141_4, wires_566_5,addr_566_5);

wire[3:0] wires_567_5;

wire[31:0] addr_567_5;

Selector_2 s567_5(wires_141_4[3], addr_141_4, wires_567_5,addr_567_5);

wire[3:0] wires_568_5;

wire[31:0] addr_568_5;

Selector_2 s568_5(wires_142_4[0], addr_142_4, wires_568_5,addr_568_5);

wire[3:0] wires_569_5;

wire[31:0] addr_569_5;

Selector_2 s569_5(wires_142_4[1], addr_142_4, wires_569_5,addr_569_5);

wire[3:0] wires_570_5;

wire[31:0] addr_570_5;

Selector_2 s570_5(wires_142_4[2], addr_142_4, wires_570_5,addr_570_5);

wire[3:0] wires_571_5;

wire[31:0] addr_571_5;

Selector_2 s571_5(wires_142_4[3], addr_142_4, wires_571_5,addr_571_5);

wire[3:0] wires_572_5;

wire[31:0] addr_572_5;

Selector_2 s572_5(wires_143_4[0], addr_143_4, wires_572_5,addr_572_5);

wire[3:0] wires_573_5;

wire[31:0] addr_573_5;

Selector_2 s573_5(wires_143_4[1], addr_143_4, wires_573_5,addr_573_5);

wire[3:0] wires_574_5;

wire[31:0] addr_574_5;

Selector_2 s574_5(wires_143_4[2], addr_143_4, wires_574_5,addr_574_5);

wire[3:0] wires_575_5;

wire[31:0] addr_575_5;

Selector_2 s575_5(wires_143_4[3], addr_143_4, wires_575_5,addr_575_5);

wire[3:0] wires_576_5;

wire[31:0] addr_576_5;

Selector_2 s576_5(wires_144_4[0], addr_144_4, wires_576_5,addr_576_5);

wire[3:0] wires_577_5;

wire[31:0] addr_577_5;

Selector_2 s577_5(wires_144_4[1], addr_144_4, wires_577_5,addr_577_5);

wire[3:0] wires_578_5;

wire[31:0] addr_578_5;

Selector_2 s578_5(wires_144_4[2], addr_144_4, wires_578_5,addr_578_5);

wire[3:0] wires_579_5;

wire[31:0] addr_579_5;

Selector_2 s579_5(wires_144_4[3], addr_144_4, wires_579_5,addr_579_5);

wire[3:0] wires_580_5;

wire[31:0] addr_580_5;

Selector_2 s580_5(wires_145_4[0], addr_145_4, wires_580_5,addr_580_5);

wire[3:0] wires_581_5;

wire[31:0] addr_581_5;

Selector_2 s581_5(wires_145_4[1], addr_145_4, wires_581_5,addr_581_5);

wire[3:0] wires_582_5;

wire[31:0] addr_582_5;

Selector_2 s582_5(wires_145_4[2], addr_145_4, wires_582_5,addr_582_5);

wire[3:0] wires_583_5;

wire[31:0] addr_583_5;

Selector_2 s583_5(wires_145_4[3], addr_145_4, wires_583_5,addr_583_5);

wire[3:0] wires_584_5;

wire[31:0] addr_584_5;

Selector_2 s584_5(wires_146_4[0], addr_146_4, wires_584_5,addr_584_5);

wire[3:0] wires_585_5;

wire[31:0] addr_585_5;

Selector_2 s585_5(wires_146_4[1], addr_146_4, wires_585_5,addr_585_5);

wire[3:0] wires_586_5;

wire[31:0] addr_586_5;

Selector_2 s586_5(wires_146_4[2], addr_146_4, wires_586_5,addr_586_5);

wire[3:0] wires_587_5;

wire[31:0] addr_587_5;

Selector_2 s587_5(wires_146_4[3], addr_146_4, wires_587_5,addr_587_5);

wire[3:0] wires_588_5;

wire[31:0] addr_588_5;

Selector_2 s588_5(wires_147_4[0], addr_147_4, wires_588_5,addr_588_5);

wire[3:0] wires_589_5;

wire[31:0] addr_589_5;

Selector_2 s589_5(wires_147_4[1], addr_147_4, wires_589_5,addr_589_5);

wire[3:0] wires_590_5;

wire[31:0] addr_590_5;

Selector_2 s590_5(wires_147_4[2], addr_147_4, wires_590_5,addr_590_5);

wire[3:0] wires_591_5;

wire[31:0] addr_591_5;

Selector_2 s591_5(wires_147_4[3], addr_147_4, wires_591_5,addr_591_5);

wire[3:0] wires_592_5;

wire[31:0] addr_592_5;

Selector_2 s592_5(wires_148_4[0], addr_148_4, wires_592_5,addr_592_5);

wire[3:0] wires_593_5;

wire[31:0] addr_593_5;

Selector_2 s593_5(wires_148_4[1], addr_148_4, wires_593_5,addr_593_5);

wire[3:0] wires_594_5;

wire[31:0] addr_594_5;

Selector_2 s594_5(wires_148_4[2], addr_148_4, wires_594_5,addr_594_5);

wire[3:0] wires_595_5;

wire[31:0] addr_595_5;

Selector_2 s595_5(wires_148_4[3], addr_148_4, wires_595_5,addr_595_5);

wire[3:0] wires_596_5;

wire[31:0] addr_596_5;

Selector_2 s596_5(wires_149_4[0], addr_149_4, wires_596_5,addr_596_5);

wire[3:0] wires_597_5;

wire[31:0] addr_597_5;

Selector_2 s597_5(wires_149_4[1], addr_149_4, wires_597_5,addr_597_5);

wire[3:0] wires_598_5;

wire[31:0] addr_598_5;

Selector_2 s598_5(wires_149_4[2], addr_149_4, wires_598_5,addr_598_5);

wire[3:0] wires_599_5;

wire[31:0] addr_599_5;

Selector_2 s599_5(wires_149_4[3], addr_149_4, wires_599_5,addr_599_5);

wire[3:0] wires_600_5;

wire[31:0] addr_600_5;

Selector_2 s600_5(wires_150_4[0], addr_150_4, wires_600_5,addr_600_5);

wire[3:0] wires_601_5;

wire[31:0] addr_601_5;

Selector_2 s601_5(wires_150_4[1], addr_150_4, wires_601_5,addr_601_5);

wire[3:0] wires_602_5;

wire[31:0] addr_602_5;

Selector_2 s602_5(wires_150_4[2], addr_150_4, wires_602_5,addr_602_5);

wire[3:0] wires_603_5;

wire[31:0] addr_603_5;

Selector_2 s603_5(wires_150_4[3], addr_150_4, wires_603_5,addr_603_5);

wire[3:0] wires_604_5;

wire[31:0] addr_604_5;

Selector_2 s604_5(wires_151_4[0], addr_151_4, wires_604_5,addr_604_5);

wire[3:0] wires_605_5;

wire[31:0] addr_605_5;

Selector_2 s605_5(wires_151_4[1], addr_151_4, wires_605_5,addr_605_5);

wire[3:0] wires_606_5;

wire[31:0] addr_606_5;

Selector_2 s606_5(wires_151_4[2], addr_151_4, wires_606_5,addr_606_5);

wire[3:0] wires_607_5;

wire[31:0] addr_607_5;

Selector_2 s607_5(wires_151_4[3], addr_151_4, wires_607_5,addr_607_5);

wire[3:0] wires_608_5;

wire[31:0] addr_608_5;

Selector_2 s608_5(wires_152_4[0], addr_152_4, wires_608_5,addr_608_5);

wire[3:0] wires_609_5;

wire[31:0] addr_609_5;

Selector_2 s609_5(wires_152_4[1], addr_152_4, wires_609_5,addr_609_5);

wire[3:0] wires_610_5;

wire[31:0] addr_610_5;

Selector_2 s610_5(wires_152_4[2], addr_152_4, wires_610_5,addr_610_5);

wire[3:0] wires_611_5;

wire[31:0] addr_611_5;

Selector_2 s611_5(wires_152_4[3], addr_152_4, wires_611_5,addr_611_5);

wire[3:0] wires_612_5;

wire[31:0] addr_612_5;

Selector_2 s612_5(wires_153_4[0], addr_153_4, wires_612_5,addr_612_5);

wire[3:0] wires_613_5;

wire[31:0] addr_613_5;

Selector_2 s613_5(wires_153_4[1], addr_153_4, wires_613_5,addr_613_5);

wire[3:0] wires_614_5;

wire[31:0] addr_614_5;

Selector_2 s614_5(wires_153_4[2], addr_153_4, wires_614_5,addr_614_5);

wire[3:0] wires_615_5;

wire[31:0] addr_615_5;

Selector_2 s615_5(wires_153_4[3], addr_153_4, wires_615_5,addr_615_5);

wire[3:0] wires_616_5;

wire[31:0] addr_616_5;

Selector_2 s616_5(wires_154_4[0], addr_154_4, wires_616_5,addr_616_5);

wire[3:0] wires_617_5;

wire[31:0] addr_617_5;

Selector_2 s617_5(wires_154_4[1], addr_154_4, wires_617_5,addr_617_5);

wire[3:0] wires_618_5;

wire[31:0] addr_618_5;

Selector_2 s618_5(wires_154_4[2], addr_154_4, wires_618_5,addr_618_5);

wire[3:0] wires_619_5;

wire[31:0] addr_619_5;

Selector_2 s619_5(wires_154_4[3], addr_154_4, wires_619_5,addr_619_5);

wire[3:0] wires_620_5;

wire[31:0] addr_620_5;

Selector_2 s620_5(wires_155_4[0], addr_155_4, wires_620_5,addr_620_5);

wire[3:0] wires_621_5;

wire[31:0] addr_621_5;

Selector_2 s621_5(wires_155_4[1], addr_155_4, wires_621_5,addr_621_5);

wire[3:0] wires_622_5;

wire[31:0] addr_622_5;

Selector_2 s622_5(wires_155_4[2], addr_155_4, wires_622_5,addr_622_5);

wire[3:0] wires_623_5;

wire[31:0] addr_623_5;

Selector_2 s623_5(wires_155_4[3], addr_155_4, wires_623_5,addr_623_5);

wire[3:0] wires_624_5;

wire[31:0] addr_624_5;

Selector_2 s624_5(wires_156_4[0], addr_156_4, wires_624_5,addr_624_5);

wire[3:0] wires_625_5;

wire[31:0] addr_625_5;

Selector_2 s625_5(wires_156_4[1], addr_156_4, wires_625_5,addr_625_5);

wire[3:0] wires_626_5;

wire[31:0] addr_626_5;

Selector_2 s626_5(wires_156_4[2], addr_156_4, wires_626_5,addr_626_5);

wire[3:0] wires_627_5;

wire[31:0] addr_627_5;

Selector_2 s627_5(wires_156_4[3], addr_156_4, wires_627_5,addr_627_5);

wire[3:0] wires_628_5;

wire[31:0] addr_628_5;

Selector_2 s628_5(wires_157_4[0], addr_157_4, wires_628_5,addr_628_5);

wire[3:0] wires_629_5;

wire[31:0] addr_629_5;

Selector_2 s629_5(wires_157_4[1], addr_157_4, wires_629_5,addr_629_5);

wire[3:0] wires_630_5;

wire[31:0] addr_630_5;

Selector_2 s630_5(wires_157_4[2], addr_157_4, wires_630_5,addr_630_5);

wire[3:0] wires_631_5;

wire[31:0] addr_631_5;

Selector_2 s631_5(wires_157_4[3], addr_157_4, wires_631_5,addr_631_5);

wire[3:0] wires_632_5;

wire[31:0] addr_632_5;

Selector_2 s632_5(wires_158_4[0], addr_158_4, wires_632_5,addr_632_5);

wire[3:0] wires_633_5;

wire[31:0] addr_633_5;

Selector_2 s633_5(wires_158_4[1], addr_158_4, wires_633_5,addr_633_5);

wire[3:0] wires_634_5;

wire[31:0] addr_634_5;

Selector_2 s634_5(wires_158_4[2], addr_158_4, wires_634_5,addr_634_5);

wire[3:0] wires_635_5;

wire[31:0] addr_635_5;

Selector_2 s635_5(wires_158_4[3], addr_158_4, wires_635_5,addr_635_5);

wire[3:0] wires_636_5;

wire[31:0] addr_636_5;

Selector_2 s636_5(wires_159_4[0], addr_159_4, wires_636_5,addr_636_5);

wire[3:0] wires_637_5;

wire[31:0] addr_637_5;

Selector_2 s637_5(wires_159_4[1], addr_159_4, wires_637_5,addr_637_5);

wire[3:0] wires_638_5;

wire[31:0] addr_638_5;

Selector_2 s638_5(wires_159_4[2], addr_159_4, wires_638_5,addr_638_5);

wire[3:0] wires_639_5;

wire[31:0] addr_639_5;

Selector_2 s639_5(wires_159_4[3], addr_159_4, wires_639_5,addr_639_5);

wire[3:0] wires_640_5;

wire[31:0] addr_640_5;

Selector_2 s640_5(wires_160_4[0], addr_160_4, wires_640_5,addr_640_5);

wire[3:0] wires_641_5;

wire[31:0] addr_641_5;

Selector_2 s641_5(wires_160_4[1], addr_160_4, wires_641_5,addr_641_5);

wire[3:0] wires_642_5;

wire[31:0] addr_642_5;

Selector_2 s642_5(wires_160_4[2], addr_160_4, wires_642_5,addr_642_5);

wire[3:0] wires_643_5;

wire[31:0] addr_643_5;

Selector_2 s643_5(wires_160_4[3], addr_160_4, wires_643_5,addr_643_5);

wire[3:0] wires_644_5;

wire[31:0] addr_644_5;

Selector_2 s644_5(wires_161_4[0], addr_161_4, wires_644_5,addr_644_5);

wire[3:0] wires_645_5;

wire[31:0] addr_645_5;

Selector_2 s645_5(wires_161_4[1], addr_161_4, wires_645_5,addr_645_5);

wire[3:0] wires_646_5;

wire[31:0] addr_646_5;

Selector_2 s646_5(wires_161_4[2], addr_161_4, wires_646_5,addr_646_5);

wire[3:0] wires_647_5;

wire[31:0] addr_647_5;

Selector_2 s647_5(wires_161_4[3], addr_161_4, wires_647_5,addr_647_5);

wire[3:0] wires_648_5;

wire[31:0] addr_648_5;

Selector_2 s648_5(wires_162_4[0], addr_162_4, wires_648_5,addr_648_5);

wire[3:0] wires_649_5;

wire[31:0] addr_649_5;

Selector_2 s649_5(wires_162_4[1], addr_162_4, wires_649_5,addr_649_5);

wire[3:0] wires_650_5;

wire[31:0] addr_650_5;

Selector_2 s650_5(wires_162_4[2], addr_162_4, wires_650_5,addr_650_5);

wire[3:0] wires_651_5;

wire[31:0] addr_651_5;

Selector_2 s651_5(wires_162_4[3], addr_162_4, wires_651_5,addr_651_5);

wire[3:0] wires_652_5;

wire[31:0] addr_652_5;

Selector_2 s652_5(wires_163_4[0], addr_163_4, wires_652_5,addr_652_5);

wire[3:0] wires_653_5;

wire[31:0] addr_653_5;

Selector_2 s653_5(wires_163_4[1], addr_163_4, wires_653_5,addr_653_5);

wire[3:0] wires_654_5;

wire[31:0] addr_654_5;

Selector_2 s654_5(wires_163_4[2], addr_163_4, wires_654_5,addr_654_5);

wire[3:0] wires_655_5;

wire[31:0] addr_655_5;

Selector_2 s655_5(wires_163_4[3], addr_163_4, wires_655_5,addr_655_5);

wire[3:0] wires_656_5;

wire[31:0] addr_656_5;

Selector_2 s656_5(wires_164_4[0], addr_164_4, wires_656_5,addr_656_5);

wire[3:0] wires_657_5;

wire[31:0] addr_657_5;

Selector_2 s657_5(wires_164_4[1], addr_164_4, wires_657_5,addr_657_5);

wire[3:0] wires_658_5;

wire[31:0] addr_658_5;

Selector_2 s658_5(wires_164_4[2], addr_164_4, wires_658_5,addr_658_5);

wire[3:0] wires_659_5;

wire[31:0] addr_659_5;

Selector_2 s659_5(wires_164_4[3], addr_164_4, wires_659_5,addr_659_5);

wire[3:0] wires_660_5;

wire[31:0] addr_660_5;

Selector_2 s660_5(wires_165_4[0], addr_165_4, wires_660_5,addr_660_5);

wire[3:0] wires_661_5;

wire[31:0] addr_661_5;

Selector_2 s661_5(wires_165_4[1], addr_165_4, wires_661_5,addr_661_5);

wire[3:0] wires_662_5;

wire[31:0] addr_662_5;

Selector_2 s662_5(wires_165_4[2], addr_165_4, wires_662_5,addr_662_5);

wire[3:0] wires_663_5;

wire[31:0] addr_663_5;

Selector_2 s663_5(wires_165_4[3], addr_165_4, wires_663_5,addr_663_5);

wire[3:0] wires_664_5;

wire[31:0] addr_664_5;

Selector_2 s664_5(wires_166_4[0], addr_166_4, wires_664_5,addr_664_5);

wire[3:0] wires_665_5;

wire[31:0] addr_665_5;

Selector_2 s665_5(wires_166_4[1], addr_166_4, wires_665_5,addr_665_5);

wire[3:0] wires_666_5;

wire[31:0] addr_666_5;

Selector_2 s666_5(wires_166_4[2], addr_166_4, wires_666_5,addr_666_5);

wire[3:0] wires_667_5;

wire[31:0] addr_667_5;

Selector_2 s667_5(wires_166_4[3], addr_166_4, wires_667_5,addr_667_5);

wire[3:0] wires_668_5;

wire[31:0] addr_668_5;

Selector_2 s668_5(wires_167_4[0], addr_167_4, wires_668_5,addr_668_5);

wire[3:0] wires_669_5;

wire[31:0] addr_669_5;

Selector_2 s669_5(wires_167_4[1], addr_167_4, wires_669_5,addr_669_5);

wire[3:0] wires_670_5;

wire[31:0] addr_670_5;

Selector_2 s670_5(wires_167_4[2], addr_167_4, wires_670_5,addr_670_5);

wire[3:0] wires_671_5;

wire[31:0] addr_671_5;

Selector_2 s671_5(wires_167_4[3], addr_167_4, wires_671_5,addr_671_5);

wire[3:0] wires_672_5;

wire[31:0] addr_672_5;

Selector_2 s672_5(wires_168_4[0], addr_168_4, wires_672_5,addr_672_5);

wire[3:0] wires_673_5;

wire[31:0] addr_673_5;

Selector_2 s673_5(wires_168_4[1], addr_168_4, wires_673_5,addr_673_5);

wire[3:0] wires_674_5;

wire[31:0] addr_674_5;

Selector_2 s674_5(wires_168_4[2], addr_168_4, wires_674_5,addr_674_5);

wire[3:0] wires_675_5;

wire[31:0] addr_675_5;

Selector_2 s675_5(wires_168_4[3], addr_168_4, wires_675_5,addr_675_5);

wire[3:0] wires_676_5;

wire[31:0] addr_676_5;

Selector_2 s676_5(wires_169_4[0], addr_169_4, wires_676_5,addr_676_5);

wire[3:0] wires_677_5;

wire[31:0] addr_677_5;

Selector_2 s677_5(wires_169_4[1], addr_169_4, wires_677_5,addr_677_5);

wire[3:0] wires_678_5;

wire[31:0] addr_678_5;

Selector_2 s678_5(wires_169_4[2], addr_169_4, wires_678_5,addr_678_5);

wire[3:0] wires_679_5;

wire[31:0] addr_679_5;

Selector_2 s679_5(wires_169_4[3], addr_169_4, wires_679_5,addr_679_5);

wire[3:0] wires_680_5;

wire[31:0] addr_680_5;

Selector_2 s680_5(wires_170_4[0], addr_170_4, wires_680_5,addr_680_5);

wire[3:0] wires_681_5;

wire[31:0] addr_681_5;

Selector_2 s681_5(wires_170_4[1], addr_170_4, wires_681_5,addr_681_5);

wire[3:0] wires_682_5;

wire[31:0] addr_682_5;

Selector_2 s682_5(wires_170_4[2], addr_170_4, wires_682_5,addr_682_5);

wire[3:0] wires_683_5;

wire[31:0] addr_683_5;

Selector_2 s683_5(wires_170_4[3], addr_170_4, wires_683_5,addr_683_5);

wire[3:0] wires_684_5;

wire[31:0] addr_684_5;

Selector_2 s684_5(wires_171_4[0], addr_171_4, wires_684_5,addr_684_5);

wire[3:0] wires_685_5;

wire[31:0] addr_685_5;

Selector_2 s685_5(wires_171_4[1], addr_171_4, wires_685_5,addr_685_5);

wire[3:0] wires_686_5;

wire[31:0] addr_686_5;

Selector_2 s686_5(wires_171_4[2], addr_171_4, wires_686_5,addr_686_5);

wire[3:0] wires_687_5;

wire[31:0] addr_687_5;

Selector_2 s687_5(wires_171_4[3], addr_171_4, wires_687_5,addr_687_5);

wire[3:0] wires_688_5;

wire[31:0] addr_688_5;

Selector_2 s688_5(wires_172_4[0], addr_172_4, wires_688_5,addr_688_5);

wire[3:0] wires_689_5;

wire[31:0] addr_689_5;

Selector_2 s689_5(wires_172_4[1], addr_172_4, wires_689_5,addr_689_5);

wire[3:0] wires_690_5;

wire[31:0] addr_690_5;

Selector_2 s690_5(wires_172_4[2], addr_172_4, wires_690_5,addr_690_5);

wire[3:0] wires_691_5;

wire[31:0] addr_691_5;

Selector_2 s691_5(wires_172_4[3], addr_172_4, wires_691_5,addr_691_5);

wire[3:0] wires_692_5;

wire[31:0] addr_692_5;

Selector_2 s692_5(wires_173_4[0], addr_173_4, wires_692_5,addr_692_5);

wire[3:0] wires_693_5;

wire[31:0] addr_693_5;

Selector_2 s693_5(wires_173_4[1], addr_173_4, wires_693_5,addr_693_5);

wire[3:0] wires_694_5;

wire[31:0] addr_694_5;

Selector_2 s694_5(wires_173_4[2], addr_173_4, wires_694_5,addr_694_5);

wire[3:0] wires_695_5;

wire[31:0] addr_695_5;

Selector_2 s695_5(wires_173_4[3], addr_173_4, wires_695_5,addr_695_5);

wire[3:0] wires_696_5;

wire[31:0] addr_696_5;

Selector_2 s696_5(wires_174_4[0], addr_174_4, wires_696_5,addr_696_5);

wire[3:0] wires_697_5;

wire[31:0] addr_697_5;

Selector_2 s697_5(wires_174_4[1], addr_174_4, wires_697_5,addr_697_5);

wire[3:0] wires_698_5;

wire[31:0] addr_698_5;

Selector_2 s698_5(wires_174_4[2], addr_174_4, wires_698_5,addr_698_5);

wire[3:0] wires_699_5;

wire[31:0] addr_699_5;

Selector_2 s699_5(wires_174_4[3], addr_174_4, wires_699_5,addr_699_5);

wire[3:0] wires_700_5;

wire[31:0] addr_700_5;

Selector_2 s700_5(wires_175_4[0], addr_175_4, wires_700_5,addr_700_5);

wire[3:0] wires_701_5;

wire[31:0] addr_701_5;

Selector_2 s701_5(wires_175_4[1], addr_175_4, wires_701_5,addr_701_5);

wire[3:0] wires_702_5;

wire[31:0] addr_702_5;

Selector_2 s702_5(wires_175_4[2], addr_175_4, wires_702_5,addr_702_5);

wire[3:0] wires_703_5;

wire[31:0] addr_703_5;

Selector_2 s703_5(wires_175_4[3], addr_175_4, wires_703_5,addr_703_5);

wire[3:0] wires_704_5;

wire[31:0] addr_704_5;

Selector_2 s704_5(wires_176_4[0], addr_176_4, wires_704_5,addr_704_5);

wire[3:0] wires_705_5;

wire[31:0] addr_705_5;

Selector_2 s705_5(wires_176_4[1], addr_176_4, wires_705_5,addr_705_5);

wire[3:0] wires_706_5;

wire[31:0] addr_706_5;

Selector_2 s706_5(wires_176_4[2], addr_176_4, wires_706_5,addr_706_5);

wire[3:0] wires_707_5;

wire[31:0] addr_707_5;

Selector_2 s707_5(wires_176_4[3], addr_176_4, wires_707_5,addr_707_5);

wire[3:0] wires_708_5;

wire[31:0] addr_708_5;

Selector_2 s708_5(wires_177_4[0], addr_177_4, wires_708_5,addr_708_5);

wire[3:0] wires_709_5;

wire[31:0] addr_709_5;

Selector_2 s709_5(wires_177_4[1], addr_177_4, wires_709_5,addr_709_5);

wire[3:0] wires_710_5;

wire[31:0] addr_710_5;

Selector_2 s710_5(wires_177_4[2], addr_177_4, wires_710_5,addr_710_5);

wire[3:0] wires_711_5;

wire[31:0] addr_711_5;

Selector_2 s711_5(wires_177_4[3], addr_177_4, wires_711_5,addr_711_5);

wire[3:0] wires_712_5;

wire[31:0] addr_712_5;

Selector_2 s712_5(wires_178_4[0], addr_178_4, wires_712_5,addr_712_5);

wire[3:0] wires_713_5;

wire[31:0] addr_713_5;

Selector_2 s713_5(wires_178_4[1], addr_178_4, wires_713_5,addr_713_5);

wire[3:0] wires_714_5;

wire[31:0] addr_714_5;

Selector_2 s714_5(wires_178_4[2], addr_178_4, wires_714_5,addr_714_5);

wire[3:0] wires_715_5;

wire[31:0] addr_715_5;

Selector_2 s715_5(wires_178_4[3], addr_178_4, wires_715_5,addr_715_5);

wire[3:0] wires_716_5;

wire[31:0] addr_716_5;

Selector_2 s716_5(wires_179_4[0], addr_179_4, wires_716_5,addr_716_5);

wire[3:0] wires_717_5;

wire[31:0] addr_717_5;

Selector_2 s717_5(wires_179_4[1], addr_179_4, wires_717_5,addr_717_5);

wire[3:0] wires_718_5;

wire[31:0] addr_718_5;

Selector_2 s718_5(wires_179_4[2], addr_179_4, wires_718_5,addr_718_5);

wire[3:0] wires_719_5;

wire[31:0] addr_719_5;

Selector_2 s719_5(wires_179_4[3], addr_179_4, wires_719_5,addr_719_5);

wire[3:0] wires_720_5;

wire[31:0] addr_720_5;

Selector_2 s720_5(wires_180_4[0], addr_180_4, wires_720_5,addr_720_5);

wire[3:0] wires_721_5;

wire[31:0] addr_721_5;

Selector_2 s721_5(wires_180_4[1], addr_180_4, wires_721_5,addr_721_5);

wire[3:0] wires_722_5;

wire[31:0] addr_722_5;

Selector_2 s722_5(wires_180_4[2], addr_180_4, wires_722_5,addr_722_5);

wire[3:0] wires_723_5;

wire[31:0] addr_723_5;

Selector_2 s723_5(wires_180_4[3], addr_180_4, wires_723_5,addr_723_5);

wire[3:0] wires_724_5;

wire[31:0] addr_724_5;

Selector_2 s724_5(wires_181_4[0], addr_181_4, wires_724_5,addr_724_5);

wire[3:0] wires_725_5;

wire[31:0] addr_725_5;

Selector_2 s725_5(wires_181_4[1], addr_181_4, wires_725_5,addr_725_5);

wire[3:0] wires_726_5;

wire[31:0] addr_726_5;

Selector_2 s726_5(wires_181_4[2], addr_181_4, wires_726_5,addr_726_5);

wire[3:0] wires_727_5;

wire[31:0] addr_727_5;

Selector_2 s727_5(wires_181_4[3], addr_181_4, wires_727_5,addr_727_5);

wire[3:0] wires_728_5;

wire[31:0] addr_728_5;

Selector_2 s728_5(wires_182_4[0], addr_182_4, wires_728_5,addr_728_5);

wire[3:0] wires_729_5;

wire[31:0] addr_729_5;

Selector_2 s729_5(wires_182_4[1], addr_182_4, wires_729_5,addr_729_5);

wire[3:0] wires_730_5;

wire[31:0] addr_730_5;

Selector_2 s730_5(wires_182_4[2], addr_182_4, wires_730_5,addr_730_5);

wire[3:0] wires_731_5;

wire[31:0] addr_731_5;

Selector_2 s731_5(wires_182_4[3], addr_182_4, wires_731_5,addr_731_5);

wire[3:0] wires_732_5;

wire[31:0] addr_732_5;

Selector_2 s732_5(wires_183_4[0], addr_183_4, wires_732_5,addr_732_5);

wire[3:0] wires_733_5;

wire[31:0] addr_733_5;

Selector_2 s733_5(wires_183_4[1], addr_183_4, wires_733_5,addr_733_5);

wire[3:0] wires_734_5;

wire[31:0] addr_734_5;

Selector_2 s734_5(wires_183_4[2], addr_183_4, wires_734_5,addr_734_5);

wire[3:0] wires_735_5;

wire[31:0] addr_735_5;

Selector_2 s735_5(wires_183_4[3], addr_183_4, wires_735_5,addr_735_5);

wire[3:0] wires_736_5;

wire[31:0] addr_736_5;

Selector_2 s736_5(wires_184_4[0], addr_184_4, wires_736_5,addr_736_5);

wire[3:0] wires_737_5;

wire[31:0] addr_737_5;

Selector_2 s737_5(wires_184_4[1], addr_184_4, wires_737_5,addr_737_5);

wire[3:0] wires_738_5;

wire[31:0] addr_738_5;

Selector_2 s738_5(wires_184_4[2], addr_184_4, wires_738_5,addr_738_5);

wire[3:0] wires_739_5;

wire[31:0] addr_739_5;

Selector_2 s739_5(wires_184_4[3], addr_184_4, wires_739_5,addr_739_5);

wire[3:0] wires_740_5;

wire[31:0] addr_740_5;

Selector_2 s740_5(wires_185_4[0], addr_185_4, wires_740_5,addr_740_5);

wire[3:0] wires_741_5;

wire[31:0] addr_741_5;

Selector_2 s741_5(wires_185_4[1], addr_185_4, wires_741_5,addr_741_5);

wire[3:0] wires_742_5;

wire[31:0] addr_742_5;

Selector_2 s742_5(wires_185_4[2], addr_185_4, wires_742_5,addr_742_5);

wire[3:0] wires_743_5;

wire[31:0] addr_743_5;

Selector_2 s743_5(wires_185_4[3], addr_185_4, wires_743_5,addr_743_5);

wire[3:0] wires_744_5;

wire[31:0] addr_744_5;

Selector_2 s744_5(wires_186_4[0], addr_186_4, wires_744_5,addr_744_5);

wire[3:0] wires_745_5;

wire[31:0] addr_745_5;

Selector_2 s745_5(wires_186_4[1], addr_186_4, wires_745_5,addr_745_5);

wire[3:0] wires_746_5;

wire[31:0] addr_746_5;

Selector_2 s746_5(wires_186_4[2], addr_186_4, wires_746_5,addr_746_5);

wire[3:0] wires_747_5;

wire[31:0] addr_747_5;

Selector_2 s747_5(wires_186_4[3], addr_186_4, wires_747_5,addr_747_5);

wire[3:0] wires_748_5;

wire[31:0] addr_748_5;

Selector_2 s748_5(wires_187_4[0], addr_187_4, wires_748_5,addr_748_5);

wire[3:0] wires_749_5;

wire[31:0] addr_749_5;

Selector_2 s749_5(wires_187_4[1], addr_187_4, wires_749_5,addr_749_5);

wire[3:0] wires_750_5;

wire[31:0] addr_750_5;

Selector_2 s750_5(wires_187_4[2], addr_187_4, wires_750_5,addr_750_5);

wire[3:0] wires_751_5;

wire[31:0] addr_751_5;

Selector_2 s751_5(wires_187_4[3], addr_187_4, wires_751_5,addr_751_5);

wire[3:0] wires_752_5;

wire[31:0] addr_752_5;

Selector_2 s752_5(wires_188_4[0], addr_188_4, wires_752_5,addr_752_5);

wire[3:0] wires_753_5;

wire[31:0] addr_753_5;

Selector_2 s753_5(wires_188_4[1], addr_188_4, wires_753_5,addr_753_5);

wire[3:0] wires_754_5;

wire[31:0] addr_754_5;

Selector_2 s754_5(wires_188_4[2], addr_188_4, wires_754_5,addr_754_5);

wire[3:0] wires_755_5;

wire[31:0] addr_755_5;

Selector_2 s755_5(wires_188_4[3], addr_188_4, wires_755_5,addr_755_5);

wire[3:0] wires_756_5;

wire[31:0] addr_756_5;

Selector_2 s756_5(wires_189_4[0], addr_189_4, wires_756_5,addr_756_5);

wire[3:0] wires_757_5;

wire[31:0] addr_757_5;

Selector_2 s757_5(wires_189_4[1], addr_189_4, wires_757_5,addr_757_5);

wire[3:0] wires_758_5;

wire[31:0] addr_758_5;

Selector_2 s758_5(wires_189_4[2], addr_189_4, wires_758_5,addr_758_5);

wire[3:0] wires_759_5;

wire[31:0] addr_759_5;

Selector_2 s759_5(wires_189_4[3], addr_189_4, wires_759_5,addr_759_5);

wire[3:0] wires_760_5;

wire[31:0] addr_760_5;

Selector_2 s760_5(wires_190_4[0], addr_190_4, wires_760_5,addr_760_5);

wire[3:0] wires_761_5;

wire[31:0] addr_761_5;

Selector_2 s761_5(wires_190_4[1], addr_190_4, wires_761_5,addr_761_5);

wire[3:0] wires_762_5;

wire[31:0] addr_762_5;

Selector_2 s762_5(wires_190_4[2], addr_190_4, wires_762_5,addr_762_5);

wire[3:0] wires_763_5;

wire[31:0] addr_763_5;

Selector_2 s763_5(wires_190_4[3], addr_190_4, wires_763_5,addr_763_5);

wire[3:0] wires_764_5;

wire[31:0] addr_764_5;

Selector_2 s764_5(wires_191_4[0], addr_191_4, wires_764_5,addr_764_5);

wire[3:0] wires_765_5;

wire[31:0] addr_765_5;

Selector_2 s765_5(wires_191_4[1], addr_191_4, wires_765_5,addr_765_5);

wire[3:0] wires_766_5;

wire[31:0] addr_766_5;

Selector_2 s766_5(wires_191_4[2], addr_191_4, wires_766_5,addr_766_5);

wire[3:0] wires_767_5;

wire[31:0] addr_767_5;

Selector_2 s767_5(wires_191_4[3], addr_191_4, wires_767_5,addr_767_5);

wire[3:0] wires_768_5;

wire[31:0] addr_768_5;

Selector_2 s768_5(wires_192_4[0], addr_192_4, wires_768_5,addr_768_5);

wire[3:0] wires_769_5;

wire[31:0] addr_769_5;

Selector_2 s769_5(wires_192_4[1], addr_192_4, wires_769_5,addr_769_5);

wire[3:0] wires_770_5;

wire[31:0] addr_770_5;

Selector_2 s770_5(wires_192_4[2], addr_192_4, wires_770_5,addr_770_5);

wire[3:0] wires_771_5;

wire[31:0] addr_771_5;

Selector_2 s771_5(wires_192_4[3], addr_192_4, wires_771_5,addr_771_5);

wire[3:0] wires_772_5;

wire[31:0] addr_772_5;

Selector_2 s772_5(wires_193_4[0], addr_193_4, wires_772_5,addr_772_5);

wire[3:0] wires_773_5;

wire[31:0] addr_773_5;

Selector_2 s773_5(wires_193_4[1], addr_193_4, wires_773_5,addr_773_5);

wire[3:0] wires_774_5;

wire[31:0] addr_774_5;

Selector_2 s774_5(wires_193_4[2], addr_193_4, wires_774_5,addr_774_5);

wire[3:0] wires_775_5;

wire[31:0] addr_775_5;

Selector_2 s775_5(wires_193_4[3], addr_193_4, wires_775_5,addr_775_5);

wire[3:0] wires_776_5;

wire[31:0] addr_776_5;

Selector_2 s776_5(wires_194_4[0], addr_194_4, wires_776_5,addr_776_5);

wire[3:0] wires_777_5;

wire[31:0] addr_777_5;

Selector_2 s777_5(wires_194_4[1], addr_194_4, wires_777_5,addr_777_5);

wire[3:0] wires_778_5;

wire[31:0] addr_778_5;

Selector_2 s778_5(wires_194_4[2], addr_194_4, wires_778_5,addr_778_5);

wire[3:0] wires_779_5;

wire[31:0] addr_779_5;

Selector_2 s779_5(wires_194_4[3], addr_194_4, wires_779_5,addr_779_5);

wire[3:0] wires_780_5;

wire[31:0] addr_780_5;

Selector_2 s780_5(wires_195_4[0], addr_195_4, wires_780_5,addr_780_5);

wire[3:0] wires_781_5;

wire[31:0] addr_781_5;

Selector_2 s781_5(wires_195_4[1], addr_195_4, wires_781_5,addr_781_5);

wire[3:0] wires_782_5;

wire[31:0] addr_782_5;

Selector_2 s782_5(wires_195_4[2], addr_195_4, wires_782_5,addr_782_5);

wire[3:0] wires_783_5;

wire[31:0] addr_783_5;

Selector_2 s783_5(wires_195_4[3], addr_195_4, wires_783_5,addr_783_5);

wire[3:0] wires_784_5;

wire[31:0] addr_784_5;

Selector_2 s784_5(wires_196_4[0], addr_196_4, wires_784_5,addr_784_5);

wire[3:0] wires_785_5;

wire[31:0] addr_785_5;

Selector_2 s785_5(wires_196_4[1], addr_196_4, wires_785_5,addr_785_5);

wire[3:0] wires_786_5;

wire[31:0] addr_786_5;

Selector_2 s786_5(wires_196_4[2], addr_196_4, wires_786_5,addr_786_5);

wire[3:0] wires_787_5;

wire[31:0] addr_787_5;

Selector_2 s787_5(wires_196_4[3], addr_196_4, wires_787_5,addr_787_5);

wire[3:0] wires_788_5;

wire[31:0] addr_788_5;

Selector_2 s788_5(wires_197_4[0], addr_197_4, wires_788_5,addr_788_5);

wire[3:0] wires_789_5;

wire[31:0] addr_789_5;

Selector_2 s789_5(wires_197_4[1], addr_197_4, wires_789_5,addr_789_5);

wire[3:0] wires_790_5;

wire[31:0] addr_790_5;

Selector_2 s790_5(wires_197_4[2], addr_197_4, wires_790_5,addr_790_5);

wire[3:0] wires_791_5;

wire[31:0] addr_791_5;

Selector_2 s791_5(wires_197_4[3], addr_197_4, wires_791_5,addr_791_5);

wire[3:0] wires_792_5;

wire[31:0] addr_792_5;

Selector_2 s792_5(wires_198_4[0], addr_198_4, wires_792_5,addr_792_5);

wire[3:0] wires_793_5;

wire[31:0] addr_793_5;

Selector_2 s793_5(wires_198_4[1], addr_198_4, wires_793_5,addr_793_5);

wire[3:0] wires_794_5;

wire[31:0] addr_794_5;

Selector_2 s794_5(wires_198_4[2], addr_198_4, wires_794_5,addr_794_5);

wire[3:0] wires_795_5;

wire[31:0] addr_795_5;

Selector_2 s795_5(wires_198_4[3], addr_198_4, wires_795_5,addr_795_5);

wire[3:0] wires_796_5;

wire[31:0] addr_796_5;

Selector_2 s796_5(wires_199_4[0], addr_199_4, wires_796_5,addr_796_5);

wire[3:0] wires_797_5;

wire[31:0] addr_797_5;

Selector_2 s797_5(wires_199_4[1], addr_199_4, wires_797_5,addr_797_5);

wire[3:0] wires_798_5;

wire[31:0] addr_798_5;

Selector_2 s798_5(wires_199_4[2], addr_199_4, wires_798_5,addr_798_5);

wire[3:0] wires_799_5;

wire[31:0] addr_799_5;

Selector_2 s799_5(wires_199_4[3], addr_199_4, wires_799_5,addr_799_5);

wire[3:0] wires_800_5;

wire[31:0] addr_800_5;

Selector_2 s800_5(wires_200_4[0], addr_200_4, wires_800_5,addr_800_5);

wire[3:0] wires_801_5;

wire[31:0] addr_801_5;

Selector_2 s801_5(wires_200_4[1], addr_200_4, wires_801_5,addr_801_5);

wire[3:0] wires_802_5;

wire[31:0] addr_802_5;

Selector_2 s802_5(wires_200_4[2], addr_200_4, wires_802_5,addr_802_5);

wire[3:0] wires_803_5;

wire[31:0] addr_803_5;

Selector_2 s803_5(wires_200_4[3], addr_200_4, wires_803_5,addr_803_5);

wire[3:0] wires_804_5;

wire[31:0] addr_804_5;

Selector_2 s804_5(wires_201_4[0], addr_201_4, wires_804_5,addr_804_5);

wire[3:0] wires_805_5;

wire[31:0] addr_805_5;

Selector_2 s805_5(wires_201_4[1], addr_201_4, wires_805_5,addr_805_5);

wire[3:0] wires_806_5;

wire[31:0] addr_806_5;

Selector_2 s806_5(wires_201_4[2], addr_201_4, wires_806_5,addr_806_5);

wire[3:0] wires_807_5;

wire[31:0] addr_807_5;

Selector_2 s807_5(wires_201_4[3], addr_201_4, wires_807_5,addr_807_5);

wire[3:0] wires_808_5;

wire[31:0] addr_808_5;

Selector_2 s808_5(wires_202_4[0], addr_202_4, wires_808_5,addr_808_5);

wire[3:0] wires_809_5;

wire[31:0] addr_809_5;

Selector_2 s809_5(wires_202_4[1], addr_202_4, wires_809_5,addr_809_5);

wire[3:0] wires_810_5;

wire[31:0] addr_810_5;

Selector_2 s810_5(wires_202_4[2], addr_202_4, wires_810_5,addr_810_5);

wire[3:0] wires_811_5;

wire[31:0] addr_811_5;

Selector_2 s811_5(wires_202_4[3], addr_202_4, wires_811_5,addr_811_5);

wire[3:0] wires_812_5;

wire[31:0] addr_812_5;

Selector_2 s812_5(wires_203_4[0], addr_203_4, wires_812_5,addr_812_5);

wire[3:0] wires_813_5;

wire[31:0] addr_813_5;

Selector_2 s813_5(wires_203_4[1], addr_203_4, wires_813_5,addr_813_5);

wire[3:0] wires_814_5;

wire[31:0] addr_814_5;

Selector_2 s814_5(wires_203_4[2], addr_203_4, wires_814_5,addr_814_5);

wire[3:0] wires_815_5;

wire[31:0] addr_815_5;

Selector_2 s815_5(wires_203_4[3], addr_203_4, wires_815_5,addr_815_5);

wire[3:0] wires_816_5;

wire[31:0] addr_816_5;

Selector_2 s816_5(wires_204_4[0], addr_204_4, wires_816_5,addr_816_5);

wire[3:0] wires_817_5;

wire[31:0] addr_817_5;

Selector_2 s817_5(wires_204_4[1], addr_204_4, wires_817_5,addr_817_5);

wire[3:0] wires_818_5;

wire[31:0] addr_818_5;

Selector_2 s818_5(wires_204_4[2], addr_204_4, wires_818_5,addr_818_5);

wire[3:0] wires_819_5;

wire[31:0] addr_819_5;

Selector_2 s819_5(wires_204_4[3], addr_204_4, wires_819_5,addr_819_5);

wire[3:0] wires_820_5;

wire[31:0] addr_820_5;

Selector_2 s820_5(wires_205_4[0], addr_205_4, wires_820_5,addr_820_5);

wire[3:0] wires_821_5;

wire[31:0] addr_821_5;

Selector_2 s821_5(wires_205_4[1], addr_205_4, wires_821_5,addr_821_5);

wire[3:0] wires_822_5;

wire[31:0] addr_822_5;

Selector_2 s822_5(wires_205_4[2], addr_205_4, wires_822_5,addr_822_5);

wire[3:0] wires_823_5;

wire[31:0] addr_823_5;

Selector_2 s823_5(wires_205_4[3], addr_205_4, wires_823_5,addr_823_5);

wire[3:0] wires_824_5;

wire[31:0] addr_824_5;

Selector_2 s824_5(wires_206_4[0], addr_206_4, wires_824_5,addr_824_5);

wire[3:0] wires_825_5;

wire[31:0] addr_825_5;

Selector_2 s825_5(wires_206_4[1], addr_206_4, wires_825_5,addr_825_5);

wire[3:0] wires_826_5;

wire[31:0] addr_826_5;

Selector_2 s826_5(wires_206_4[2], addr_206_4, wires_826_5,addr_826_5);

wire[3:0] wires_827_5;

wire[31:0] addr_827_5;

Selector_2 s827_5(wires_206_4[3], addr_206_4, wires_827_5,addr_827_5);

wire[3:0] wires_828_5;

wire[31:0] addr_828_5;

Selector_2 s828_5(wires_207_4[0], addr_207_4, wires_828_5,addr_828_5);

wire[3:0] wires_829_5;

wire[31:0] addr_829_5;

Selector_2 s829_5(wires_207_4[1], addr_207_4, wires_829_5,addr_829_5);

wire[3:0] wires_830_5;

wire[31:0] addr_830_5;

Selector_2 s830_5(wires_207_4[2], addr_207_4, wires_830_5,addr_830_5);

wire[3:0] wires_831_5;

wire[31:0] addr_831_5;

Selector_2 s831_5(wires_207_4[3], addr_207_4, wires_831_5,addr_831_5);

wire[3:0] wires_832_5;

wire[31:0] addr_832_5;

Selector_2 s832_5(wires_208_4[0], addr_208_4, wires_832_5,addr_832_5);

wire[3:0] wires_833_5;

wire[31:0] addr_833_5;

Selector_2 s833_5(wires_208_4[1], addr_208_4, wires_833_5,addr_833_5);

wire[3:0] wires_834_5;

wire[31:0] addr_834_5;

Selector_2 s834_5(wires_208_4[2], addr_208_4, wires_834_5,addr_834_5);

wire[3:0] wires_835_5;

wire[31:0] addr_835_5;

Selector_2 s835_5(wires_208_4[3], addr_208_4, wires_835_5,addr_835_5);

wire[3:0] wires_836_5;

wire[31:0] addr_836_5;

Selector_2 s836_5(wires_209_4[0], addr_209_4, wires_836_5,addr_836_5);

wire[3:0] wires_837_5;

wire[31:0] addr_837_5;

Selector_2 s837_5(wires_209_4[1], addr_209_4, wires_837_5,addr_837_5);

wire[3:0] wires_838_5;

wire[31:0] addr_838_5;

Selector_2 s838_5(wires_209_4[2], addr_209_4, wires_838_5,addr_838_5);

wire[3:0] wires_839_5;

wire[31:0] addr_839_5;

Selector_2 s839_5(wires_209_4[3], addr_209_4, wires_839_5,addr_839_5);

wire[3:0] wires_840_5;

wire[31:0] addr_840_5;

Selector_2 s840_5(wires_210_4[0], addr_210_4, wires_840_5,addr_840_5);

wire[3:0] wires_841_5;

wire[31:0] addr_841_5;

Selector_2 s841_5(wires_210_4[1], addr_210_4, wires_841_5,addr_841_5);

wire[3:0] wires_842_5;

wire[31:0] addr_842_5;

Selector_2 s842_5(wires_210_4[2], addr_210_4, wires_842_5,addr_842_5);

wire[3:0] wires_843_5;

wire[31:0] addr_843_5;

Selector_2 s843_5(wires_210_4[3], addr_210_4, wires_843_5,addr_843_5);

wire[3:0] wires_844_5;

wire[31:0] addr_844_5;

Selector_2 s844_5(wires_211_4[0], addr_211_4, wires_844_5,addr_844_5);

wire[3:0] wires_845_5;

wire[31:0] addr_845_5;

Selector_2 s845_5(wires_211_4[1], addr_211_4, wires_845_5,addr_845_5);

wire[3:0] wires_846_5;

wire[31:0] addr_846_5;

Selector_2 s846_5(wires_211_4[2], addr_211_4, wires_846_5,addr_846_5);

wire[3:0] wires_847_5;

wire[31:0] addr_847_5;

Selector_2 s847_5(wires_211_4[3], addr_211_4, wires_847_5,addr_847_5);

wire[3:0] wires_848_5;

wire[31:0] addr_848_5;

Selector_2 s848_5(wires_212_4[0], addr_212_4, wires_848_5,addr_848_5);

wire[3:0] wires_849_5;

wire[31:0] addr_849_5;

Selector_2 s849_5(wires_212_4[1], addr_212_4, wires_849_5,addr_849_5);

wire[3:0] wires_850_5;

wire[31:0] addr_850_5;

Selector_2 s850_5(wires_212_4[2], addr_212_4, wires_850_5,addr_850_5);

wire[3:0] wires_851_5;

wire[31:0] addr_851_5;

Selector_2 s851_5(wires_212_4[3], addr_212_4, wires_851_5,addr_851_5);

wire[3:0] wires_852_5;

wire[31:0] addr_852_5;

Selector_2 s852_5(wires_213_4[0], addr_213_4, wires_852_5,addr_852_5);

wire[3:0] wires_853_5;

wire[31:0] addr_853_5;

Selector_2 s853_5(wires_213_4[1], addr_213_4, wires_853_5,addr_853_5);

wire[3:0] wires_854_5;

wire[31:0] addr_854_5;

Selector_2 s854_5(wires_213_4[2], addr_213_4, wires_854_5,addr_854_5);

wire[3:0] wires_855_5;

wire[31:0] addr_855_5;

Selector_2 s855_5(wires_213_4[3], addr_213_4, wires_855_5,addr_855_5);

wire[3:0] wires_856_5;

wire[31:0] addr_856_5;

Selector_2 s856_5(wires_214_4[0], addr_214_4, wires_856_5,addr_856_5);

wire[3:0] wires_857_5;

wire[31:0] addr_857_5;

Selector_2 s857_5(wires_214_4[1], addr_214_4, wires_857_5,addr_857_5);

wire[3:0] wires_858_5;

wire[31:0] addr_858_5;

Selector_2 s858_5(wires_214_4[2], addr_214_4, wires_858_5,addr_858_5);

wire[3:0] wires_859_5;

wire[31:0] addr_859_5;

Selector_2 s859_5(wires_214_4[3], addr_214_4, wires_859_5,addr_859_5);

wire[3:0] wires_860_5;

wire[31:0] addr_860_5;

Selector_2 s860_5(wires_215_4[0], addr_215_4, wires_860_5,addr_860_5);

wire[3:0] wires_861_5;

wire[31:0] addr_861_5;

Selector_2 s861_5(wires_215_4[1], addr_215_4, wires_861_5,addr_861_5);

wire[3:0] wires_862_5;

wire[31:0] addr_862_5;

Selector_2 s862_5(wires_215_4[2], addr_215_4, wires_862_5,addr_862_5);

wire[3:0] wires_863_5;

wire[31:0] addr_863_5;

Selector_2 s863_5(wires_215_4[3], addr_215_4, wires_863_5,addr_863_5);

wire[3:0] wires_864_5;

wire[31:0] addr_864_5;

Selector_2 s864_5(wires_216_4[0], addr_216_4, wires_864_5,addr_864_5);

wire[3:0] wires_865_5;

wire[31:0] addr_865_5;

Selector_2 s865_5(wires_216_4[1], addr_216_4, wires_865_5,addr_865_5);

wire[3:0] wires_866_5;

wire[31:0] addr_866_5;

Selector_2 s866_5(wires_216_4[2], addr_216_4, wires_866_5,addr_866_5);

wire[3:0] wires_867_5;

wire[31:0] addr_867_5;

Selector_2 s867_5(wires_216_4[3], addr_216_4, wires_867_5,addr_867_5);

wire[3:0] wires_868_5;

wire[31:0] addr_868_5;

Selector_2 s868_5(wires_217_4[0], addr_217_4, wires_868_5,addr_868_5);

wire[3:0] wires_869_5;

wire[31:0] addr_869_5;

Selector_2 s869_5(wires_217_4[1], addr_217_4, wires_869_5,addr_869_5);

wire[3:0] wires_870_5;

wire[31:0] addr_870_5;

Selector_2 s870_5(wires_217_4[2], addr_217_4, wires_870_5,addr_870_5);

wire[3:0] wires_871_5;

wire[31:0] addr_871_5;

Selector_2 s871_5(wires_217_4[3], addr_217_4, wires_871_5,addr_871_5);

wire[3:0] wires_872_5;

wire[31:0] addr_872_5;

Selector_2 s872_5(wires_218_4[0], addr_218_4, wires_872_5,addr_872_5);

wire[3:0] wires_873_5;

wire[31:0] addr_873_5;

Selector_2 s873_5(wires_218_4[1], addr_218_4, wires_873_5,addr_873_5);

wire[3:0] wires_874_5;

wire[31:0] addr_874_5;

Selector_2 s874_5(wires_218_4[2], addr_218_4, wires_874_5,addr_874_5);

wire[3:0] wires_875_5;

wire[31:0] addr_875_5;

Selector_2 s875_5(wires_218_4[3], addr_218_4, wires_875_5,addr_875_5);

wire[3:0] wires_876_5;

wire[31:0] addr_876_5;

Selector_2 s876_5(wires_219_4[0], addr_219_4, wires_876_5,addr_876_5);

wire[3:0] wires_877_5;

wire[31:0] addr_877_5;

Selector_2 s877_5(wires_219_4[1], addr_219_4, wires_877_5,addr_877_5);

wire[3:0] wires_878_5;

wire[31:0] addr_878_5;

Selector_2 s878_5(wires_219_4[2], addr_219_4, wires_878_5,addr_878_5);

wire[3:0] wires_879_5;

wire[31:0] addr_879_5;

Selector_2 s879_5(wires_219_4[3], addr_219_4, wires_879_5,addr_879_5);

wire[3:0] wires_880_5;

wire[31:0] addr_880_5;

Selector_2 s880_5(wires_220_4[0], addr_220_4, wires_880_5,addr_880_5);

wire[3:0] wires_881_5;

wire[31:0] addr_881_5;

Selector_2 s881_5(wires_220_4[1], addr_220_4, wires_881_5,addr_881_5);

wire[3:0] wires_882_5;

wire[31:0] addr_882_5;

Selector_2 s882_5(wires_220_4[2], addr_220_4, wires_882_5,addr_882_5);

wire[3:0] wires_883_5;

wire[31:0] addr_883_5;

Selector_2 s883_5(wires_220_4[3], addr_220_4, wires_883_5,addr_883_5);

wire[3:0] wires_884_5;

wire[31:0] addr_884_5;

Selector_2 s884_5(wires_221_4[0], addr_221_4, wires_884_5,addr_884_5);

wire[3:0] wires_885_5;

wire[31:0] addr_885_5;

Selector_2 s885_5(wires_221_4[1], addr_221_4, wires_885_5,addr_885_5);

wire[3:0] wires_886_5;

wire[31:0] addr_886_5;

Selector_2 s886_5(wires_221_4[2], addr_221_4, wires_886_5,addr_886_5);

wire[3:0] wires_887_5;

wire[31:0] addr_887_5;

Selector_2 s887_5(wires_221_4[3], addr_221_4, wires_887_5,addr_887_5);

wire[3:0] wires_888_5;

wire[31:0] addr_888_5;

Selector_2 s888_5(wires_222_4[0], addr_222_4, wires_888_5,addr_888_5);

wire[3:0] wires_889_5;

wire[31:0] addr_889_5;

Selector_2 s889_5(wires_222_4[1], addr_222_4, wires_889_5,addr_889_5);

wire[3:0] wires_890_5;

wire[31:0] addr_890_5;

Selector_2 s890_5(wires_222_4[2], addr_222_4, wires_890_5,addr_890_5);

wire[3:0] wires_891_5;

wire[31:0] addr_891_5;

Selector_2 s891_5(wires_222_4[3], addr_222_4, wires_891_5,addr_891_5);

wire[3:0] wires_892_5;

wire[31:0] addr_892_5;

Selector_2 s892_5(wires_223_4[0], addr_223_4, wires_892_5,addr_892_5);

wire[3:0] wires_893_5;

wire[31:0] addr_893_5;

Selector_2 s893_5(wires_223_4[1], addr_223_4, wires_893_5,addr_893_5);

wire[3:0] wires_894_5;

wire[31:0] addr_894_5;

Selector_2 s894_5(wires_223_4[2], addr_223_4, wires_894_5,addr_894_5);

wire[3:0] wires_895_5;

wire[31:0] addr_895_5;

Selector_2 s895_5(wires_223_4[3], addr_223_4, wires_895_5,addr_895_5);

wire[3:0] wires_896_5;

wire[31:0] addr_896_5;

Selector_2 s896_5(wires_224_4[0], addr_224_4, wires_896_5,addr_896_5);

wire[3:0] wires_897_5;

wire[31:0] addr_897_5;

Selector_2 s897_5(wires_224_4[1], addr_224_4, wires_897_5,addr_897_5);

wire[3:0] wires_898_5;

wire[31:0] addr_898_5;

Selector_2 s898_5(wires_224_4[2], addr_224_4, wires_898_5,addr_898_5);

wire[3:0] wires_899_5;

wire[31:0] addr_899_5;

Selector_2 s899_5(wires_224_4[3], addr_224_4, wires_899_5,addr_899_5);

wire[3:0] wires_900_5;

wire[31:0] addr_900_5;

Selector_2 s900_5(wires_225_4[0], addr_225_4, wires_900_5,addr_900_5);

wire[3:0] wires_901_5;

wire[31:0] addr_901_5;

Selector_2 s901_5(wires_225_4[1], addr_225_4, wires_901_5,addr_901_5);

wire[3:0] wires_902_5;

wire[31:0] addr_902_5;

Selector_2 s902_5(wires_225_4[2], addr_225_4, wires_902_5,addr_902_5);

wire[3:0] wires_903_5;

wire[31:0] addr_903_5;

Selector_2 s903_5(wires_225_4[3], addr_225_4, wires_903_5,addr_903_5);

wire[3:0] wires_904_5;

wire[31:0] addr_904_5;

Selector_2 s904_5(wires_226_4[0], addr_226_4, wires_904_5,addr_904_5);

wire[3:0] wires_905_5;

wire[31:0] addr_905_5;

Selector_2 s905_5(wires_226_4[1], addr_226_4, wires_905_5,addr_905_5);

wire[3:0] wires_906_5;

wire[31:0] addr_906_5;

Selector_2 s906_5(wires_226_4[2], addr_226_4, wires_906_5,addr_906_5);

wire[3:0] wires_907_5;

wire[31:0] addr_907_5;

Selector_2 s907_5(wires_226_4[3], addr_226_4, wires_907_5,addr_907_5);

wire[3:0] wires_908_5;

wire[31:0] addr_908_5;

Selector_2 s908_5(wires_227_4[0], addr_227_4, wires_908_5,addr_908_5);

wire[3:0] wires_909_5;

wire[31:0] addr_909_5;

Selector_2 s909_5(wires_227_4[1], addr_227_4, wires_909_5,addr_909_5);

wire[3:0] wires_910_5;

wire[31:0] addr_910_5;

Selector_2 s910_5(wires_227_4[2], addr_227_4, wires_910_5,addr_910_5);

wire[3:0] wires_911_5;

wire[31:0] addr_911_5;

Selector_2 s911_5(wires_227_4[3], addr_227_4, wires_911_5,addr_911_5);

wire[3:0] wires_912_5;

wire[31:0] addr_912_5;

Selector_2 s912_5(wires_228_4[0], addr_228_4, wires_912_5,addr_912_5);

wire[3:0] wires_913_5;

wire[31:0] addr_913_5;

Selector_2 s913_5(wires_228_4[1], addr_228_4, wires_913_5,addr_913_5);

wire[3:0] wires_914_5;

wire[31:0] addr_914_5;

Selector_2 s914_5(wires_228_4[2], addr_228_4, wires_914_5,addr_914_5);

wire[3:0] wires_915_5;

wire[31:0] addr_915_5;

Selector_2 s915_5(wires_228_4[3], addr_228_4, wires_915_5,addr_915_5);

wire[3:0] wires_916_5;

wire[31:0] addr_916_5;

Selector_2 s916_5(wires_229_4[0], addr_229_4, wires_916_5,addr_916_5);

wire[3:0] wires_917_5;

wire[31:0] addr_917_5;

Selector_2 s917_5(wires_229_4[1], addr_229_4, wires_917_5,addr_917_5);

wire[3:0] wires_918_5;

wire[31:0] addr_918_5;

Selector_2 s918_5(wires_229_4[2], addr_229_4, wires_918_5,addr_918_5);

wire[3:0] wires_919_5;

wire[31:0] addr_919_5;

Selector_2 s919_5(wires_229_4[3], addr_229_4, wires_919_5,addr_919_5);

wire[3:0] wires_920_5;

wire[31:0] addr_920_5;

Selector_2 s920_5(wires_230_4[0], addr_230_4, wires_920_5,addr_920_5);

wire[3:0] wires_921_5;

wire[31:0] addr_921_5;

Selector_2 s921_5(wires_230_4[1], addr_230_4, wires_921_5,addr_921_5);

wire[3:0] wires_922_5;

wire[31:0] addr_922_5;

Selector_2 s922_5(wires_230_4[2], addr_230_4, wires_922_5,addr_922_5);

wire[3:0] wires_923_5;

wire[31:0] addr_923_5;

Selector_2 s923_5(wires_230_4[3], addr_230_4, wires_923_5,addr_923_5);

wire[3:0] wires_924_5;

wire[31:0] addr_924_5;

Selector_2 s924_5(wires_231_4[0], addr_231_4, wires_924_5,addr_924_5);

wire[3:0] wires_925_5;

wire[31:0] addr_925_5;

Selector_2 s925_5(wires_231_4[1], addr_231_4, wires_925_5,addr_925_5);

wire[3:0] wires_926_5;

wire[31:0] addr_926_5;

Selector_2 s926_5(wires_231_4[2], addr_231_4, wires_926_5,addr_926_5);

wire[3:0] wires_927_5;

wire[31:0] addr_927_5;

Selector_2 s927_5(wires_231_4[3], addr_231_4, wires_927_5,addr_927_5);

wire[3:0] wires_928_5;

wire[31:0] addr_928_5;

Selector_2 s928_5(wires_232_4[0], addr_232_4, wires_928_5,addr_928_5);

wire[3:0] wires_929_5;

wire[31:0] addr_929_5;

Selector_2 s929_5(wires_232_4[1], addr_232_4, wires_929_5,addr_929_5);

wire[3:0] wires_930_5;

wire[31:0] addr_930_5;

Selector_2 s930_5(wires_232_4[2], addr_232_4, wires_930_5,addr_930_5);

wire[3:0] wires_931_5;

wire[31:0] addr_931_5;

Selector_2 s931_5(wires_232_4[3], addr_232_4, wires_931_5,addr_931_5);

wire[3:0] wires_932_5;

wire[31:0] addr_932_5;

Selector_2 s932_5(wires_233_4[0], addr_233_4, wires_932_5,addr_932_5);

wire[3:0] wires_933_5;

wire[31:0] addr_933_5;

Selector_2 s933_5(wires_233_4[1], addr_233_4, wires_933_5,addr_933_5);

wire[3:0] wires_934_5;

wire[31:0] addr_934_5;

Selector_2 s934_5(wires_233_4[2], addr_233_4, wires_934_5,addr_934_5);

wire[3:0] wires_935_5;

wire[31:0] addr_935_5;

Selector_2 s935_5(wires_233_4[3], addr_233_4, wires_935_5,addr_935_5);

wire[3:0] wires_936_5;

wire[31:0] addr_936_5;

Selector_2 s936_5(wires_234_4[0], addr_234_4, wires_936_5,addr_936_5);

wire[3:0] wires_937_5;

wire[31:0] addr_937_5;

Selector_2 s937_5(wires_234_4[1], addr_234_4, wires_937_5,addr_937_5);

wire[3:0] wires_938_5;

wire[31:0] addr_938_5;

Selector_2 s938_5(wires_234_4[2], addr_234_4, wires_938_5,addr_938_5);

wire[3:0] wires_939_5;

wire[31:0] addr_939_5;

Selector_2 s939_5(wires_234_4[3], addr_234_4, wires_939_5,addr_939_5);

wire[3:0] wires_940_5;

wire[31:0] addr_940_5;

Selector_2 s940_5(wires_235_4[0], addr_235_4, wires_940_5,addr_940_5);

wire[3:0] wires_941_5;

wire[31:0] addr_941_5;

Selector_2 s941_5(wires_235_4[1], addr_235_4, wires_941_5,addr_941_5);

wire[3:0] wires_942_5;

wire[31:0] addr_942_5;

Selector_2 s942_5(wires_235_4[2], addr_235_4, wires_942_5,addr_942_5);

wire[3:0] wires_943_5;

wire[31:0] addr_943_5;

Selector_2 s943_5(wires_235_4[3], addr_235_4, wires_943_5,addr_943_5);

wire[3:0] wires_944_5;

wire[31:0] addr_944_5;

Selector_2 s944_5(wires_236_4[0], addr_236_4, wires_944_5,addr_944_5);

wire[3:0] wires_945_5;

wire[31:0] addr_945_5;

Selector_2 s945_5(wires_236_4[1], addr_236_4, wires_945_5,addr_945_5);

wire[3:0] wires_946_5;

wire[31:0] addr_946_5;

Selector_2 s946_5(wires_236_4[2], addr_236_4, wires_946_5,addr_946_5);

wire[3:0] wires_947_5;

wire[31:0] addr_947_5;

Selector_2 s947_5(wires_236_4[3], addr_236_4, wires_947_5,addr_947_5);

wire[3:0] wires_948_5;

wire[31:0] addr_948_5;

Selector_2 s948_5(wires_237_4[0], addr_237_4, wires_948_5,addr_948_5);

wire[3:0] wires_949_5;

wire[31:0] addr_949_5;

Selector_2 s949_5(wires_237_4[1], addr_237_4, wires_949_5,addr_949_5);

wire[3:0] wires_950_5;

wire[31:0] addr_950_5;

Selector_2 s950_5(wires_237_4[2], addr_237_4, wires_950_5,addr_950_5);

wire[3:0] wires_951_5;

wire[31:0] addr_951_5;

Selector_2 s951_5(wires_237_4[3], addr_237_4, wires_951_5,addr_951_5);

wire[3:0] wires_952_5;

wire[31:0] addr_952_5;

Selector_2 s952_5(wires_238_4[0], addr_238_4, wires_952_5,addr_952_5);

wire[3:0] wires_953_5;

wire[31:0] addr_953_5;

Selector_2 s953_5(wires_238_4[1], addr_238_4, wires_953_5,addr_953_5);

wire[3:0] wires_954_5;

wire[31:0] addr_954_5;

Selector_2 s954_5(wires_238_4[2], addr_238_4, wires_954_5,addr_954_5);

wire[3:0] wires_955_5;

wire[31:0] addr_955_5;

Selector_2 s955_5(wires_238_4[3], addr_238_4, wires_955_5,addr_955_5);

wire[3:0] wires_956_5;

wire[31:0] addr_956_5;

Selector_2 s956_5(wires_239_4[0], addr_239_4, wires_956_5,addr_956_5);

wire[3:0] wires_957_5;

wire[31:0] addr_957_5;

Selector_2 s957_5(wires_239_4[1], addr_239_4, wires_957_5,addr_957_5);

wire[3:0] wires_958_5;

wire[31:0] addr_958_5;

Selector_2 s958_5(wires_239_4[2], addr_239_4, wires_958_5,addr_958_5);

wire[3:0] wires_959_5;

wire[31:0] addr_959_5;

Selector_2 s959_5(wires_239_4[3], addr_239_4, wires_959_5,addr_959_5);

wire[3:0] wires_960_5;

wire[31:0] addr_960_5;

Selector_2 s960_5(wires_240_4[0], addr_240_4, wires_960_5,addr_960_5);

wire[3:0] wires_961_5;

wire[31:0] addr_961_5;

Selector_2 s961_5(wires_240_4[1], addr_240_4, wires_961_5,addr_961_5);

wire[3:0] wires_962_5;

wire[31:0] addr_962_5;

Selector_2 s962_5(wires_240_4[2], addr_240_4, wires_962_5,addr_962_5);

wire[3:0] wires_963_5;

wire[31:0] addr_963_5;

Selector_2 s963_5(wires_240_4[3], addr_240_4, wires_963_5,addr_963_5);

wire[3:0] wires_964_5;

wire[31:0] addr_964_5;

Selector_2 s964_5(wires_241_4[0], addr_241_4, wires_964_5,addr_964_5);

wire[3:0] wires_965_5;

wire[31:0] addr_965_5;

Selector_2 s965_5(wires_241_4[1], addr_241_4, wires_965_5,addr_965_5);

wire[3:0] wires_966_5;

wire[31:0] addr_966_5;

Selector_2 s966_5(wires_241_4[2], addr_241_4, wires_966_5,addr_966_5);

wire[3:0] wires_967_5;

wire[31:0] addr_967_5;

Selector_2 s967_5(wires_241_4[3], addr_241_4, wires_967_5,addr_967_5);

wire[3:0] wires_968_5;

wire[31:0] addr_968_5;

Selector_2 s968_5(wires_242_4[0], addr_242_4, wires_968_5,addr_968_5);

wire[3:0] wires_969_5;

wire[31:0] addr_969_5;

Selector_2 s969_5(wires_242_4[1], addr_242_4, wires_969_5,addr_969_5);

wire[3:0] wires_970_5;

wire[31:0] addr_970_5;

Selector_2 s970_5(wires_242_4[2], addr_242_4, wires_970_5,addr_970_5);

wire[3:0] wires_971_5;

wire[31:0] addr_971_5;

Selector_2 s971_5(wires_242_4[3], addr_242_4, wires_971_5,addr_971_5);

wire[3:0] wires_972_5;

wire[31:0] addr_972_5;

Selector_2 s972_5(wires_243_4[0], addr_243_4, wires_972_5,addr_972_5);

wire[3:0] wires_973_5;

wire[31:0] addr_973_5;

Selector_2 s973_5(wires_243_4[1], addr_243_4, wires_973_5,addr_973_5);

wire[3:0] wires_974_5;

wire[31:0] addr_974_5;

Selector_2 s974_5(wires_243_4[2], addr_243_4, wires_974_5,addr_974_5);

wire[3:0] wires_975_5;

wire[31:0] addr_975_5;

Selector_2 s975_5(wires_243_4[3], addr_243_4, wires_975_5,addr_975_5);

wire[3:0] wires_976_5;

wire[31:0] addr_976_5;

Selector_2 s976_5(wires_244_4[0], addr_244_4, wires_976_5,addr_976_5);

wire[3:0] wires_977_5;

wire[31:0] addr_977_5;

Selector_2 s977_5(wires_244_4[1], addr_244_4, wires_977_5,addr_977_5);

wire[3:0] wires_978_5;

wire[31:0] addr_978_5;

Selector_2 s978_5(wires_244_4[2], addr_244_4, wires_978_5,addr_978_5);

wire[3:0] wires_979_5;

wire[31:0] addr_979_5;

Selector_2 s979_5(wires_244_4[3], addr_244_4, wires_979_5,addr_979_5);

wire[3:0] wires_980_5;

wire[31:0] addr_980_5;

Selector_2 s980_5(wires_245_4[0], addr_245_4, wires_980_5,addr_980_5);

wire[3:0] wires_981_5;

wire[31:0] addr_981_5;

Selector_2 s981_5(wires_245_4[1], addr_245_4, wires_981_5,addr_981_5);

wire[3:0] wires_982_5;

wire[31:0] addr_982_5;

Selector_2 s982_5(wires_245_4[2], addr_245_4, wires_982_5,addr_982_5);

wire[3:0] wires_983_5;

wire[31:0] addr_983_5;

Selector_2 s983_5(wires_245_4[3], addr_245_4, wires_983_5,addr_983_5);

wire[3:0] wires_984_5;

wire[31:0] addr_984_5;

Selector_2 s984_5(wires_246_4[0], addr_246_4, wires_984_5,addr_984_5);

wire[3:0] wires_985_5;

wire[31:0] addr_985_5;

Selector_2 s985_5(wires_246_4[1], addr_246_4, wires_985_5,addr_985_5);

wire[3:0] wires_986_5;

wire[31:0] addr_986_5;

Selector_2 s986_5(wires_246_4[2], addr_246_4, wires_986_5,addr_986_5);

wire[3:0] wires_987_5;

wire[31:0] addr_987_5;

Selector_2 s987_5(wires_246_4[3], addr_246_4, wires_987_5,addr_987_5);

wire[3:0] wires_988_5;

wire[31:0] addr_988_5;

Selector_2 s988_5(wires_247_4[0], addr_247_4, wires_988_5,addr_988_5);

wire[3:0] wires_989_5;

wire[31:0] addr_989_5;

Selector_2 s989_5(wires_247_4[1], addr_247_4, wires_989_5,addr_989_5);

wire[3:0] wires_990_5;

wire[31:0] addr_990_5;

Selector_2 s990_5(wires_247_4[2], addr_247_4, wires_990_5,addr_990_5);

wire[3:0] wires_991_5;

wire[31:0] addr_991_5;

Selector_2 s991_5(wires_247_4[3], addr_247_4, wires_991_5,addr_991_5);

wire[3:0] wires_992_5;

wire[31:0] addr_992_5;

Selector_2 s992_5(wires_248_4[0], addr_248_4, wires_992_5,addr_992_5);

wire[3:0] wires_993_5;

wire[31:0] addr_993_5;

Selector_2 s993_5(wires_248_4[1], addr_248_4, wires_993_5,addr_993_5);

wire[3:0] wires_994_5;

wire[31:0] addr_994_5;

Selector_2 s994_5(wires_248_4[2], addr_248_4, wires_994_5,addr_994_5);

wire[3:0] wires_995_5;

wire[31:0] addr_995_5;

Selector_2 s995_5(wires_248_4[3], addr_248_4, wires_995_5,addr_995_5);

wire[3:0] wires_996_5;

wire[31:0] addr_996_5;

Selector_2 s996_5(wires_249_4[0], addr_249_4, wires_996_5,addr_996_5);

wire[3:0] wires_997_5;

wire[31:0] addr_997_5;

Selector_2 s997_5(wires_249_4[1], addr_249_4, wires_997_5,addr_997_5);

wire[3:0] wires_998_5;

wire[31:0] addr_998_5;

Selector_2 s998_5(wires_249_4[2], addr_249_4, wires_998_5,addr_998_5);

wire[3:0] wires_999_5;

wire[31:0] addr_999_5;

Selector_2 s999_5(wires_249_4[3], addr_249_4, wires_999_5,addr_999_5);

wire[3:0] wires_1000_5;

wire[31:0] addr_1000_5;

Selector_2 s1000_5(wires_250_4[0], addr_250_4, wires_1000_5,addr_1000_5);

wire[3:0] wires_1001_5;

wire[31:0] addr_1001_5;

Selector_2 s1001_5(wires_250_4[1], addr_250_4, wires_1001_5,addr_1001_5);

wire[3:0] wires_1002_5;

wire[31:0] addr_1002_5;

Selector_2 s1002_5(wires_250_4[2], addr_250_4, wires_1002_5,addr_1002_5);

wire[3:0] wires_1003_5;

wire[31:0] addr_1003_5;

Selector_2 s1003_5(wires_250_4[3], addr_250_4, wires_1003_5,addr_1003_5);

wire[3:0] wires_1004_5;

wire[31:0] addr_1004_5;

Selector_2 s1004_5(wires_251_4[0], addr_251_4, wires_1004_5,addr_1004_5);

wire[3:0] wires_1005_5;

wire[31:0] addr_1005_5;

Selector_2 s1005_5(wires_251_4[1], addr_251_4, wires_1005_5,addr_1005_5);

wire[3:0] wires_1006_5;

wire[31:0] addr_1006_5;

Selector_2 s1006_5(wires_251_4[2], addr_251_4, wires_1006_5,addr_1006_5);

wire[3:0] wires_1007_5;

wire[31:0] addr_1007_5;

Selector_2 s1007_5(wires_251_4[3], addr_251_4, wires_1007_5,addr_1007_5);

wire[3:0] wires_1008_5;

wire[31:0] addr_1008_5;

Selector_2 s1008_5(wires_252_4[0], addr_252_4, wires_1008_5,addr_1008_5);

wire[3:0] wires_1009_5;

wire[31:0] addr_1009_5;

Selector_2 s1009_5(wires_252_4[1], addr_252_4, wires_1009_5,addr_1009_5);

wire[3:0] wires_1010_5;

wire[31:0] addr_1010_5;

Selector_2 s1010_5(wires_252_4[2], addr_252_4, wires_1010_5,addr_1010_5);

wire[3:0] wires_1011_5;

wire[31:0] addr_1011_5;

Selector_2 s1011_5(wires_252_4[3], addr_252_4, wires_1011_5,addr_1011_5);

wire[3:0] wires_1012_5;

wire[31:0] addr_1012_5;

Selector_2 s1012_5(wires_253_4[0], addr_253_4, wires_1012_5,addr_1012_5);

wire[3:0] wires_1013_5;

wire[31:0] addr_1013_5;

Selector_2 s1013_5(wires_253_4[1], addr_253_4, wires_1013_5,addr_1013_5);

wire[3:0] wires_1014_5;

wire[31:0] addr_1014_5;

Selector_2 s1014_5(wires_253_4[2], addr_253_4, wires_1014_5,addr_1014_5);

wire[3:0] wires_1015_5;

wire[31:0] addr_1015_5;

Selector_2 s1015_5(wires_253_4[3], addr_253_4, wires_1015_5,addr_1015_5);

wire[3:0] wires_1016_5;

wire[31:0] addr_1016_5;

Selector_2 s1016_5(wires_254_4[0], addr_254_4, wires_1016_5,addr_1016_5);

wire[3:0] wires_1017_5;

wire[31:0] addr_1017_5;

Selector_2 s1017_5(wires_254_4[1], addr_254_4, wires_1017_5,addr_1017_5);

wire[3:0] wires_1018_5;

wire[31:0] addr_1018_5;

Selector_2 s1018_5(wires_254_4[2], addr_254_4, wires_1018_5,addr_1018_5);

wire[3:0] wires_1019_5;

wire[31:0] addr_1019_5;

Selector_2 s1019_5(wires_254_4[3], addr_254_4, wires_1019_5,addr_1019_5);

wire[3:0] wires_1020_5;

wire[31:0] addr_1020_5;

Selector_2 s1020_5(wires_255_4[0], addr_255_4, wires_1020_5,addr_1020_5);

wire[3:0] wires_1021_5;

wire[31:0] addr_1021_5;

Selector_2 s1021_5(wires_255_4[1], addr_255_4, wires_1021_5,addr_1021_5);

wire[3:0] wires_1022_5;

wire[31:0] addr_1022_5;

Selector_2 s1022_5(wires_255_4[2], addr_255_4, wires_1022_5,addr_1022_5);

wire[3:0] wires_1023_5;

wire[31:0] addr_1023_5;

Selector_2 s1023_5(wires_255_4[3], addr_255_4, wires_1023_5,addr_1023_5);

wire[3:0] wires_0_6;

wire[31:0] addr_0_6;

Selector_2 s0_6(wires_0_5[0], addr_0_5, wires_0_6,addr_0_6);

wire[3:0] wires_1_6;

wire[31:0] addr_1_6;

Selector_2 s1_6(wires_0_5[1], addr_0_5, wires_1_6,addr_1_6);

wire[3:0] wires_2_6;

wire[31:0] addr_2_6;

Selector_2 s2_6(wires_0_5[2], addr_0_5, wires_2_6,addr_2_6);

wire[3:0] wires_3_6;

wire[31:0] addr_3_6;

Selector_2 s3_6(wires_0_5[3], addr_0_5, wires_3_6,addr_3_6);

wire[3:0] wires_4_6;

wire[31:0] addr_4_6;

Selector_2 s4_6(wires_1_5[0], addr_1_5, wires_4_6,addr_4_6);

wire[3:0] wires_5_6;

wire[31:0] addr_5_6;

Selector_2 s5_6(wires_1_5[1], addr_1_5, wires_5_6,addr_5_6);

wire[3:0] wires_6_6;

wire[31:0] addr_6_6;

Selector_2 s6_6(wires_1_5[2], addr_1_5, wires_6_6,addr_6_6);

wire[3:0] wires_7_6;

wire[31:0] addr_7_6;

Selector_2 s7_6(wires_1_5[3], addr_1_5, wires_7_6,addr_7_6);

wire[3:0] wires_8_6;

wire[31:0] addr_8_6;

Selector_2 s8_6(wires_2_5[0], addr_2_5, wires_8_6,addr_8_6);

wire[3:0] wires_9_6;

wire[31:0] addr_9_6;

Selector_2 s9_6(wires_2_5[1], addr_2_5, wires_9_6,addr_9_6);

wire[3:0] wires_10_6;

wire[31:0] addr_10_6;

Selector_2 s10_6(wires_2_5[2], addr_2_5, wires_10_6,addr_10_6);

wire[3:0] wires_11_6;

wire[31:0] addr_11_6;

Selector_2 s11_6(wires_2_5[3], addr_2_5, wires_11_6,addr_11_6);

wire[3:0] wires_12_6;

wire[31:0] addr_12_6;

Selector_2 s12_6(wires_3_5[0], addr_3_5, wires_12_6,addr_12_6);

wire[3:0] wires_13_6;

wire[31:0] addr_13_6;

Selector_2 s13_6(wires_3_5[1], addr_3_5, wires_13_6,addr_13_6);

wire[3:0] wires_14_6;

wire[31:0] addr_14_6;

Selector_2 s14_6(wires_3_5[2], addr_3_5, wires_14_6,addr_14_6);

wire[3:0] wires_15_6;

wire[31:0] addr_15_6;

Selector_2 s15_6(wires_3_5[3], addr_3_5, wires_15_6,addr_15_6);

wire[3:0] wires_16_6;

wire[31:0] addr_16_6;

Selector_2 s16_6(wires_4_5[0], addr_4_5, wires_16_6,addr_16_6);

wire[3:0] wires_17_6;

wire[31:0] addr_17_6;

Selector_2 s17_6(wires_4_5[1], addr_4_5, wires_17_6,addr_17_6);

wire[3:0] wires_18_6;

wire[31:0] addr_18_6;

Selector_2 s18_6(wires_4_5[2], addr_4_5, wires_18_6,addr_18_6);

wire[3:0] wires_19_6;

wire[31:0] addr_19_6;

Selector_2 s19_6(wires_4_5[3], addr_4_5, wires_19_6,addr_19_6);

wire[3:0] wires_20_6;

wire[31:0] addr_20_6;

Selector_2 s20_6(wires_5_5[0], addr_5_5, wires_20_6,addr_20_6);

wire[3:0] wires_21_6;

wire[31:0] addr_21_6;

Selector_2 s21_6(wires_5_5[1], addr_5_5, wires_21_6,addr_21_6);

wire[3:0] wires_22_6;

wire[31:0] addr_22_6;

Selector_2 s22_6(wires_5_5[2], addr_5_5, wires_22_6,addr_22_6);

wire[3:0] wires_23_6;

wire[31:0] addr_23_6;

Selector_2 s23_6(wires_5_5[3], addr_5_5, wires_23_6,addr_23_6);

wire[3:0] wires_24_6;

wire[31:0] addr_24_6;

Selector_2 s24_6(wires_6_5[0], addr_6_5, wires_24_6,addr_24_6);

wire[3:0] wires_25_6;

wire[31:0] addr_25_6;

Selector_2 s25_6(wires_6_5[1], addr_6_5, wires_25_6,addr_25_6);

wire[3:0] wires_26_6;

wire[31:0] addr_26_6;

Selector_2 s26_6(wires_6_5[2], addr_6_5, wires_26_6,addr_26_6);

wire[3:0] wires_27_6;

wire[31:0] addr_27_6;

Selector_2 s27_6(wires_6_5[3], addr_6_5, wires_27_6,addr_27_6);

wire[3:0] wires_28_6;

wire[31:0] addr_28_6;

Selector_2 s28_6(wires_7_5[0], addr_7_5, wires_28_6,addr_28_6);

wire[3:0] wires_29_6;

wire[31:0] addr_29_6;

Selector_2 s29_6(wires_7_5[1], addr_7_5, wires_29_6,addr_29_6);

wire[3:0] wires_30_6;

wire[31:0] addr_30_6;

Selector_2 s30_6(wires_7_5[2], addr_7_5, wires_30_6,addr_30_6);

wire[3:0] wires_31_6;

wire[31:0] addr_31_6;

Selector_2 s31_6(wires_7_5[3], addr_7_5, wires_31_6,addr_31_6);

wire[3:0] wires_32_6;

wire[31:0] addr_32_6;

Selector_2 s32_6(wires_8_5[0], addr_8_5, wires_32_6,addr_32_6);

wire[3:0] wires_33_6;

wire[31:0] addr_33_6;

Selector_2 s33_6(wires_8_5[1], addr_8_5, wires_33_6,addr_33_6);

wire[3:0] wires_34_6;

wire[31:0] addr_34_6;

Selector_2 s34_6(wires_8_5[2], addr_8_5, wires_34_6,addr_34_6);

wire[3:0] wires_35_6;

wire[31:0] addr_35_6;

Selector_2 s35_6(wires_8_5[3], addr_8_5, wires_35_6,addr_35_6);

wire[3:0] wires_36_6;

wire[31:0] addr_36_6;

Selector_2 s36_6(wires_9_5[0], addr_9_5, wires_36_6,addr_36_6);

wire[3:0] wires_37_6;

wire[31:0] addr_37_6;

Selector_2 s37_6(wires_9_5[1], addr_9_5, wires_37_6,addr_37_6);

wire[3:0] wires_38_6;

wire[31:0] addr_38_6;

Selector_2 s38_6(wires_9_5[2], addr_9_5, wires_38_6,addr_38_6);

wire[3:0] wires_39_6;

wire[31:0] addr_39_6;

Selector_2 s39_6(wires_9_5[3], addr_9_5, wires_39_6,addr_39_6);

wire[3:0] wires_40_6;

wire[31:0] addr_40_6;

Selector_2 s40_6(wires_10_5[0], addr_10_5, wires_40_6,addr_40_6);

wire[3:0] wires_41_6;

wire[31:0] addr_41_6;

Selector_2 s41_6(wires_10_5[1], addr_10_5, wires_41_6,addr_41_6);

wire[3:0] wires_42_6;

wire[31:0] addr_42_6;

Selector_2 s42_6(wires_10_5[2], addr_10_5, wires_42_6,addr_42_6);

wire[3:0] wires_43_6;

wire[31:0] addr_43_6;

Selector_2 s43_6(wires_10_5[3], addr_10_5, wires_43_6,addr_43_6);

wire[3:0] wires_44_6;

wire[31:0] addr_44_6;

Selector_2 s44_6(wires_11_5[0], addr_11_5, wires_44_6,addr_44_6);

wire[3:0] wires_45_6;

wire[31:0] addr_45_6;

Selector_2 s45_6(wires_11_5[1], addr_11_5, wires_45_6,addr_45_6);

wire[3:0] wires_46_6;

wire[31:0] addr_46_6;

Selector_2 s46_6(wires_11_5[2], addr_11_5, wires_46_6,addr_46_6);

wire[3:0] wires_47_6;

wire[31:0] addr_47_6;

Selector_2 s47_6(wires_11_5[3], addr_11_5, wires_47_6,addr_47_6);

wire[3:0] wires_48_6;

wire[31:0] addr_48_6;

Selector_2 s48_6(wires_12_5[0], addr_12_5, wires_48_6,addr_48_6);

wire[3:0] wires_49_6;

wire[31:0] addr_49_6;

Selector_2 s49_6(wires_12_5[1], addr_12_5, wires_49_6,addr_49_6);

wire[3:0] wires_50_6;

wire[31:0] addr_50_6;

Selector_2 s50_6(wires_12_5[2], addr_12_5, wires_50_6,addr_50_6);

wire[3:0] wires_51_6;

wire[31:0] addr_51_6;

Selector_2 s51_6(wires_12_5[3], addr_12_5, wires_51_6,addr_51_6);

wire[3:0] wires_52_6;

wire[31:0] addr_52_6;

Selector_2 s52_6(wires_13_5[0], addr_13_5, wires_52_6,addr_52_6);

wire[3:0] wires_53_6;

wire[31:0] addr_53_6;

Selector_2 s53_6(wires_13_5[1], addr_13_5, wires_53_6,addr_53_6);

wire[3:0] wires_54_6;

wire[31:0] addr_54_6;

Selector_2 s54_6(wires_13_5[2], addr_13_5, wires_54_6,addr_54_6);

wire[3:0] wires_55_6;

wire[31:0] addr_55_6;

Selector_2 s55_6(wires_13_5[3], addr_13_5, wires_55_6,addr_55_6);

wire[3:0] wires_56_6;

wire[31:0] addr_56_6;

Selector_2 s56_6(wires_14_5[0], addr_14_5, wires_56_6,addr_56_6);

wire[3:0] wires_57_6;

wire[31:0] addr_57_6;

Selector_2 s57_6(wires_14_5[1], addr_14_5, wires_57_6,addr_57_6);

wire[3:0] wires_58_6;

wire[31:0] addr_58_6;

Selector_2 s58_6(wires_14_5[2], addr_14_5, wires_58_6,addr_58_6);

wire[3:0] wires_59_6;

wire[31:0] addr_59_6;

Selector_2 s59_6(wires_14_5[3], addr_14_5, wires_59_6,addr_59_6);

wire[3:0] wires_60_6;

wire[31:0] addr_60_6;

Selector_2 s60_6(wires_15_5[0], addr_15_5, wires_60_6,addr_60_6);

wire[3:0] wires_61_6;

wire[31:0] addr_61_6;

Selector_2 s61_6(wires_15_5[1], addr_15_5, wires_61_6,addr_61_6);

wire[3:0] wires_62_6;

wire[31:0] addr_62_6;

Selector_2 s62_6(wires_15_5[2], addr_15_5, wires_62_6,addr_62_6);

wire[3:0] wires_63_6;

wire[31:0] addr_63_6;

Selector_2 s63_6(wires_15_5[3], addr_15_5, wires_63_6,addr_63_6);

wire[3:0] wires_64_6;

wire[31:0] addr_64_6;

Selector_2 s64_6(wires_16_5[0], addr_16_5, wires_64_6,addr_64_6);

wire[3:0] wires_65_6;

wire[31:0] addr_65_6;

Selector_2 s65_6(wires_16_5[1], addr_16_5, wires_65_6,addr_65_6);

wire[3:0] wires_66_6;

wire[31:0] addr_66_6;

Selector_2 s66_6(wires_16_5[2], addr_16_5, wires_66_6,addr_66_6);

wire[3:0] wires_67_6;

wire[31:0] addr_67_6;

Selector_2 s67_6(wires_16_5[3], addr_16_5, wires_67_6,addr_67_6);

wire[3:0] wires_68_6;

wire[31:0] addr_68_6;

Selector_2 s68_6(wires_17_5[0], addr_17_5, wires_68_6,addr_68_6);

wire[3:0] wires_69_6;

wire[31:0] addr_69_6;

Selector_2 s69_6(wires_17_5[1], addr_17_5, wires_69_6,addr_69_6);

wire[3:0] wires_70_6;

wire[31:0] addr_70_6;

Selector_2 s70_6(wires_17_5[2], addr_17_5, wires_70_6,addr_70_6);

wire[3:0] wires_71_6;

wire[31:0] addr_71_6;

Selector_2 s71_6(wires_17_5[3], addr_17_5, wires_71_6,addr_71_6);

wire[3:0] wires_72_6;

wire[31:0] addr_72_6;

Selector_2 s72_6(wires_18_5[0], addr_18_5, wires_72_6,addr_72_6);

wire[3:0] wires_73_6;

wire[31:0] addr_73_6;

Selector_2 s73_6(wires_18_5[1], addr_18_5, wires_73_6,addr_73_6);

wire[3:0] wires_74_6;

wire[31:0] addr_74_6;

Selector_2 s74_6(wires_18_5[2], addr_18_5, wires_74_6,addr_74_6);

wire[3:0] wires_75_6;

wire[31:0] addr_75_6;

Selector_2 s75_6(wires_18_5[3], addr_18_5, wires_75_6,addr_75_6);

wire[3:0] wires_76_6;

wire[31:0] addr_76_6;

Selector_2 s76_6(wires_19_5[0], addr_19_5, wires_76_6,addr_76_6);

wire[3:0] wires_77_6;

wire[31:0] addr_77_6;

Selector_2 s77_6(wires_19_5[1], addr_19_5, wires_77_6,addr_77_6);

wire[3:0] wires_78_6;

wire[31:0] addr_78_6;

Selector_2 s78_6(wires_19_5[2], addr_19_5, wires_78_6,addr_78_6);

wire[3:0] wires_79_6;

wire[31:0] addr_79_6;

Selector_2 s79_6(wires_19_5[3], addr_19_5, wires_79_6,addr_79_6);

wire[3:0] wires_80_6;

wire[31:0] addr_80_6;

Selector_2 s80_6(wires_20_5[0], addr_20_5, wires_80_6,addr_80_6);

wire[3:0] wires_81_6;

wire[31:0] addr_81_6;

Selector_2 s81_6(wires_20_5[1], addr_20_5, wires_81_6,addr_81_6);

wire[3:0] wires_82_6;

wire[31:0] addr_82_6;

Selector_2 s82_6(wires_20_5[2], addr_20_5, wires_82_6,addr_82_6);

wire[3:0] wires_83_6;

wire[31:0] addr_83_6;

Selector_2 s83_6(wires_20_5[3], addr_20_5, wires_83_6,addr_83_6);

wire[3:0] wires_84_6;

wire[31:0] addr_84_6;

Selector_2 s84_6(wires_21_5[0], addr_21_5, wires_84_6,addr_84_6);

wire[3:0] wires_85_6;

wire[31:0] addr_85_6;

Selector_2 s85_6(wires_21_5[1], addr_21_5, wires_85_6,addr_85_6);

wire[3:0] wires_86_6;

wire[31:0] addr_86_6;

Selector_2 s86_6(wires_21_5[2], addr_21_5, wires_86_6,addr_86_6);

wire[3:0] wires_87_6;

wire[31:0] addr_87_6;

Selector_2 s87_6(wires_21_5[3], addr_21_5, wires_87_6,addr_87_6);

wire[3:0] wires_88_6;

wire[31:0] addr_88_6;

Selector_2 s88_6(wires_22_5[0], addr_22_5, wires_88_6,addr_88_6);

wire[3:0] wires_89_6;

wire[31:0] addr_89_6;

Selector_2 s89_6(wires_22_5[1], addr_22_5, wires_89_6,addr_89_6);

wire[3:0] wires_90_6;

wire[31:0] addr_90_6;

Selector_2 s90_6(wires_22_5[2], addr_22_5, wires_90_6,addr_90_6);

wire[3:0] wires_91_6;

wire[31:0] addr_91_6;

Selector_2 s91_6(wires_22_5[3], addr_22_5, wires_91_6,addr_91_6);

wire[3:0] wires_92_6;

wire[31:0] addr_92_6;

Selector_2 s92_6(wires_23_5[0], addr_23_5, wires_92_6,addr_92_6);

wire[3:0] wires_93_6;

wire[31:0] addr_93_6;

Selector_2 s93_6(wires_23_5[1], addr_23_5, wires_93_6,addr_93_6);

wire[3:0] wires_94_6;

wire[31:0] addr_94_6;

Selector_2 s94_6(wires_23_5[2], addr_23_5, wires_94_6,addr_94_6);

wire[3:0] wires_95_6;

wire[31:0] addr_95_6;

Selector_2 s95_6(wires_23_5[3], addr_23_5, wires_95_6,addr_95_6);

wire[3:0] wires_96_6;

wire[31:0] addr_96_6;

Selector_2 s96_6(wires_24_5[0], addr_24_5, wires_96_6,addr_96_6);

wire[3:0] wires_97_6;

wire[31:0] addr_97_6;

Selector_2 s97_6(wires_24_5[1], addr_24_5, wires_97_6,addr_97_6);

wire[3:0] wires_98_6;

wire[31:0] addr_98_6;

Selector_2 s98_6(wires_24_5[2], addr_24_5, wires_98_6,addr_98_6);

wire[3:0] wires_99_6;

wire[31:0] addr_99_6;

Selector_2 s99_6(wires_24_5[3], addr_24_5, wires_99_6,addr_99_6);

wire[3:0] wires_100_6;

wire[31:0] addr_100_6;

Selector_2 s100_6(wires_25_5[0], addr_25_5, wires_100_6,addr_100_6);

wire[3:0] wires_101_6;

wire[31:0] addr_101_6;

Selector_2 s101_6(wires_25_5[1], addr_25_5, wires_101_6,addr_101_6);

wire[3:0] wires_102_6;

wire[31:0] addr_102_6;

Selector_2 s102_6(wires_25_5[2], addr_25_5, wires_102_6,addr_102_6);

wire[3:0] wires_103_6;

wire[31:0] addr_103_6;

Selector_2 s103_6(wires_25_5[3], addr_25_5, wires_103_6,addr_103_6);

wire[3:0] wires_104_6;

wire[31:0] addr_104_6;

Selector_2 s104_6(wires_26_5[0], addr_26_5, wires_104_6,addr_104_6);

wire[3:0] wires_105_6;

wire[31:0] addr_105_6;

Selector_2 s105_6(wires_26_5[1], addr_26_5, wires_105_6,addr_105_6);

wire[3:0] wires_106_6;

wire[31:0] addr_106_6;

Selector_2 s106_6(wires_26_5[2], addr_26_5, wires_106_6,addr_106_6);

wire[3:0] wires_107_6;

wire[31:0] addr_107_6;

Selector_2 s107_6(wires_26_5[3], addr_26_5, wires_107_6,addr_107_6);

wire[3:0] wires_108_6;

wire[31:0] addr_108_6;

Selector_2 s108_6(wires_27_5[0], addr_27_5, wires_108_6,addr_108_6);

wire[3:0] wires_109_6;

wire[31:0] addr_109_6;

Selector_2 s109_6(wires_27_5[1], addr_27_5, wires_109_6,addr_109_6);

wire[3:0] wires_110_6;

wire[31:0] addr_110_6;

Selector_2 s110_6(wires_27_5[2], addr_27_5, wires_110_6,addr_110_6);

wire[3:0] wires_111_6;

wire[31:0] addr_111_6;

Selector_2 s111_6(wires_27_5[3], addr_27_5, wires_111_6,addr_111_6);

wire[3:0] wires_112_6;

wire[31:0] addr_112_6;

Selector_2 s112_6(wires_28_5[0], addr_28_5, wires_112_6,addr_112_6);

wire[3:0] wires_113_6;

wire[31:0] addr_113_6;

Selector_2 s113_6(wires_28_5[1], addr_28_5, wires_113_6,addr_113_6);

wire[3:0] wires_114_6;

wire[31:0] addr_114_6;

Selector_2 s114_6(wires_28_5[2], addr_28_5, wires_114_6,addr_114_6);

wire[3:0] wires_115_6;

wire[31:0] addr_115_6;

Selector_2 s115_6(wires_28_5[3], addr_28_5, wires_115_6,addr_115_6);

wire[3:0] wires_116_6;

wire[31:0] addr_116_6;

Selector_2 s116_6(wires_29_5[0], addr_29_5, wires_116_6,addr_116_6);

wire[3:0] wires_117_6;

wire[31:0] addr_117_6;

Selector_2 s117_6(wires_29_5[1], addr_29_5, wires_117_6,addr_117_6);

wire[3:0] wires_118_6;

wire[31:0] addr_118_6;

Selector_2 s118_6(wires_29_5[2], addr_29_5, wires_118_6,addr_118_6);

wire[3:0] wires_119_6;

wire[31:0] addr_119_6;

Selector_2 s119_6(wires_29_5[3], addr_29_5, wires_119_6,addr_119_6);

wire[3:0] wires_120_6;

wire[31:0] addr_120_6;

Selector_2 s120_6(wires_30_5[0], addr_30_5, wires_120_6,addr_120_6);

wire[3:0] wires_121_6;

wire[31:0] addr_121_6;

Selector_2 s121_6(wires_30_5[1], addr_30_5, wires_121_6,addr_121_6);

wire[3:0] wires_122_6;

wire[31:0] addr_122_6;

Selector_2 s122_6(wires_30_5[2], addr_30_5, wires_122_6,addr_122_6);

wire[3:0] wires_123_6;

wire[31:0] addr_123_6;

Selector_2 s123_6(wires_30_5[3], addr_30_5, wires_123_6,addr_123_6);

wire[3:0] wires_124_6;

wire[31:0] addr_124_6;

Selector_2 s124_6(wires_31_5[0], addr_31_5, wires_124_6,addr_124_6);

wire[3:0] wires_125_6;

wire[31:0] addr_125_6;

Selector_2 s125_6(wires_31_5[1], addr_31_5, wires_125_6,addr_125_6);

wire[3:0] wires_126_6;

wire[31:0] addr_126_6;

Selector_2 s126_6(wires_31_5[2], addr_31_5, wires_126_6,addr_126_6);

wire[3:0] wires_127_6;

wire[31:0] addr_127_6;

Selector_2 s127_6(wires_31_5[3], addr_31_5, wires_127_6,addr_127_6);

wire[3:0] wires_128_6;

wire[31:0] addr_128_6;

Selector_2 s128_6(wires_32_5[0], addr_32_5, wires_128_6,addr_128_6);

wire[3:0] wires_129_6;

wire[31:0] addr_129_6;

Selector_2 s129_6(wires_32_5[1], addr_32_5, wires_129_6,addr_129_6);

wire[3:0] wires_130_6;

wire[31:0] addr_130_6;

Selector_2 s130_6(wires_32_5[2], addr_32_5, wires_130_6,addr_130_6);

wire[3:0] wires_131_6;

wire[31:0] addr_131_6;

Selector_2 s131_6(wires_32_5[3], addr_32_5, wires_131_6,addr_131_6);

wire[3:0] wires_132_6;

wire[31:0] addr_132_6;

Selector_2 s132_6(wires_33_5[0], addr_33_5, wires_132_6,addr_132_6);

wire[3:0] wires_133_6;

wire[31:0] addr_133_6;

Selector_2 s133_6(wires_33_5[1], addr_33_5, wires_133_6,addr_133_6);

wire[3:0] wires_134_6;

wire[31:0] addr_134_6;

Selector_2 s134_6(wires_33_5[2], addr_33_5, wires_134_6,addr_134_6);

wire[3:0] wires_135_6;

wire[31:0] addr_135_6;

Selector_2 s135_6(wires_33_5[3], addr_33_5, wires_135_6,addr_135_6);

wire[3:0] wires_136_6;

wire[31:0] addr_136_6;

Selector_2 s136_6(wires_34_5[0], addr_34_5, wires_136_6,addr_136_6);

wire[3:0] wires_137_6;

wire[31:0] addr_137_6;

Selector_2 s137_6(wires_34_5[1], addr_34_5, wires_137_6,addr_137_6);

wire[3:0] wires_138_6;

wire[31:0] addr_138_6;

Selector_2 s138_6(wires_34_5[2], addr_34_5, wires_138_6,addr_138_6);

wire[3:0] wires_139_6;

wire[31:0] addr_139_6;

Selector_2 s139_6(wires_34_5[3], addr_34_5, wires_139_6,addr_139_6);

wire[3:0] wires_140_6;

wire[31:0] addr_140_6;

Selector_2 s140_6(wires_35_5[0], addr_35_5, wires_140_6,addr_140_6);

wire[3:0] wires_141_6;

wire[31:0] addr_141_6;

Selector_2 s141_6(wires_35_5[1], addr_35_5, wires_141_6,addr_141_6);

wire[3:0] wires_142_6;

wire[31:0] addr_142_6;

Selector_2 s142_6(wires_35_5[2], addr_35_5, wires_142_6,addr_142_6);

wire[3:0] wires_143_6;

wire[31:0] addr_143_6;

Selector_2 s143_6(wires_35_5[3], addr_35_5, wires_143_6,addr_143_6);

wire[3:0] wires_144_6;

wire[31:0] addr_144_6;

Selector_2 s144_6(wires_36_5[0], addr_36_5, wires_144_6,addr_144_6);

wire[3:0] wires_145_6;

wire[31:0] addr_145_6;

Selector_2 s145_6(wires_36_5[1], addr_36_5, wires_145_6,addr_145_6);

wire[3:0] wires_146_6;

wire[31:0] addr_146_6;

Selector_2 s146_6(wires_36_5[2], addr_36_5, wires_146_6,addr_146_6);

wire[3:0] wires_147_6;

wire[31:0] addr_147_6;

Selector_2 s147_6(wires_36_5[3], addr_36_5, wires_147_6,addr_147_6);

wire[3:0] wires_148_6;

wire[31:0] addr_148_6;

Selector_2 s148_6(wires_37_5[0], addr_37_5, wires_148_6,addr_148_6);

wire[3:0] wires_149_6;

wire[31:0] addr_149_6;

Selector_2 s149_6(wires_37_5[1], addr_37_5, wires_149_6,addr_149_6);

wire[3:0] wires_150_6;

wire[31:0] addr_150_6;

Selector_2 s150_6(wires_37_5[2], addr_37_5, wires_150_6,addr_150_6);

wire[3:0] wires_151_6;

wire[31:0] addr_151_6;

Selector_2 s151_6(wires_37_5[3], addr_37_5, wires_151_6,addr_151_6);

wire[3:0] wires_152_6;

wire[31:0] addr_152_6;

Selector_2 s152_6(wires_38_5[0], addr_38_5, wires_152_6,addr_152_6);

wire[3:0] wires_153_6;

wire[31:0] addr_153_6;

Selector_2 s153_6(wires_38_5[1], addr_38_5, wires_153_6,addr_153_6);

wire[3:0] wires_154_6;

wire[31:0] addr_154_6;

Selector_2 s154_6(wires_38_5[2], addr_38_5, wires_154_6,addr_154_6);

wire[3:0] wires_155_6;

wire[31:0] addr_155_6;

Selector_2 s155_6(wires_38_5[3], addr_38_5, wires_155_6,addr_155_6);

wire[3:0] wires_156_6;

wire[31:0] addr_156_6;

Selector_2 s156_6(wires_39_5[0], addr_39_5, wires_156_6,addr_156_6);

wire[3:0] wires_157_6;

wire[31:0] addr_157_6;

Selector_2 s157_6(wires_39_5[1], addr_39_5, wires_157_6,addr_157_6);

wire[3:0] wires_158_6;

wire[31:0] addr_158_6;

Selector_2 s158_6(wires_39_5[2], addr_39_5, wires_158_6,addr_158_6);

wire[3:0] wires_159_6;

wire[31:0] addr_159_6;

Selector_2 s159_6(wires_39_5[3], addr_39_5, wires_159_6,addr_159_6);

wire[3:0] wires_160_6;

wire[31:0] addr_160_6;

Selector_2 s160_6(wires_40_5[0], addr_40_5, wires_160_6,addr_160_6);

wire[3:0] wires_161_6;

wire[31:0] addr_161_6;

Selector_2 s161_6(wires_40_5[1], addr_40_5, wires_161_6,addr_161_6);

wire[3:0] wires_162_6;

wire[31:0] addr_162_6;

Selector_2 s162_6(wires_40_5[2], addr_40_5, wires_162_6,addr_162_6);

wire[3:0] wires_163_6;

wire[31:0] addr_163_6;

Selector_2 s163_6(wires_40_5[3], addr_40_5, wires_163_6,addr_163_6);

wire[3:0] wires_164_6;

wire[31:0] addr_164_6;

Selector_2 s164_6(wires_41_5[0], addr_41_5, wires_164_6,addr_164_6);

wire[3:0] wires_165_6;

wire[31:0] addr_165_6;

Selector_2 s165_6(wires_41_5[1], addr_41_5, wires_165_6,addr_165_6);

wire[3:0] wires_166_6;

wire[31:0] addr_166_6;

Selector_2 s166_6(wires_41_5[2], addr_41_5, wires_166_6,addr_166_6);

wire[3:0] wires_167_6;

wire[31:0] addr_167_6;

Selector_2 s167_6(wires_41_5[3], addr_41_5, wires_167_6,addr_167_6);

wire[3:0] wires_168_6;

wire[31:0] addr_168_6;

Selector_2 s168_6(wires_42_5[0], addr_42_5, wires_168_6,addr_168_6);

wire[3:0] wires_169_6;

wire[31:0] addr_169_6;

Selector_2 s169_6(wires_42_5[1], addr_42_5, wires_169_6,addr_169_6);

wire[3:0] wires_170_6;

wire[31:0] addr_170_6;

Selector_2 s170_6(wires_42_5[2], addr_42_5, wires_170_6,addr_170_6);

wire[3:0] wires_171_6;

wire[31:0] addr_171_6;

Selector_2 s171_6(wires_42_5[3], addr_42_5, wires_171_6,addr_171_6);

wire[3:0] wires_172_6;

wire[31:0] addr_172_6;

Selector_2 s172_6(wires_43_5[0], addr_43_5, wires_172_6,addr_172_6);

wire[3:0] wires_173_6;

wire[31:0] addr_173_6;

Selector_2 s173_6(wires_43_5[1], addr_43_5, wires_173_6,addr_173_6);

wire[3:0] wires_174_6;

wire[31:0] addr_174_6;

Selector_2 s174_6(wires_43_5[2], addr_43_5, wires_174_6,addr_174_6);

wire[3:0] wires_175_6;

wire[31:0] addr_175_6;

Selector_2 s175_6(wires_43_5[3], addr_43_5, wires_175_6,addr_175_6);

wire[3:0] wires_176_6;

wire[31:0] addr_176_6;

Selector_2 s176_6(wires_44_5[0], addr_44_5, wires_176_6,addr_176_6);

wire[3:0] wires_177_6;

wire[31:0] addr_177_6;

Selector_2 s177_6(wires_44_5[1], addr_44_5, wires_177_6,addr_177_6);

wire[3:0] wires_178_6;

wire[31:0] addr_178_6;

Selector_2 s178_6(wires_44_5[2], addr_44_5, wires_178_6,addr_178_6);

wire[3:0] wires_179_6;

wire[31:0] addr_179_6;

Selector_2 s179_6(wires_44_5[3], addr_44_5, wires_179_6,addr_179_6);

wire[3:0] wires_180_6;

wire[31:0] addr_180_6;

Selector_2 s180_6(wires_45_5[0], addr_45_5, wires_180_6,addr_180_6);

wire[3:0] wires_181_6;

wire[31:0] addr_181_6;

Selector_2 s181_6(wires_45_5[1], addr_45_5, wires_181_6,addr_181_6);

wire[3:0] wires_182_6;

wire[31:0] addr_182_6;

Selector_2 s182_6(wires_45_5[2], addr_45_5, wires_182_6,addr_182_6);

wire[3:0] wires_183_6;

wire[31:0] addr_183_6;

Selector_2 s183_6(wires_45_5[3], addr_45_5, wires_183_6,addr_183_6);

wire[3:0] wires_184_6;

wire[31:0] addr_184_6;

Selector_2 s184_6(wires_46_5[0], addr_46_5, wires_184_6,addr_184_6);

wire[3:0] wires_185_6;

wire[31:0] addr_185_6;

Selector_2 s185_6(wires_46_5[1], addr_46_5, wires_185_6,addr_185_6);

wire[3:0] wires_186_6;

wire[31:0] addr_186_6;

Selector_2 s186_6(wires_46_5[2], addr_46_5, wires_186_6,addr_186_6);

wire[3:0] wires_187_6;

wire[31:0] addr_187_6;

Selector_2 s187_6(wires_46_5[3], addr_46_5, wires_187_6,addr_187_6);

wire[3:0] wires_188_6;

wire[31:0] addr_188_6;

Selector_2 s188_6(wires_47_5[0], addr_47_5, wires_188_6,addr_188_6);

wire[3:0] wires_189_6;

wire[31:0] addr_189_6;

Selector_2 s189_6(wires_47_5[1], addr_47_5, wires_189_6,addr_189_6);

wire[3:0] wires_190_6;

wire[31:0] addr_190_6;

Selector_2 s190_6(wires_47_5[2], addr_47_5, wires_190_6,addr_190_6);

wire[3:0] wires_191_6;

wire[31:0] addr_191_6;

Selector_2 s191_6(wires_47_5[3], addr_47_5, wires_191_6,addr_191_6);

wire[3:0] wires_192_6;

wire[31:0] addr_192_6;

Selector_2 s192_6(wires_48_5[0], addr_48_5, wires_192_6,addr_192_6);

wire[3:0] wires_193_6;

wire[31:0] addr_193_6;

Selector_2 s193_6(wires_48_5[1], addr_48_5, wires_193_6,addr_193_6);

wire[3:0] wires_194_6;

wire[31:0] addr_194_6;

Selector_2 s194_6(wires_48_5[2], addr_48_5, wires_194_6,addr_194_6);

wire[3:0] wires_195_6;

wire[31:0] addr_195_6;

Selector_2 s195_6(wires_48_5[3], addr_48_5, wires_195_6,addr_195_6);

wire[3:0] wires_196_6;

wire[31:0] addr_196_6;

Selector_2 s196_6(wires_49_5[0], addr_49_5, wires_196_6,addr_196_6);

wire[3:0] wires_197_6;

wire[31:0] addr_197_6;

Selector_2 s197_6(wires_49_5[1], addr_49_5, wires_197_6,addr_197_6);

wire[3:0] wires_198_6;

wire[31:0] addr_198_6;

Selector_2 s198_6(wires_49_5[2], addr_49_5, wires_198_6,addr_198_6);

wire[3:0] wires_199_6;

wire[31:0] addr_199_6;

Selector_2 s199_6(wires_49_5[3], addr_49_5, wires_199_6,addr_199_6);

wire[3:0] wires_200_6;

wire[31:0] addr_200_6;

Selector_2 s200_6(wires_50_5[0], addr_50_5, wires_200_6,addr_200_6);

wire[3:0] wires_201_6;

wire[31:0] addr_201_6;

Selector_2 s201_6(wires_50_5[1], addr_50_5, wires_201_6,addr_201_6);

wire[3:0] wires_202_6;

wire[31:0] addr_202_6;

Selector_2 s202_6(wires_50_5[2], addr_50_5, wires_202_6,addr_202_6);

wire[3:0] wires_203_6;

wire[31:0] addr_203_6;

Selector_2 s203_6(wires_50_5[3], addr_50_5, wires_203_6,addr_203_6);

wire[3:0] wires_204_6;

wire[31:0] addr_204_6;

Selector_2 s204_6(wires_51_5[0], addr_51_5, wires_204_6,addr_204_6);

wire[3:0] wires_205_6;

wire[31:0] addr_205_6;

Selector_2 s205_6(wires_51_5[1], addr_51_5, wires_205_6,addr_205_6);

wire[3:0] wires_206_6;

wire[31:0] addr_206_6;

Selector_2 s206_6(wires_51_5[2], addr_51_5, wires_206_6,addr_206_6);

wire[3:0] wires_207_6;

wire[31:0] addr_207_6;

Selector_2 s207_6(wires_51_5[3], addr_51_5, wires_207_6,addr_207_6);

wire[3:0] wires_208_6;

wire[31:0] addr_208_6;

Selector_2 s208_6(wires_52_5[0], addr_52_5, wires_208_6,addr_208_6);

wire[3:0] wires_209_6;

wire[31:0] addr_209_6;

Selector_2 s209_6(wires_52_5[1], addr_52_5, wires_209_6,addr_209_6);

wire[3:0] wires_210_6;

wire[31:0] addr_210_6;

Selector_2 s210_6(wires_52_5[2], addr_52_5, wires_210_6,addr_210_6);

wire[3:0] wires_211_6;

wire[31:0] addr_211_6;

Selector_2 s211_6(wires_52_5[3], addr_52_5, wires_211_6,addr_211_6);

wire[3:0] wires_212_6;

wire[31:0] addr_212_6;

Selector_2 s212_6(wires_53_5[0], addr_53_5, wires_212_6,addr_212_6);

wire[3:0] wires_213_6;

wire[31:0] addr_213_6;

Selector_2 s213_6(wires_53_5[1], addr_53_5, wires_213_6,addr_213_6);

wire[3:0] wires_214_6;

wire[31:0] addr_214_6;

Selector_2 s214_6(wires_53_5[2], addr_53_5, wires_214_6,addr_214_6);

wire[3:0] wires_215_6;

wire[31:0] addr_215_6;

Selector_2 s215_6(wires_53_5[3], addr_53_5, wires_215_6,addr_215_6);

wire[3:0] wires_216_6;

wire[31:0] addr_216_6;

Selector_2 s216_6(wires_54_5[0], addr_54_5, wires_216_6,addr_216_6);

wire[3:0] wires_217_6;

wire[31:0] addr_217_6;

Selector_2 s217_6(wires_54_5[1], addr_54_5, wires_217_6,addr_217_6);

wire[3:0] wires_218_6;

wire[31:0] addr_218_6;

Selector_2 s218_6(wires_54_5[2], addr_54_5, wires_218_6,addr_218_6);

wire[3:0] wires_219_6;

wire[31:0] addr_219_6;

Selector_2 s219_6(wires_54_5[3], addr_54_5, wires_219_6,addr_219_6);

wire[3:0] wires_220_6;

wire[31:0] addr_220_6;

Selector_2 s220_6(wires_55_5[0], addr_55_5, wires_220_6,addr_220_6);

wire[3:0] wires_221_6;

wire[31:0] addr_221_6;

Selector_2 s221_6(wires_55_5[1], addr_55_5, wires_221_6,addr_221_6);

wire[3:0] wires_222_6;

wire[31:0] addr_222_6;

Selector_2 s222_6(wires_55_5[2], addr_55_5, wires_222_6,addr_222_6);

wire[3:0] wires_223_6;

wire[31:0] addr_223_6;

Selector_2 s223_6(wires_55_5[3], addr_55_5, wires_223_6,addr_223_6);

wire[3:0] wires_224_6;

wire[31:0] addr_224_6;

Selector_2 s224_6(wires_56_5[0], addr_56_5, wires_224_6,addr_224_6);

wire[3:0] wires_225_6;

wire[31:0] addr_225_6;

Selector_2 s225_6(wires_56_5[1], addr_56_5, wires_225_6,addr_225_6);

wire[3:0] wires_226_6;

wire[31:0] addr_226_6;

Selector_2 s226_6(wires_56_5[2], addr_56_5, wires_226_6,addr_226_6);

wire[3:0] wires_227_6;

wire[31:0] addr_227_6;

Selector_2 s227_6(wires_56_5[3], addr_56_5, wires_227_6,addr_227_6);

wire[3:0] wires_228_6;

wire[31:0] addr_228_6;

Selector_2 s228_6(wires_57_5[0], addr_57_5, wires_228_6,addr_228_6);

wire[3:0] wires_229_6;

wire[31:0] addr_229_6;

Selector_2 s229_6(wires_57_5[1], addr_57_5, wires_229_6,addr_229_6);

wire[3:0] wires_230_6;

wire[31:0] addr_230_6;

Selector_2 s230_6(wires_57_5[2], addr_57_5, wires_230_6,addr_230_6);

wire[3:0] wires_231_6;

wire[31:0] addr_231_6;

Selector_2 s231_6(wires_57_5[3], addr_57_5, wires_231_6,addr_231_6);

wire[3:0] wires_232_6;

wire[31:0] addr_232_6;

Selector_2 s232_6(wires_58_5[0], addr_58_5, wires_232_6,addr_232_6);

wire[3:0] wires_233_6;

wire[31:0] addr_233_6;

Selector_2 s233_6(wires_58_5[1], addr_58_5, wires_233_6,addr_233_6);

wire[3:0] wires_234_6;

wire[31:0] addr_234_6;

Selector_2 s234_6(wires_58_5[2], addr_58_5, wires_234_6,addr_234_6);

wire[3:0] wires_235_6;

wire[31:0] addr_235_6;

Selector_2 s235_6(wires_58_5[3], addr_58_5, wires_235_6,addr_235_6);

wire[3:0] wires_236_6;

wire[31:0] addr_236_6;

Selector_2 s236_6(wires_59_5[0], addr_59_5, wires_236_6,addr_236_6);

wire[3:0] wires_237_6;

wire[31:0] addr_237_6;

Selector_2 s237_6(wires_59_5[1], addr_59_5, wires_237_6,addr_237_6);

wire[3:0] wires_238_6;

wire[31:0] addr_238_6;

Selector_2 s238_6(wires_59_5[2], addr_59_5, wires_238_6,addr_238_6);

wire[3:0] wires_239_6;

wire[31:0] addr_239_6;

Selector_2 s239_6(wires_59_5[3], addr_59_5, wires_239_6,addr_239_6);

wire[3:0] wires_240_6;

wire[31:0] addr_240_6;

Selector_2 s240_6(wires_60_5[0], addr_60_5, wires_240_6,addr_240_6);

wire[3:0] wires_241_6;

wire[31:0] addr_241_6;

Selector_2 s241_6(wires_60_5[1], addr_60_5, wires_241_6,addr_241_6);

wire[3:0] wires_242_6;

wire[31:0] addr_242_6;

Selector_2 s242_6(wires_60_5[2], addr_60_5, wires_242_6,addr_242_6);

wire[3:0] wires_243_6;

wire[31:0] addr_243_6;

Selector_2 s243_6(wires_60_5[3], addr_60_5, wires_243_6,addr_243_6);

wire[3:0] wires_244_6;

wire[31:0] addr_244_6;

Selector_2 s244_6(wires_61_5[0], addr_61_5, wires_244_6,addr_244_6);

wire[3:0] wires_245_6;

wire[31:0] addr_245_6;

Selector_2 s245_6(wires_61_5[1], addr_61_5, wires_245_6,addr_245_6);

wire[3:0] wires_246_6;

wire[31:0] addr_246_6;

Selector_2 s246_6(wires_61_5[2], addr_61_5, wires_246_6,addr_246_6);

wire[3:0] wires_247_6;

wire[31:0] addr_247_6;

Selector_2 s247_6(wires_61_5[3], addr_61_5, wires_247_6,addr_247_6);

wire[3:0] wires_248_6;

wire[31:0] addr_248_6;

Selector_2 s248_6(wires_62_5[0], addr_62_5, wires_248_6,addr_248_6);

wire[3:0] wires_249_6;

wire[31:0] addr_249_6;

Selector_2 s249_6(wires_62_5[1], addr_62_5, wires_249_6,addr_249_6);

wire[3:0] wires_250_6;

wire[31:0] addr_250_6;

Selector_2 s250_6(wires_62_5[2], addr_62_5, wires_250_6,addr_250_6);

wire[3:0] wires_251_6;

wire[31:0] addr_251_6;

Selector_2 s251_6(wires_62_5[3], addr_62_5, wires_251_6,addr_251_6);

wire[3:0] wires_252_6;

wire[31:0] addr_252_6;

Selector_2 s252_6(wires_63_5[0], addr_63_5, wires_252_6,addr_252_6);

wire[3:0] wires_253_6;

wire[31:0] addr_253_6;

Selector_2 s253_6(wires_63_5[1], addr_63_5, wires_253_6,addr_253_6);

wire[3:0] wires_254_6;

wire[31:0] addr_254_6;

Selector_2 s254_6(wires_63_5[2], addr_63_5, wires_254_6,addr_254_6);

wire[3:0] wires_255_6;

wire[31:0] addr_255_6;

Selector_2 s255_6(wires_63_5[3], addr_63_5, wires_255_6,addr_255_6);

wire[3:0] wires_256_6;

wire[31:0] addr_256_6;

Selector_2 s256_6(wires_64_5[0], addr_64_5, wires_256_6,addr_256_6);

wire[3:0] wires_257_6;

wire[31:0] addr_257_6;

Selector_2 s257_6(wires_64_5[1], addr_64_5, wires_257_6,addr_257_6);

wire[3:0] wires_258_6;

wire[31:0] addr_258_6;

Selector_2 s258_6(wires_64_5[2], addr_64_5, wires_258_6,addr_258_6);

wire[3:0] wires_259_6;

wire[31:0] addr_259_6;

Selector_2 s259_6(wires_64_5[3], addr_64_5, wires_259_6,addr_259_6);

wire[3:0] wires_260_6;

wire[31:0] addr_260_6;

Selector_2 s260_6(wires_65_5[0], addr_65_5, wires_260_6,addr_260_6);

wire[3:0] wires_261_6;

wire[31:0] addr_261_6;

Selector_2 s261_6(wires_65_5[1], addr_65_5, wires_261_6,addr_261_6);

wire[3:0] wires_262_6;

wire[31:0] addr_262_6;

Selector_2 s262_6(wires_65_5[2], addr_65_5, wires_262_6,addr_262_6);

wire[3:0] wires_263_6;

wire[31:0] addr_263_6;

Selector_2 s263_6(wires_65_5[3], addr_65_5, wires_263_6,addr_263_6);

wire[3:0] wires_264_6;

wire[31:0] addr_264_6;

Selector_2 s264_6(wires_66_5[0], addr_66_5, wires_264_6,addr_264_6);

wire[3:0] wires_265_6;

wire[31:0] addr_265_6;

Selector_2 s265_6(wires_66_5[1], addr_66_5, wires_265_6,addr_265_6);

wire[3:0] wires_266_6;

wire[31:0] addr_266_6;

Selector_2 s266_6(wires_66_5[2], addr_66_5, wires_266_6,addr_266_6);

wire[3:0] wires_267_6;

wire[31:0] addr_267_6;

Selector_2 s267_6(wires_66_5[3], addr_66_5, wires_267_6,addr_267_6);

wire[3:0] wires_268_6;

wire[31:0] addr_268_6;

Selector_2 s268_6(wires_67_5[0], addr_67_5, wires_268_6,addr_268_6);

wire[3:0] wires_269_6;

wire[31:0] addr_269_6;

Selector_2 s269_6(wires_67_5[1], addr_67_5, wires_269_6,addr_269_6);

wire[3:0] wires_270_6;

wire[31:0] addr_270_6;

Selector_2 s270_6(wires_67_5[2], addr_67_5, wires_270_6,addr_270_6);

wire[3:0] wires_271_6;

wire[31:0] addr_271_6;

Selector_2 s271_6(wires_67_5[3], addr_67_5, wires_271_6,addr_271_6);

wire[3:0] wires_272_6;

wire[31:0] addr_272_6;

Selector_2 s272_6(wires_68_5[0], addr_68_5, wires_272_6,addr_272_6);

wire[3:0] wires_273_6;

wire[31:0] addr_273_6;

Selector_2 s273_6(wires_68_5[1], addr_68_5, wires_273_6,addr_273_6);

wire[3:0] wires_274_6;

wire[31:0] addr_274_6;

Selector_2 s274_6(wires_68_5[2], addr_68_5, wires_274_6,addr_274_6);

wire[3:0] wires_275_6;

wire[31:0] addr_275_6;

Selector_2 s275_6(wires_68_5[3], addr_68_5, wires_275_6,addr_275_6);

wire[3:0] wires_276_6;

wire[31:0] addr_276_6;

Selector_2 s276_6(wires_69_5[0], addr_69_5, wires_276_6,addr_276_6);

wire[3:0] wires_277_6;

wire[31:0] addr_277_6;

Selector_2 s277_6(wires_69_5[1], addr_69_5, wires_277_6,addr_277_6);

wire[3:0] wires_278_6;

wire[31:0] addr_278_6;

Selector_2 s278_6(wires_69_5[2], addr_69_5, wires_278_6,addr_278_6);

wire[3:0] wires_279_6;

wire[31:0] addr_279_6;

Selector_2 s279_6(wires_69_5[3], addr_69_5, wires_279_6,addr_279_6);

wire[3:0] wires_280_6;

wire[31:0] addr_280_6;

Selector_2 s280_6(wires_70_5[0], addr_70_5, wires_280_6,addr_280_6);

wire[3:0] wires_281_6;

wire[31:0] addr_281_6;

Selector_2 s281_6(wires_70_5[1], addr_70_5, wires_281_6,addr_281_6);

wire[3:0] wires_282_6;

wire[31:0] addr_282_6;

Selector_2 s282_6(wires_70_5[2], addr_70_5, wires_282_6,addr_282_6);

wire[3:0] wires_283_6;

wire[31:0] addr_283_6;

Selector_2 s283_6(wires_70_5[3], addr_70_5, wires_283_6,addr_283_6);

wire[3:0] wires_284_6;

wire[31:0] addr_284_6;

Selector_2 s284_6(wires_71_5[0], addr_71_5, wires_284_6,addr_284_6);

wire[3:0] wires_285_6;

wire[31:0] addr_285_6;

Selector_2 s285_6(wires_71_5[1], addr_71_5, wires_285_6,addr_285_6);

wire[3:0] wires_286_6;

wire[31:0] addr_286_6;

Selector_2 s286_6(wires_71_5[2], addr_71_5, wires_286_6,addr_286_6);

wire[3:0] wires_287_6;

wire[31:0] addr_287_6;

Selector_2 s287_6(wires_71_5[3], addr_71_5, wires_287_6,addr_287_6);

wire[3:0] wires_288_6;

wire[31:0] addr_288_6;

Selector_2 s288_6(wires_72_5[0], addr_72_5, wires_288_6,addr_288_6);

wire[3:0] wires_289_6;

wire[31:0] addr_289_6;

Selector_2 s289_6(wires_72_5[1], addr_72_5, wires_289_6,addr_289_6);

wire[3:0] wires_290_6;

wire[31:0] addr_290_6;

Selector_2 s290_6(wires_72_5[2], addr_72_5, wires_290_6,addr_290_6);

wire[3:0] wires_291_6;

wire[31:0] addr_291_6;

Selector_2 s291_6(wires_72_5[3], addr_72_5, wires_291_6,addr_291_6);

wire[3:0] wires_292_6;

wire[31:0] addr_292_6;

Selector_2 s292_6(wires_73_5[0], addr_73_5, wires_292_6,addr_292_6);

wire[3:0] wires_293_6;

wire[31:0] addr_293_6;

Selector_2 s293_6(wires_73_5[1], addr_73_5, wires_293_6,addr_293_6);

wire[3:0] wires_294_6;

wire[31:0] addr_294_6;

Selector_2 s294_6(wires_73_5[2], addr_73_5, wires_294_6,addr_294_6);

wire[3:0] wires_295_6;

wire[31:0] addr_295_6;

Selector_2 s295_6(wires_73_5[3], addr_73_5, wires_295_6,addr_295_6);

wire[3:0] wires_296_6;

wire[31:0] addr_296_6;

Selector_2 s296_6(wires_74_5[0], addr_74_5, wires_296_6,addr_296_6);

wire[3:0] wires_297_6;

wire[31:0] addr_297_6;

Selector_2 s297_6(wires_74_5[1], addr_74_5, wires_297_6,addr_297_6);

wire[3:0] wires_298_6;

wire[31:0] addr_298_6;

Selector_2 s298_6(wires_74_5[2], addr_74_5, wires_298_6,addr_298_6);

wire[3:0] wires_299_6;

wire[31:0] addr_299_6;

Selector_2 s299_6(wires_74_5[3], addr_74_5, wires_299_6,addr_299_6);

wire[3:0] wires_300_6;

wire[31:0] addr_300_6;

Selector_2 s300_6(wires_75_5[0], addr_75_5, wires_300_6,addr_300_6);

wire[3:0] wires_301_6;

wire[31:0] addr_301_6;

Selector_2 s301_6(wires_75_5[1], addr_75_5, wires_301_6,addr_301_6);

wire[3:0] wires_302_6;

wire[31:0] addr_302_6;

Selector_2 s302_6(wires_75_5[2], addr_75_5, wires_302_6,addr_302_6);

wire[3:0] wires_303_6;

wire[31:0] addr_303_6;

Selector_2 s303_6(wires_75_5[3], addr_75_5, wires_303_6,addr_303_6);

wire[3:0] wires_304_6;

wire[31:0] addr_304_6;

Selector_2 s304_6(wires_76_5[0], addr_76_5, wires_304_6,addr_304_6);

wire[3:0] wires_305_6;

wire[31:0] addr_305_6;

Selector_2 s305_6(wires_76_5[1], addr_76_5, wires_305_6,addr_305_6);

wire[3:0] wires_306_6;

wire[31:0] addr_306_6;

Selector_2 s306_6(wires_76_5[2], addr_76_5, wires_306_6,addr_306_6);

wire[3:0] wires_307_6;

wire[31:0] addr_307_6;

Selector_2 s307_6(wires_76_5[3], addr_76_5, wires_307_6,addr_307_6);

wire[3:0] wires_308_6;

wire[31:0] addr_308_6;

Selector_2 s308_6(wires_77_5[0], addr_77_5, wires_308_6,addr_308_6);

wire[3:0] wires_309_6;

wire[31:0] addr_309_6;

Selector_2 s309_6(wires_77_5[1], addr_77_5, wires_309_6,addr_309_6);

wire[3:0] wires_310_6;

wire[31:0] addr_310_6;

Selector_2 s310_6(wires_77_5[2], addr_77_5, wires_310_6,addr_310_6);

wire[3:0] wires_311_6;

wire[31:0] addr_311_6;

Selector_2 s311_6(wires_77_5[3], addr_77_5, wires_311_6,addr_311_6);

wire[3:0] wires_312_6;

wire[31:0] addr_312_6;

Selector_2 s312_6(wires_78_5[0], addr_78_5, wires_312_6,addr_312_6);

wire[3:0] wires_313_6;

wire[31:0] addr_313_6;

Selector_2 s313_6(wires_78_5[1], addr_78_5, wires_313_6,addr_313_6);

wire[3:0] wires_314_6;

wire[31:0] addr_314_6;

Selector_2 s314_6(wires_78_5[2], addr_78_5, wires_314_6,addr_314_6);

wire[3:0] wires_315_6;

wire[31:0] addr_315_6;

Selector_2 s315_6(wires_78_5[3], addr_78_5, wires_315_6,addr_315_6);

wire[3:0] wires_316_6;

wire[31:0] addr_316_6;

Selector_2 s316_6(wires_79_5[0], addr_79_5, wires_316_6,addr_316_6);

wire[3:0] wires_317_6;

wire[31:0] addr_317_6;

Selector_2 s317_6(wires_79_5[1], addr_79_5, wires_317_6,addr_317_6);

wire[3:0] wires_318_6;

wire[31:0] addr_318_6;

Selector_2 s318_6(wires_79_5[2], addr_79_5, wires_318_6,addr_318_6);

wire[3:0] wires_319_6;

wire[31:0] addr_319_6;

Selector_2 s319_6(wires_79_5[3], addr_79_5, wires_319_6,addr_319_6);

wire[3:0] wires_320_6;

wire[31:0] addr_320_6;

Selector_2 s320_6(wires_80_5[0], addr_80_5, wires_320_6,addr_320_6);

wire[3:0] wires_321_6;

wire[31:0] addr_321_6;

Selector_2 s321_6(wires_80_5[1], addr_80_5, wires_321_6,addr_321_6);

wire[3:0] wires_322_6;

wire[31:0] addr_322_6;

Selector_2 s322_6(wires_80_5[2], addr_80_5, wires_322_6,addr_322_6);

wire[3:0] wires_323_6;

wire[31:0] addr_323_6;

Selector_2 s323_6(wires_80_5[3], addr_80_5, wires_323_6,addr_323_6);

wire[3:0] wires_324_6;

wire[31:0] addr_324_6;

Selector_2 s324_6(wires_81_5[0], addr_81_5, wires_324_6,addr_324_6);

wire[3:0] wires_325_6;

wire[31:0] addr_325_6;

Selector_2 s325_6(wires_81_5[1], addr_81_5, wires_325_6,addr_325_6);

wire[3:0] wires_326_6;

wire[31:0] addr_326_6;

Selector_2 s326_6(wires_81_5[2], addr_81_5, wires_326_6,addr_326_6);

wire[3:0] wires_327_6;

wire[31:0] addr_327_6;

Selector_2 s327_6(wires_81_5[3], addr_81_5, wires_327_6,addr_327_6);

wire[3:0] wires_328_6;

wire[31:0] addr_328_6;

Selector_2 s328_6(wires_82_5[0], addr_82_5, wires_328_6,addr_328_6);

wire[3:0] wires_329_6;

wire[31:0] addr_329_6;

Selector_2 s329_6(wires_82_5[1], addr_82_5, wires_329_6,addr_329_6);

wire[3:0] wires_330_6;

wire[31:0] addr_330_6;

Selector_2 s330_6(wires_82_5[2], addr_82_5, wires_330_6,addr_330_6);

wire[3:0] wires_331_6;

wire[31:0] addr_331_6;

Selector_2 s331_6(wires_82_5[3], addr_82_5, wires_331_6,addr_331_6);

wire[3:0] wires_332_6;

wire[31:0] addr_332_6;

Selector_2 s332_6(wires_83_5[0], addr_83_5, wires_332_6,addr_332_6);

wire[3:0] wires_333_6;

wire[31:0] addr_333_6;

Selector_2 s333_6(wires_83_5[1], addr_83_5, wires_333_6,addr_333_6);

wire[3:0] wires_334_6;

wire[31:0] addr_334_6;

Selector_2 s334_6(wires_83_5[2], addr_83_5, wires_334_6,addr_334_6);

wire[3:0] wires_335_6;

wire[31:0] addr_335_6;

Selector_2 s335_6(wires_83_5[3], addr_83_5, wires_335_6,addr_335_6);

wire[3:0] wires_336_6;

wire[31:0] addr_336_6;

Selector_2 s336_6(wires_84_5[0], addr_84_5, wires_336_6,addr_336_6);

wire[3:0] wires_337_6;

wire[31:0] addr_337_6;

Selector_2 s337_6(wires_84_5[1], addr_84_5, wires_337_6,addr_337_6);

wire[3:0] wires_338_6;

wire[31:0] addr_338_6;

Selector_2 s338_6(wires_84_5[2], addr_84_5, wires_338_6,addr_338_6);

wire[3:0] wires_339_6;

wire[31:0] addr_339_6;

Selector_2 s339_6(wires_84_5[3], addr_84_5, wires_339_6,addr_339_6);

wire[3:0] wires_340_6;

wire[31:0] addr_340_6;

Selector_2 s340_6(wires_85_5[0], addr_85_5, wires_340_6,addr_340_6);

wire[3:0] wires_341_6;

wire[31:0] addr_341_6;

Selector_2 s341_6(wires_85_5[1], addr_85_5, wires_341_6,addr_341_6);

wire[3:0] wires_342_6;

wire[31:0] addr_342_6;

Selector_2 s342_6(wires_85_5[2], addr_85_5, wires_342_6,addr_342_6);

wire[3:0] wires_343_6;

wire[31:0] addr_343_6;

Selector_2 s343_6(wires_85_5[3], addr_85_5, wires_343_6,addr_343_6);

wire[3:0] wires_344_6;

wire[31:0] addr_344_6;

Selector_2 s344_6(wires_86_5[0], addr_86_5, wires_344_6,addr_344_6);

wire[3:0] wires_345_6;

wire[31:0] addr_345_6;

Selector_2 s345_6(wires_86_5[1], addr_86_5, wires_345_6,addr_345_6);

wire[3:0] wires_346_6;

wire[31:0] addr_346_6;

Selector_2 s346_6(wires_86_5[2], addr_86_5, wires_346_6,addr_346_6);

wire[3:0] wires_347_6;

wire[31:0] addr_347_6;

Selector_2 s347_6(wires_86_5[3], addr_86_5, wires_347_6,addr_347_6);

wire[3:0] wires_348_6;

wire[31:0] addr_348_6;

Selector_2 s348_6(wires_87_5[0], addr_87_5, wires_348_6,addr_348_6);

wire[3:0] wires_349_6;

wire[31:0] addr_349_6;

Selector_2 s349_6(wires_87_5[1], addr_87_5, wires_349_6,addr_349_6);

wire[3:0] wires_350_6;

wire[31:0] addr_350_6;

Selector_2 s350_6(wires_87_5[2], addr_87_5, wires_350_6,addr_350_6);

wire[3:0] wires_351_6;

wire[31:0] addr_351_6;

Selector_2 s351_6(wires_87_5[3], addr_87_5, wires_351_6,addr_351_6);

wire[3:0] wires_352_6;

wire[31:0] addr_352_6;

Selector_2 s352_6(wires_88_5[0], addr_88_5, wires_352_6,addr_352_6);

wire[3:0] wires_353_6;

wire[31:0] addr_353_6;

Selector_2 s353_6(wires_88_5[1], addr_88_5, wires_353_6,addr_353_6);

wire[3:0] wires_354_6;

wire[31:0] addr_354_6;

Selector_2 s354_6(wires_88_5[2], addr_88_5, wires_354_6,addr_354_6);

wire[3:0] wires_355_6;

wire[31:0] addr_355_6;

Selector_2 s355_6(wires_88_5[3], addr_88_5, wires_355_6,addr_355_6);

wire[3:0] wires_356_6;

wire[31:0] addr_356_6;

Selector_2 s356_6(wires_89_5[0], addr_89_5, wires_356_6,addr_356_6);

wire[3:0] wires_357_6;

wire[31:0] addr_357_6;

Selector_2 s357_6(wires_89_5[1], addr_89_5, wires_357_6,addr_357_6);

wire[3:0] wires_358_6;

wire[31:0] addr_358_6;

Selector_2 s358_6(wires_89_5[2], addr_89_5, wires_358_6,addr_358_6);

wire[3:0] wires_359_6;

wire[31:0] addr_359_6;

Selector_2 s359_6(wires_89_5[3], addr_89_5, wires_359_6,addr_359_6);

wire[3:0] wires_360_6;

wire[31:0] addr_360_6;

Selector_2 s360_6(wires_90_5[0], addr_90_5, wires_360_6,addr_360_6);

wire[3:0] wires_361_6;

wire[31:0] addr_361_6;

Selector_2 s361_6(wires_90_5[1], addr_90_5, wires_361_6,addr_361_6);

wire[3:0] wires_362_6;

wire[31:0] addr_362_6;

Selector_2 s362_6(wires_90_5[2], addr_90_5, wires_362_6,addr_362_6);

wire[3:0] wires_363_6;

wire[31:0] addr_363_6;

Selector_2 s363_6(wires_90_5[3], addr_90_5, wires_363_6,addr_363_6);

wire[3:0] wires_364_6;

wire[31:0] addr_364_6;

Selector_2 s364_6(wires_91_5[0], addr_91_5, wires_364_6,addr_364_6);

wire[3:0] wires_365_6;

wire[31:0] addr_365_6;

Selector_2 s365_6(wires_91_5[1], addr_91_5, wires_365_6,addr_365_6);

wire[3:0] wires_366_6;

wire[31:0] addr_366_6;

Selector_2 s366_6(wires_91_5[2], addr_91_5, wires_366_6,addr_366_6);

wire[3:0] wires_367_6;

wire[31:0] addr_367_6;

Selector_2 s367_6(wires_91_5[3], addr_91_5, wires_367_6,addr_367_6);

wire[3:0] wires_368_6;

wire[31:0] addr_368_6;

Selector_2 s368_6(wires_92_5[0], addr_92_5, wires_368_6,addr_368_6);

wire[3:0] wires_369_6;

wire[31:0] addr_369_6;

Selector_2 s369_6(wires_92_5[1], addr_92_5, wires_369_6,addr_369_6);

wire[3:0] wires_370_6;

wire[31:0] addr_370_6;

Selector_2 s370_6(wires_92_5[2], addr_92_5, wires_370_6,addr_370_6);

wire[3:0] wires_371_6;

wire[31:0] addr_371_6;

Selector_2 s371_6(wires_92_5[3], addr_92_5, wires_371_6,addr_371_6);

wire[3:0] wires_372_6;

wire[31:0] addr_372_6;

Selector_2 s372_6(wires_93_5[0], addr_93_5, wires_372_6,addr_372_6);

wire[3:0] wires_373_6;

wire[31:0] addr_373_6;

Selector_2 s373_6(wires_93_5[1], addr_93_5, wires_373_6,addr_373_6);

wire[3:0] wires_374_6;

wire[31:0] addr_374_6;

Selector_2 s374_6(wires_93_5[2], addr_93_5, wires_374_6,addr_374_6);

wire[3:0] wires_375_6;

wire[31:0] addr_375_6;

Selector_2 s375_6(wires_93_5[3], addr_93_5, wires_375_6,addr_375_6);

wire[3:0] wires_376_6;

wire[31:0] addr_376_6;

Selector_2 s376_6(wires_94_5[0], addr_94_5, wires_376_6,addr_376_6);

wire[3:0] wires_377_6;

wire[31:0] addr_377_6;

Selector_2 s377_6(wires_94_5[1], addr_94_5, wires_377_6,addr_377_6);

wire[3:0] wires_378_6;

wire[31:0] addr_378_6;

Selector_2 s378_6(wires_94_5[2], addr_94_5, wires_378_6,addr_378_6);

wire[3:0] wires_379_6;

wire[31:0] addr_379_6;

Selector_2 s379_6(wires_94_5[3], addr_94_5, wires_379_6,addr_379_6);

wire[3:0] wires_380_6;

wire[31:0] addr_380_6;

Selector_2 s380_6(wires_95_5[0], addr_95_5, wires_380_6,addr_380_6);

wire[3:0] wires_381_6;

wire[31:0] addr_381_6;

Selector_2 s381_6(wires_95_5[1], addr_95_5, wires_381_6,addr_381_6);

wire[3:0] wires_382_6;

wire[31:0] addr_382_6;

Selector_2 s382_6(wires_95_5[2], addr_95_5, wires_382_6,addr_382_6);

wire[3:0] wires_383_6;

wire[31:0] addr_383_6;

Selector_2 s383_6(wires_95_5[3], addr_95_5, wires_383_6,addr_383_6);

wire[3:0] wires_384_6;

wire[31:0] addr_384_6;

Selector_2 s384_6(wires_96_5[0], addr_96_5, wires_384_6,addr_384_6);

wire[3:0] wires_385_6;

wire[31:0] addr_385_6;

Selector_2 s385_6(wires_96_5[1], addr_96_5, wires_385_6,addr_385_6);

wire[3:0] wires_386_6;

wire[31:0] addr_386_6;

Selector_2 s386_6(wires_96_5[2], addr_96_5, wires_386_6,addr_386_6);

wire[3:0] wires_387_6;

wire[31:0] addr_387_6;

Selector_2 s387_6(wires_96_5[3], addr_96_5, wires_387_6,addr_387_6);

wire[3:0] wires_388_6;

wire[31:0] addr_388_6;

Selector_2 s388_6(wires_97_5[0], addr_97_5, wires_388_6,addr_388_6);

wire[3:0] wires_389_6;

wire[31:0] addr_389_6;

Selector_2 s389_6(wires_97_5[1], addr_97_5, wires_389_6,addr_389_6);

wire[3:0] wires_390_6;

wire[31:0] addr_390_6;

Selector_2 s390_6(wires_97_5[2], addr_97_5, wires_390_6,addr_390_6);

wire[3:0] wires_391_6;

wire[31:0] addr_391_6;

Selector_2 s391_6(wires_97_5[3], addr_97_5, wires_391_6,addr_391_6);

wire[3:0] wires_392_6;

wire[31:0] addr_392_6;

Selector_2 s392_6(wires_98_5[0], addr_98_5, wires_392_6,addr_392_6);

wire[3:0] wires_393_6;

wire[31:0] addr_393_6;

Selector_2 s393_6(wires_98_5[1], addr_98_5, wires_393_6,addr_393_6);

wire[3:0] wires_394_6;

wire[31:0] addr_394_6;

Selector_2 s394_6(wires_98_5[2], addr_98_5, wires_394_6,addr_394_6);

wire[3:0] wires_395_6;

wire[31:0] addr_395_6;

Selector_2 s395_6(wires_98_5[3], addr_98_5, wires_395_6,addr_395_6);

wire[3:0] wires_396_6;

wire[31:0] addr_396_6;

Selector_2 s396_6(wires_99_5[0], addr_99_5, wires_396_6,addr_396_6);

wire[3:0] wires_397_6;

wire[31:0] addr_397_6;

Selector_2 s397_6(wires_99_5[1], addr_99_5, wires_397_6,addr_397_6);

wire[3:0] wires_398_6;

wire[31:0] addr_398_6;

Selector_2 s398_6(wires_99_5[2], addr_99_5, wires_398_6,addr_398_6);

wire[3:0] wires_399_6;

wire[31:0] addr_399_6;

Selector_2 s399_6(wires_99_5[3], addr_99_5, wires_399_6,addr_399_6);

wire[3:0] wires_400_6;

wire[31:0] addr_400_6;

Selector_2 s400_6(wires_100_5[0], addr_100_5, wires_400_6,addr_400_6);

wire[3:0] wires_401_6;

wire[31:0] addr_401_6;

Selector_2 s401_6(wires_100_5[1], addr_100_5, wires_401_6,addr_401_6);

wire[3:0] wires_402_6;

wire[31:0] addr_402_6;

Selector_2 s402_6(wires_100_5[2], addr_100_5, wires_402_6,addr_402_6);

wire[3:0] wires_403_6;

wire[31:0] addr_403_6;

Selector_2 s403_6(wires_100_5[3], addr_100_5, wires_403_6,addr_403_6);

wire[3:0] wires_404_6;

wire[31:0] addr_404_6;

Selector_2 s404_6(wires_101_5[0], addr_101_5, wires_404_6,addr_404_6);

wire[3:0] wires_405_6;

wire[31:0] addr_405_6;

Selector_2 s405_6(wires_101_5[1], addr_101_5, wires_405_6,addr_405_6);

wire[3:0] wires_406_6;

wire[31:0] addr_406_6;

Selector_2 s406_6(wires_101_5[2], addr_101_5, wires_406_6,addr_406_6);

wire[3:0] wires_407_6;

wire[31:0] addr_407_6;

Selector_2 s407_6(wires_101_5[3], addr_101_5, wires_407_6,addr_407_6);

wire[3:0] wires_408_6;

wire[31:0] addr_408_6;

Selector_2 s408_6(wires_102_5[0], addr_102_5, wires_408_6,addr_408_6);

wire[3:0] wires_409_6;

wire[31:0] addr_409_6;

Selector_2 s409_6(wires_102_5[1], addr_102_5, wires_409_6,addr_409_6);

wire[3:0] wires_410_6;

wire[31:0] addr_410_6;

Selector_2 s410_6(wires_102_5[2], addr_102_5, wires_410_6,addr_410_6);

wire[3:0] wires_411_6;

wire[31:0] addr_411_6;

Selector_2 s411_6(wires_102_5[3], addr_102_5, wires_411_6,addr_411_6);

wire[3:0] wires_412_6;

wire[31:0] addr_412_6;

Selector_2 s412_6(wires_103_5[0], addr_103_5, wires_412_6,addr_412_6);

wire[3:0] wires_413_6;

wire[31:0] addr_413_6;

Selector_2 s413_6(wires_103_5[1], addr_103_5, wires_413_6,addr_413_6);

wire[3:0] wires_414_6;

wire[31:0] addr_414_6;

Selector_2 s414_6(wires_103_5[2], addr_103_5, wires_414_6,addr_414_6);

wire[3:0] wires_415_6;

wire[31:0] addr_415_6;

Selector_2 s415_6(wires_103_5[3], addr_103_5, wires_415_6,addr_415_6);

wire[3:0] wires_416_6;

wire[31:0] addr_416_6;

Selector_2 s416_6(wires_104_5[0], addr_104_5, wires_416_6,addr_416_6);

wire[3:0] wires_417_6;

wire[31:0] addr_417_6;

Selector_2 s417_6(wires_104_5[1], addr_104_5, wires_417_6,addr_417_6);

wire[3:0] wires_418_6;

wire[31:0] addr_418_6;

Selector_2 s418_6(wires_104_5[2], addr_104_5, wires_418_6,addr_418_6);

wire[3:0] wires_419_6;

wire[31:0] addr_419_6;

Selector_2 s419_6(wires_104_5[3], addr_104_5, wires_419_6,addr_419_6);

wire[3:0] wires_420_6;

wire[31:0] addr_420_6;

Selector_2 s420_6(wires_105_5[0], addr_105_5, wires_420_6,addr_420_6);

wire[3:0] wires_421_6;

wire[31:0] addr_421_6;

Selector_2 s421_6(wires_105_5[1], addr_105_5, wires_421_6,addr_421_6);

wire[3:0] wires_422_6;

wire[31:0] addr_422_6;

Selector_2 s422_6(wires_105_5[2], addr_105_5, wires_422_6,addr_422_6);

wire[3:0] wires_423_6;

wire[31:0] addr_423_6;

Selector_2 s423_6(wires_105_5[3], addr_105_5, wires_423_6,addr_423_6);

wire[3:0] wires_424_6;

wire[31:0] addr_424_6;

Selector_2 s424_6(wires_106_5[0], addr_106_5, wires_424_6,addr_424_6);

wire[3:0] wires_425_6;

wire[31:0] addr_425_6;

Selector_2 s425_6(wires_106_5[1], addr_106_5, wires_425_6,addr_425_6);

wire[3:0] wires_426_6;

wire[31:0] addr_426_6;

Selector_2 s426_6(wires_106_5[2], addr_106_5, wires_426_6,addr_426_6);

wire[3:0] wires_427_6;

wire[31:0] addr_427_6;

Selector_2 s427_6(wires_106_5[3], addr_106_5, wires_427_6,addr_427_6);

wire[3:0] wires_428_6;

wire[31:0] addr_428_6;

Selector_2 s428_6(wires_107_5[0], addr_107_5, wires_428_6,addr_428_6);

wire[3:0] wires_429_6;

wire[31:0] addr_429_6;

Selector_2 s429_6(wires_107_5[1], addr_107_5, wires_429_6,addr_429_6);

wire[3:0] wires_430_6;

wire[31:0] addr_430_6;

Selector_2 s430_6(wires_107_5[2], addr_107_5, wires_430_6,addr_430_6);

wire[3:0] wires_431_6;

wire[31:0] addr_431_6;

Selector_2 s431_6(wires_107_5[3], addr_107_5, wires_431_6,addr_431_6);

wire[3:0] wires_432_6;

wire[31:0] addr_432_6;

Selector_2 s432_6(wires_108_5[0], addr_108_5, wires_432_6,addr_432_6);

wire[3:0] wires_433_6;

wire[31:0] addr_433_6;

Selector_2 s433_6(wires_108_5[1], addr_108_5, wires_433_6,addr_433_6);

wire[3:0] wires_434_6;

wire[31:0] addr_434_6;

Selector_2 s434_6(wires_108_5[2], addr_108_5, wires_434_6,addr_434_6);

wire[3:0] wires_435_6;

wire[31:0] addr_435_6;

Selector_2 s435_6(wires_108_5[3], addr_108_5, wires_435_6,addr_435_6);

wire[3:0] wires_436_6;

wire[31:0] addr_436_6;

Selector_2 s436_6(wires_109_5[0], addr_109_5, wires_436_6,addr_436_6);

wire[3:0] wires_437_6;

wire[31:0] addr_437_6;

Selector_2 s437_6(wires_109_5[1], addr_109_5, wires_437_6,addr_437_6);

wire[3:0] wires_438_6;

wire[31:0] addr_438_6;

Selector_2 s438_6(wires_109_5[2], addr_109_5, wires_438_6,addr_438_6);

wire[3:0] wires_439_6;

wire[31:0] addr_439_6;

Selector_2 s439_6(wires_109_5[3], addr_109_5, wires_439_6,addr_439_6);

wire[3:0] wires_440_6;

wire[31:0] addr_440_6;

Selector_2 s440_6(wires_110_5[0], addr_110_5, wires_440_6,addr_440_6);

wire[3:0] wires_441_6;

wire[31:0] addr_441_6;

Selector_2 s441_6(wires_110_5[1], addr_110_5, wires_441_6,addr_441_6);

wire[3:0] wires_442_6;

wire[31:0] addr_442_6;

Selector_2 s442_6(wires_110_5[2], addr_110_5, wires_442_6,addr_442_6);

wire[3:0] wires_443_6;

wire[31:0] addr_443_6;

Selector_2 s443_6(wires_110_5[3], addr_110_5, wires_443_6,addr_443_6);

wire[3:0] wires_444_6;

wire[31:0] addr_444_6;

Selector_2 s444_6(wires_111_5[0], addr_111_5, wires_444_6,addr_444_6);

wire[3:0] wires_445_6;

wire[31:0] addr_445_6;

Selector_2 s445_6(wires_111_5[1], addr_111_5, wires_445_6,addr_445_6);

wire[3:0] wires_446_6;

wire[31:0] addr_446_6;

Selector_2 s446_6(wires_111_5[2], addr_111_5, wires_446_6,addr_446_6);

wire[3:0] wires_447_6;

wire[31:0] addr_447_6;

Selector_2 s447_6(wires_111_5[3], addr_111_5, wires_447_6,addr_447_6);

wire[3:0] wires_448_6;

wire[31:0] addr_448_6;

Selector_2 s448_6(wires_112_5[0], addr_112_5, wires_448_6,addr_448_6);

wire[3:0] wires_449_6;

wire[31:0] addr_449_6;

Selector_2 s449_6(wires_112_5[1], addr_112_5, wires_449_6,addr_449_6);

wire[3:0] wires_450_6;

wire[31:0] addr_450_6;

Selector_2 s450_6(wires_112_5[2], addr_112_5, wires_450_6,addr_450_6);

wire[3:0] wires_451_6;

wire[31:0] addr_451_6;

Selector_2 s451_6(wires_112_5[3], addr_112_5, wires_451_6,addr_451_6);

wire[3:0] wires_452_6;

wire[31:0] addr_452_6;

Selector_2 s452_6(wires_113_5[0], addr_113_5, wires_452_6,addr_452_6);

wire[3:0] wires_453_6;

wire[31:0] addr_453_6;

Selector_2 s453_6(wires_113_5[1], addr_113_5, wires_453_6,addr_453_6);

wire[3:0] wires_454_6;

wire[31:0] addr_454_6;

Selector_2 s454_6(wires_113_5[2], addr_113_5, wires_454_6,addr_454_6);

wire[3:0] wires_455_6;

wire[31:0] addr_455_6;

Selector_2 s455_6(wires_113_5[3], addr_113_5, wires_455_6,addr_455_6);

wire[3:0] wires_456_6;

wire[31:0] addr_456_6;

Selector_2 s456_6(wires_114_5[0], addr_114_5, wires_456_6,addr_456_6);

wire[3:0] wires_457_6;

wire[31:0] addr_457_6;

Selector_2 s457_6(wires_114_5[1], addr_114_5, wires_457_6,addr_457_6);

wire[3:0] wires_458_6;

wire[31:0] addr_458_6;

Selector_2 s458_6(wires_114_5[2], addr_114_5, wires_458_6,addr_458_6);

wire[3:0] wires_459_6;

wire[31:0] addr_459_6;

Selector_2 s459_6(wires_114_5[3], addr_114_5, wires_459_6,addr_459_6);

wire[3:0] wires_460_6;

wire[31:0] addr_460_6;

Selector_2 s460_6(wires_115_5[0], addr_115_5, wires_460_6,addr_460_6);

wire[3:0] wires_461_6;

wire[31:0] addr_461_6;

Selector_2 s461_6(wires_115_5[1], addr_115_5, wires_461_6,addr_461_6);

wire[3:0] wires_462_6;

wire[31:0] addr_462_6;

Selector_2 s462_6(wires_115_5[2], addr_115_5, wires_462_6,addr_462_6);

wire[3:0] wires_463_6;

wire[31:0] addr_463_6;

Selector_2 s463_6(wires_115_5[3], addr_115_5, wires_463_6,addr_463_6);

wire[3:0] wires_464_6;

wire[31:0] addr_464_6;

Selector_2 s464_6(wires_116_5[0], addr_116_5, wires_464_6,addr_464_6);

wire[3:0] wires_465_6;

wire[31:0] addr_465_6;

Selector_2 s465_6(wires_116_5[1], addr_116_5, wires_465_6,addr_465_6);

wire[3:0] wires_466_6;

wire[31:0] addr_466_6;

Selector_2 s466_6(wires_116_5[2], addr_116_5, wires_466_6,addr_466_6);

wire[3:0] wires_467_6;

wire[31:0] addr_467_6;

Selector_2 s467_6(wires_116_5[3], addr_116_5, wires_467_6,addr_467_6);

wire[3:0] wires_468_6;

wire[31:0] addr_468_6;

Selector_2 s468_6(wires_117_5[0], addr_117_5, wires_468_6,addr_468_6);

wire[3:0] wires_469_6;

wire[31:0] addr_469_6;

Selector_2 s469_6(wires_117_5[1], addr_117_5, wires_469_6,addr_469_6);

wire[3:0] wires_470_6;

wire[31:0] addr_470_6;

Selector_2 s470_6(wires_117_5[2], addr_117_5, wires_470_6,addr_470_6);

wire[3:0] wires_471_6;

wire[31:0] addr_471_6;

Selector_2 s471_6(wires_117_5[3], addr_117_5, wires_471_6,addr_471_6);

wire[3:0] wires_472_6;

wire[31:0] addr_472_6;

Selector_2 s472_6(wires_118_5[0], addr_118_5, wires_472_6,addr_472_6);

wire[3:0] wires_473_6;

wire[31:0] addr_473_6;

Selector_2 s473_6(wires_118_5[1], addr_118_5, wires_473_6,addr_473_6);

wire[3:0] wires_474_6;

wire[31:0] addr_474_6;

Selector_2 s474_6(wires_118_5[2], addr_118_5, wires_474_6,addr_474_6);

wire[3:0] wires_475_6;

wire[31:0] addr_475_6;

Selector_2 s475_6(wires_118_5[3], addr_118_5, wires_475_6,addr_475_6);

wire[3:0] wires_476_6;

wire[31:0] addr_476_6;

Selector_2 s476_6(wires_119_5[0], addr_119_5, wires_476_6,addr_476_6);

wire[3:0] wires_477_6;

wire[31:0] addr_477_6;

Selector_2 s477_6(wires_119_5[1], addr_119_5, wires_477_6,addr_477_6);

wire[3:0] wires_478_6;

wire[31:0] addr_478_6;

Selector_2 s478_6(wires_119_5[2], addr_119_5, wires_478_6,addr_478_6);

wire[3:0] wires_479_6;

wire[31:0] addr_479_6;

Selector_2 s479_6(wires_119_5[3], addr_119_5, wires_479_6,addr_479_6);

wire[3:0] wires_480_6;

wire[31:0] addr_480_6;

Selector_2 s480_6(wires_120_5[0], addr_120_5, wires_480_6,addr_480_6);

wire[3:0] wires_481_6;

wire[31:0] addr_481_6;

Selector_2 s481_6(wires_120_5[1], addr_120_5, wires_481_6,addr_481_6);

wire[3:0] wires_482_6;

wire[31:0] addr_482_6;

Selector_2 s482_6(wires_120_5[2], addr_120_5, wires_482_6,addr_482_6);

wire[3:0] wires_483_6;

wire[31:0] addr_483_6;

Selector_2 s483_6(wires_120_5[3], addr_120_5, wires_483_6,addr_483_6);

wire[3:0] wires_484_6;

wire[31:0] addr_484_6;

Selector_2 s484_6(wires_121_5[0], addr_121_5, wires_484_6,addr_484_6);

wire[3:0] wires_485_6;

wire[31:0] addr_485_6;

Selector_2 s485_6(wires_121_5[1], addr_121_5, wires_485_6,addr_485_6);

wire[3:0] wires_486_6;

wire[31:0] addr_486_6;

Selector_2 s486_6(wires_121_5[2], addr_121_5, wires_486_6,addr_486_6);

wire[3:0] wires_487_6;

wire[31:0] addr_487_6;

Selector_2 s487_6(wires_121_5[3], addr_121_5, wires_487_6,addr_487_6);

wire[3:0] wires_488_6;

wire[31:0] addr_488_6;

Selector_2 s488_6(wires_122_5[0], addr_122_5, wires_488_6,addr_488_6);

wire[3:0] wires_489_6;

wire[31:0] addr_489_6;

Selector_2 s489_6(wires_122_5[1], addr_122_5, wires_489_6,addr_489_6);

wire[3:0] wires_490_6;

wire[31:0] addr_490_6;

Selector_2 s490_6(wires_122_5[2], addr_122_5, wires_490_6,addr_490_6);

wire[3:0] wires_491_6;

wire[31:0] addr_491_6;

Selector_2 s491_6(wires_122_5[3], addr_122_5, wires_491_6,addr_491_6);

wire[3:0] wires_492_6;

wire[31:0] addr_492_6;

Selector_2 s492_6(wires_123_5[0], addr_123_5, wires_492_6,addr_492_6);

wire[3:0] wires_493_6;

wire[31:0] addr_493_6;

Selector_2 s493_6(wires_123_5[1], addr_123_5, wires_493_6,addr_493_6);

wire[3:0] wires_494_6;

wire[31:0] addr_494_6;

Selector_2 s494_6(wires_123_5[2], addr_123_5, wires_494_6,addr_494_6);

wire[3:0] wires_495_6;

wire[31:0] addr_495_6;

Selector_2 s495_6(wires_123_5[3], addr_123_5, wires_495_6,addr_495_6);

wire[3:0] wires_496_6;

wire[31:0] addr_496_6;

Selector_2 s496_6(wires_124_5[0], addr_124_5, wires_496_6,addr_496_6);

wire[3:0] wires_497_6;

wire[31:0] addr_497_6;

Selector_2 s497_6(wires_124_5[1], addr_124_5, wires_497_6,addr_497_6);

wire[3:0] wires_498_6;

wire[31:0] addr_498_6;

Selector_2 s498_6(wires_124_5[2], addr_124_5, wires_498_6,addr_498_6);

wire[3:0] wires_499_6;

wire[31:0] addr_499_6;

Selector_2 s499_6(wires_124_5[3], addr_124_5, wires_499_6,addr_499_6);

wire[3:0] wires_500_6;

wire[31:0] addr_500_6;

Selector_2 s500_6(wires_125_5[0], addr_125_5, wires_500_6,addr_500_6);

wire[3:0] wires_501_6;

wire[31:0] addr_501_6;

Selector_2 s501_6(wires_125_5[1], addr_125_5, wires_501_6,addr_501_6);

wire[3:0] wires_502_6;

wire[31:0] addr_502_6;

Selector_2 s502_6(wires_125_5[2], addr_125_5, wires_502_6,addr_502_6);

wire[3:0] wires_503_6;

wire[31:0] addr_503_6;

Selector_2 s503_6(wires_125_5[3], addr_125_5, wires_503_6,addr_503_6);

wire[3:0] wires_504_6;

wire[31:0] addr_504_6;

Selector_2 s504_6(wires_126_5[0], addr_126_5, wires_504_6,addr_504_6);

wire[3:0] wires_505_6;

wire[31:0] addr_505_6;

Selector_2 s505_6(wires_126_5[1], addr_126_5, wires_505_6,addr_505_6);

wire[3:0] wires_506_6;

wire[31:0] addr_506_6;

Selector_2 s506_6(wires_126_5[2], addr_126_5, wires_506_6,addr_506_6);

wire[3:0] wires_507_6;

wire[31:0] addr_507_6;

Selector_2 s507_6(wires_126_5[3], addr_126_5, wires_507_6,addr_507_6);

wire[3:0] wires_508_6;

wire[31:0] addr_508_6;

Selector_2 s508_6(wires_127_5[0], addr_127_5, wires_508_6,addr_508_6);

wire[3:0] wires_509_6;

wire[31:0] addr_509_6;

Selector_2 s509_6(wires_127_5[1], addr_127_5, wires_509_6,addr_509_6);

wire[3:0] wires_510_6;

wire[31:0] addr_510_6;

Selector_2 s510_6(wires_127_5[2], addr_127_5, wires_510_6,addr_510_6);

wire[3:0] wires_511_6;

wire[31:0] addr_511_6;

Selector_2 s511_6(wires_127_5[3], addr_127_5, wires_511_6,addr_511_6);

wire[3:0] wires_512_6;

wire[31:0] addr_512_6;

Selector_2 s512_6(wires_128_5[0], addr_128_5, wires_512_6,addr_512_6);

wire[3:0] wires_513_6;

wire[31:0] addr_513_6;

Selector_2 s513_6(wires_128_5[1], addr_128_5, wires_513_6,addr_513_6);

wire[3:0] wires_514_6;

wire[31:0] addr_514_6;

Selector_2 s514_6(wires_128_5[2], addr_128_5, wires_514_6,addr_514_6);

wire[3:0] wires_515_6;

wire[31:0] addr_515_6;

Selector_2 s515_6(wires_128_5[3], addr_128_5, wires_515_6,addr_515_6);

wire[3:0] wires_516_6;

wire[31:0] addr_516_6;

Selector_2 s516_6(wires_129_5[0], addr_129_5, wires_516_6,addr_516_6);

wire[3:0] wires_517_6;

wire[31:0] addr_517_6;

Selector_2 s517_6(wires_129_5[1], addr_129_5, wires_517_6,addr_517_6);

wire[3:0] wires_518_6;

wire[31:0] addr_518_6;

Selector_2 s518_6(wires_129_5[2], addr_129_5, wires_518_6,addr_518_6);

wire[3:0] wires_519_6;

wire[31:0] addr_519_6;

Selector_2 s519_6(wires_129_5[3], addr_129_5, wires_519_6,addr_519_6);

wire[3:0] wires_520_6;

wire[31:0] addr_520_6;

Selector_2 s520_6(wires_130_5[0], addr_130_5, wires_520_6,addr_520_6);

wire[3:0] wires_521_6;

wire[31:0] addr_521_6;

Selector_2 s521_6(wires_130_5[1], addr_130_5, wires_521_6,addr_521_6);

wire[3:0] wires_522_6;

wire[31:0] addr_522_6;

Selector_2 s522_6(wires_130_5[2], addr_130_5, wires_522_6,addr_522_6);

wire[3:0] wires_523_6;

wire[31:0] addr_523_6;

Selector_2 s523_6(wires_130_5[3], addr_130_5, wires_523_6,addr_523_6);

wire[3:0] wires_524_6;

wire[31:0] addr_524_6;

Selector_2 s524_6(wires_131_5[0], addr_131_5, wires_524_6,addr_524_6);

wire[3:0] wires_525_6;

wire[31:0] addr_525_6;

Selector_2 s525_6(wires_131_5[1], addr_131_5, wires_525_6,addr_525_6);

wire[3:0] wires_526_6;

wire[31:0] addr_526_6;

Selector_2 s526_6(wires_131_5[2], addr_131_5, wires_526_6,addr_526_6);

wire[3:0] wires_527_6;

wire[31:0] addr_527_6;

Selector_2 s527_6(wires_131_5[3], addr_131_5, wires_527_6,addr_527_6);

wire[3:0] wires_528_6;

wire[31:0] addr_528_6;

Selector_2 s528_6(wires_132_5[0], addr_132_5, wires_528_6,addr_528_6);

wire[3:0] wires_529_6;

wire[31:0] addr_529_6;

Selector_2 s529_6(wires_132_5[1], addr_132_5, wires_529_6,addr_529_6);

wire[3:0] wires_530_6;

wire[31:0] addr_530_6;

Selector_2 s530_6(wires_132_5[2], addr_132_5, wires_530_6,addr_530_6);

wire[3:0] wires_531_6;

wire[31:0] addr_531_6;

Selector_2 s531_6(wires_132_5[3], addr_132_5, wires_531_6,addr_531_6);

wire[3:0] wires_532_6;

wire[31:0] addr_532_6;

Selector_2 s532_6(wires_133_5[0], addr_133_5, wires_532_6,addr_532_6);

wire[3:0] wires_533_6;

wire[31:0] addr_533_6;

Selector_2 s533_6(wires_133_5[1], addr_133_5, wires_533_6,addr_533_6);

wire[3:0] wires_534_6;

wire[31:0] addr_534_6;

Selector_2 s534_6(wires_133_5[2], addr_133_5, wires_534_6,addr_534_6);

wire[3:0] wires_535_6;

wire[31:0] addr_535_6;

Selector_2 s535_6(wires_133_5[3], addr_133_5, wires_535_6,addr_535_6);

wire[3:0] wires_536_6;

wire[31:0] addr_536_6;

Selector_2 s536_6(wires_134_5[0], addr_134_5, wires_536_6,addr_536_6);

wire[3:0] wires_537_6;

wire[31:0] addr_537_6;

Selector_2 s537_6(wires_134_5[1], addr_134_5, wires_537_6,addr_537_6);

wire[3:0] wires_538_6;

wire[31:0] addr_538_6;

Selector_2 s538_6(wires_134_5[2], addr_134_5, wires_538_6,addr_538_6);

wire[3:0] wires_539_6;

wire[31:0] addr_539_6;

Selector_2 s539_6(wires_134_5[3], addr_134_5, wires_539_6,addr_539_6);

wire[3:0] wires_540_6;

wire[31:0] addr_540_6;

Selector_2 s540_6(wires_135_5[0], addr_135_5, wires_540_6,addr_540_6);

wire[3:0] wires_541_6;

wire[31:0] addr_541_6;

Selector_2 s541_6(wires_135_5[1], addr_135_5, wires_541_6,addr_541_6);

wire[3:0] wires_542_6;

wire[31:0] addr_542_6;

Selector_2 s542_6(wires_135_5[2], addr_135_5, wires_542_6,addr_542_6);

wire[3:0] wires_543_6;

wire[31:0] addr_543_6;

Selector_2 s543_6(wires_135_5[3], addr_135_5, wires_543_6,addr_543_6);

wire[3:0] wires_544_6;

wire[31:0] addr_544_6;

Selector_2 s544_6(wires_136_5[0], addr_136_5, wires_544_6,addr_544_6);

wire[3:0] wires_545_6;

wire[31:0] addr_545_6;

Selector_2 s545_6(wires_136_5[1], addr_136_5, wires_545_6,addr_545_6);

wire[3:0] wires_546_6;

wire[31:0] addr_546_6;

Selector_2 s546_6(wires_136_5[2], addr_136_5, wires_546_6,addr_546_6);

wire[3:0] wires_547_6;

wire[31:0] addr_547_6;

Selector_2 s547_6(wires_136_5[3], addr_136_5, wires_547_6,addr_547_6);

wire[3:0] wires_548_6;

wire[31:0] addr_548_6;

Selector_2 s548_6(wires_137_5[0], addr_137_5, wires_548_6,addr_548_6);

wire[3:0] wires_549_6;

wire[31:0] addr_549_6;

Selector_2 s549_6(wires_137_5[1], addr_137_5, wires_549_6,addr_549_6);

wire[3:0] wires_550_6;

wire[31:0] addr_550_6;

Selector_2 s550_6(wires_137_5[2], addr_137_5, wires_550_6,addr_550_6);

wire[3:0] wires_551_6;

wire[31:0] addr_551_6;

Selector_2 s551_6(wires_137_5[3], addr_137_5, wires_551_6,addr_551_6);

wire[3:0] wires_552_6;

wire[31:0] addr_552_6;

Selector_2 s552_6(wires_138_5[0], addr_138_5, wires_552_6,addr_552_6);

wire[3:0] wires_553_6;

wire[31:0] addr_553_6;

Selector_2 s553_6(wires_138_5[1], addr_138_5, wires_553_6,addr_553_6);

wire[3:0] wires_554_6;

wire[31:0] addr_554_6;

Selector_2 s554_6(wires_138_5[2], addr_138_5, wires_554_6,addr_554_6);

wire[3:0] wires_555_6;

wire[31:0] addr_555_6;

Selector_2 s555_6(wires_138_5[3], addr_138_5, wires_555_6,addr_555_6);

wire[3:0] wires_556_6;

wire[31:0] addr_556_6;

Selector_2 s556_6(wires_139_5[0], addr_139_5, wires_556_6,addr_556_6);

wire[3:0] wires_557_6;

wire[31:0] addr_557_6;

Selector_2 s557_6(wires_139_5[1], addr_139_5, wires_557_6,addr_557_6);

wire[3:0] wires_558_6;

wire[31:0] addr_558_6;

Selector_2 s558_6(wires_139_5[2], addr_139_5, wires_558_6,addr_558_6);

wire[3:0] wires_559_6;

wire[31:0] addr_559_6;

Selector_2 s559_6(wires_139_5[3], addr_139_5, wires_559_6,addr_559_6);

wire[3:0] wires_560_6;

wire[31:0] addr_560_6;

Selector_2 s560_6(wires_140_5[0], addr_140_5, wires_560_6,addr_560_6);

wire[3:0] wires_561_6;

wire[31:0] addr_561_6;

Selector_2 s561_6(wires_140_5[1], addr_140_5, wires_561_6,addr_561_6);

wire[3:0] wires_562_6;

wire[31:0] addr_562_6;

Selector_2 s562_6(wires_140_5[2], addr_140_5, wires_562_6,addr_562_6);

wire[3:0] wires_563_6;

wire[31:0] addr_563_6;

Selector_2 s563_6(wires_140_5[3], addr_140_5, wires_563_6,addr_563_6);

wire[3:0] wires_564_6;

wire[31:0] addr_564_6;

Selector_2 s564_6(wires_141_5[0], addr_141_5, wires_564_6,addr_564_6);

wire[3:0] wires_565_6;

wire[31:0] addr_565_6;

Selector_2 s565_6(wires_141_5[1], addr_141_5, wires_565_6,addr_565_6);

wire[3:0] wires_566_6;

wire[31:0] addr_566_6;

Selector_2 s566_6(wires_141_5[2], addr_141_5, wires_566_6,addr_566_6);

wire[3:0] wires_567_6;

wire[31:0] addr_567_6;

Selector_2 s567_6(wires_141_5[3], addr_141_5, wires_567_6,addr_567_6);

wire[3:0] wires_568_6;

wire[31:0] addr_568_6;

Selector_2 s568_6(wires_142_5[0], addr_142_5, wires_568_6,addr_568_6);

wire[3:0] wires_569_6;

wire[31:0] addr_569_6;

Selector_2 s569_6(wires_142_5[1], addr_142_5, wires_569_6,addr_569_6);

wire[3:0] wires_570_6;

wire[31:0] addr_570_6;

Selector_2 s570_6(wires_142_5[2], addr_142_5, wires_570_6,addr_570_6);

wire[3:0] wires_571_6;

wire[31:0] addr_571_6;

Selector_2 s571_6(wires_142_5[3], addr_142_5, wires_571_6,addr_571_6);

wire[3:0] wires_572_6;

wire[31:0] addr_572_6;

Selector_2 s572_6(wires_143_5[0], addr_143_5, wires_572_6,addr_572_6);

wire[3:0] wires_573_6;

wire[31:0] addr_573_6;

Selector_2 s573_6(wires_143_5[1], addr_143_5, wires_573_6,addr_573_6);

wire[3:0] wires_574_6;

wire[31:0] addr_574_6;

Selector_2 s574_6(wires_143_5[2], addr_143_5, wires_574_6,addr_574_6);

wire[3:0] wires_575_6;

wire[31:0] addr_575_6;

Selector_2 s575_6(wires_143_5[3], addr_143_5, wires_575_6,addr_575_6);

wire[3:0] wires_576_6;

wire[31:0] addr_576_6;

Selector_2 s576_6(wires_144_5[0], addr_144_5, wires_576_6,addr_576_6);

wire[3:0] wires_577_6;

wire[31:0] addr_577_6;

Selector_2 s577_6(wires_144_5[1], addr_144_5, wires_577_6,addr_577_6);

wire[3:0] wires_578_6;

wire[31:0] addr_578_6;

Selector_2 s578_6(wires_144_5[2], addr_144_5, wires_578_6,addr_578_6);

wire[3:0] wires_579_6;

wire[31:0] addr_579_6;

Selector_2 s579_6(wires_144_5[3], addr_144_5, wires_579_6,addr_579_6);

wire[3:0] wires_580_6;

wire[31:0] addr_580_6;

Selector_2 s580_6(wires_145_5[0], addr_145_5, wires_580_6,addr_580_6);

wire[3:0] wires_581_6;

wire[31:0] addr_581_6;

Selector_2 s581_6(wires_145_5[1], addr_145_5, wires_581_6,addr_581_6);

wire[3:0] wires_582_6;

wire[31:0] addr_582_6;

Selector_2 s582_6(wires_145_5[2], addr_145_5, wires_582_6,addr_582_6);

wire[3:0] wires_583_6;

wire[31:0] addr_583_6;

Selector_2 s583_6(wires_145_5[3], addr_145_5, wires_583_6,addr_583_6);

wire[3:0] wires_584_6;

wire[31:0] addr_584_6;

Selector_2 s584_6(wires_146_5[0], addr_146_5, wires_584_6,addr_584_6);

wire[3:0] wires_585_6;

wire[31:0] addr_585_6;

Selector_2 s585_6(wires_146_5[1], addr_146_5, wires_585_6,addr_585_6);

wire[3:0] wires_586_6;

wire[31:0] addr_586_6;

Selector_2 s586_6(wires_146_5[2], addr_146_5, wires_586_6,addr_586_6);

wire[3:0] wires_587_6;

wire[31:0] addr_587_6;

Selector_2 s587_6(wires_146_5[3], addr_146_5, wires_587_6,addr_587_6);

wire[3:0] wires_588_6;

wire[31:0] addr_588_6;

Selector_2 s588_6(wires_147_5[0], addr_147_5, wires_588_6,addr_588_6);

wire[3:0] wires_589_6;

wire[31:0] addr_589_6;

Selector_2 s589_6(wires_147_5[1], addr_147_5, wires_589_6,addr_589_6);

wire[3:0] wires_590_6;

wire[31:0] addr_590_6;

Selector_2 s590_6(wires_147_5[2], addr_147_5, wires_590_6,addr_590_6);

wire[3:0] wires_591_6;

wire[31:0] addr_591_6;

Selector_2 s591_6(wires_147_5[3], addr_147_5, wires_591_6,addr_591_6);

wire[3:0] wires_592_6;

wire[31:0] addr_592_6;

Selector_2 s592_6(wires_148_5[0], addr_148_5, wires_592_6,addr_592_6);

wire[3:0] wires_593_6;

wire[31:0] addr_593_6;

Selector_2 s593_6(wires_148_5[1], addr_148_5, wires_593_6,addr_593_6);

wire[3:0] wires_594_6;

wire[31:0] addr_594_6;

Selector_2 s594_6(wires_148_5[2], addr_148_5, wires_594_6,addr_594_6);

wire[3:0] wires_595_6;

wire[31:0] addr_595_6;

Selector_2 s595_6(wires_148_5[3], addr_148_5, wires_595_6,addr_595_6);

wire[3:0] wires_596_6;

wire[31:0] addr_596_6;

Selector_2 s596_6(wires_149_5[0], addr_149_5, wires_596_6,addr_596_6);

wire[3:0] wires_597_6;

wire[31:0] addr_597_6;

Selector_2 s597_6(wires_149_5[1], addr_149_5, wires_597_6,addr_597_6);

wire[3:0] wires_598_6;

wire[31:0] addr_598_6;

Selector_2 s598_6(wires_149_5[2], addr_149_5, wires_598_6,addr_598_6);

wire[3:0] wires_599_6;

wire[31:0] addr_599_6;

Selector_2 s599_6(wires_149_5[3], addr_149_5, wires_599_6,addr_599_6);

wire[3:0] wires_600_6;

wire[31:0] addr_600_6;

Selector_2 s600_6(wires_150_5[0], addr_150_5, wires_600_6,addr_600_6);

wire[3:0] wires_601_6;

wire[31:0] addr_601_6;

Selector_2 s601_6(wires_150_5[1], addr_150_5, wires_601_6,addr_601_6);

wire[3:0] wires_602_6;

wire[31:0] addr_602_6;

Selector_2 s602_6(wires_150_5[2], addr_150_5, wires_602_6,addr_602_6);

wire[3:0] wires_603_6;

wire[31:0] addr_603_6;

Selector_2 s603_6(wires_150_5[3], addr_150_5, wires_603_6,addr_603_6);

wire[3:0] wires_604_6;

wire[31:0] addr_604_6;

Selector_2 s604_6(wires_151_5[0], addr_151_5, wires_604_6,addr_604_6);

wire[3:0] wires_605_6;

wire[31:0] addr_605_6;

Selector_2 s605_6(wires_151_5[1], addr_151_5, wires_605_6,addr_605_6);

wire[3:0] wires_606_6;

wire[31:0] addr_606_6;

Selector_2 s606_6(wires_151_5[2], addr_151_5, wires_606_6,addr_606_6);

wire[3:0] wires_607_6;

wire[31:0] addr_607_6;

Selector_2 s607_6(wires_151_5[3], addr_151_5, wires_607_6,addr_607_6);

wire[3:0] wires_608_6;

wire[31:0] addr_608_6;

Selector_2 s608_6(wires_152_5[0], addr_152_5, wires_608_6,addr_608_6);

wire[3:0] wires_609_6;

wire[31:0] addr_609_6;

Selector_2 s609_6(wires_152_5[1], addr_152_5, wires_609_6,addr_609_6);

wire[3:0] wires_610_6;

wire[31:0] addr_610_6;

Selector_2 s610_6(wires_152_5[2], addr_152_5, wires_610_6,addr_610_6);

wire[3:0] wires_611_6;

wire[31:0] addr_611_6;

Selector_2 s611_6(wires_152_5[3], addr_152_5, wires_611_6,addr_611_6);

wire[3:0] wires_612_6;

wire[31:0] addr_612_6;

Selector_2 s612_6(wires_153_5[0], addr_153_5, wires_612_6,addr_612_6);

wire[3:0] wires_613_6;

wire[31:0] addr_613_6;

Selector_2 s613_6(wires_153_5[1], addr_153_5, wires_613_6,addr_613_6);

wire[3:0] wires_614_6;

wire[31:0] addr_614_6;

Selector_2 s614_6(wires_153_5[2], addr_153_5, wires_614_6,addr_614_6);

wire[3:0] wires_615_6;

wire[31:0] addr_615_6;

Selector_2 s615_6(wires_153_5[3], addr_153_5, wires_615_6,addr_615_6);

wire[3:0] wires_616_6;

wire[31:0] addr_616_6;

Selector_2 s616_6(wires_154_5[0], addr_154_5, wires_616_6,addr_616_6);

wire[3:0] wires_617_6;

wire[31:0] addr_617_6;

Selector_2 s617_6(wires_154_5[1], addr_154_5, wires_617_6,addr_617_6);

wire[3:0] wires_618_6;

wire[31:0] addr_618_6;

Selector_2 s618_6(wires_154_5[2], addr_154_5, wires_618_6,addr_618_6);

wire[3:0] wires_619_6;

wire[31:0] addr_619_6;

Selector_2 s619_6(wires_154_5[3], addr_154_5, wires_619_6,addr_619_6);

wire[3:0] wires_620_6;

wire[31:0] addr_620_6;

Selector_2 s620_6(wires_155_5[0], addr_155_5, wires_620_6,addr_620_6);

wire[3:0] wires_621_6;

wire[31:0] addr_621_6;

Selector_2 s621_6(wires_155_5[1], addr_155_5, wires_621_6,addr_621_6);

wire[3:0] wires_622_6;

wire[31:0] addr_622_6;

Selector_2 s622_6(wires_155_5[2], addr_155_5, wires_622_6,addr_622_6);

wire[3:0] wires_623_6;

wire[31:0] addr_623_6;

Selector_2 s623_6(wires_155_5[3], addr_155_5, wires_623_6,addr_623_6);

wire[3:0] wires_624_6;

wire[31:0] addr_624_6;

Selector_2 s624_6(wires_156_5[0], addr_156_5, wires_624_6,addr_624_6);

wire[3:0] wires_625_6;

wire[31:0] addr_625_6;

Selector_2 s625_6(wires_156_5[1], addr_156_5, wires_625_6,addr_625_6);

wire[3:0] wires_626_6;

wire[31:0] addr_626_6;

Selector_2 s626_6(wires_156_5[2], addr_156_5, wires_626_6,addr_626_6);

wire[3:0] wires_627_6;

wire[31:0] addr_627_6;

Selector_2 s627_6(wires_156_5[3], addr_156_5, wires_627_6,addr_627_6);

wire[3:0] wires_628_6;

wire[31:0] addr_628_6;

Selector_2 s628_6(wires_157_5[0], addr_157_5, wires_628_6,addr_628_6);

wire[3:0] wires_629_6;

wire[31:0] addr_629_6;

Selector_2 s629_6(wires_157_5[1], addr_157_5, wires_629_6,addr_629_6);

wire[3:0] wires_630_6;

wire[31:0] addr_630_6;

Selector_2 s630_6(wires_157_5[2], addr_157_5, wires_630_6,addr_630_6);

wire[3:0] wires_631_6;

wire[31:0] addr_631_6;

Selector_2 s631_6(wires_157_5[3], addr_157_5, wires_631_6,addr_631_6);

wire[3:0] wires_632_6;

wire[31:0] addr_632_6;

Selector_2 s632_6(wires_158_5[0], addr_158_5, wires_632_6,addr_632_6);

wire[3:0] wires_633_6;

wire[31:0] addr_633_6;

Selector_2 s633_6(wires_158_5[1], addr_158_5, wires_633_6,addr_633_6);

wire[3:0] wires_634_6;

wire[31:0] addr_634_6;

Selector_2 s634_6(wires_158_5[2], addr_158_5, wires_634_6,addr_634_6);

wire[3:0] wires_635_6;

wire[31:0] addr_635_6;

Selector_2 s635_6(wires_158_5[3], addr_158_5, wires_635_6,addr_635_6);

wire[3:0] wires_636_6;

wire[31:0] addr_636_6;

Selector_2 s636_6(wires_159_5[0], addr_159_5, wires_636_6,addr_636_6);

wire[3:0] wires_637_6;

wire[31:0] addr_637_6;

Selector_2 s637_6(wires_159_5[1], addr_159_5, wires_637_6,addr_637_6);

wire[3:0] wires_638_6;

wire[31:0] addr_638_6;

Selector_2 s638_6(wires_159_5[2], addr_159_5, wires_638_6,addr_638_6);

wire[3:0] wires_639_6;

wire[31:0] addr_639_6;

Selector_2 s639_6(wires_159_5[3], addr_159_5, wires_639_6,addr_639_6);

wire[3:0] wires_640_6;

wire[31:0] addr_640_6;

Selector_2 s640_6(wires_160_5[0], addr_160_5, wires_640_6,addr_640_6);

wire[3:0] wires_641_6;

wire[31:0] addr_641_6;

Selector_2 s641_6(wires_160_5[1], addr_160_5, wires_641_6,addr_641_6);

wire[3:0] wires_642_6;

wire[31:0] addr_642_6;

Selector_2 s642_6(wires_160_5[2], addr_160_5, wires_642_6,addr_642_6);

wire[3:0] wires_643_6;

wire[31:0] addr_643_6;

Selector_2 s643_6(wires_160_5[3], addr_160_5, wires_643_6,addr_643_6);

wire[3:0] wires_644_6;

wire[31:0] addr_644_6;

Selector_2 s644_6(wires_161_5[0], addr_161_5, wires_644_6,addr_644_6);

wire[3:0] wires_645_6;

wire[31:0] addr_645_6;

Selector_2 s645_6(wires_161_5[1], addr_161_5, wires_645_6,addr_645_6);

wire[3:0] wires_646_6;

wire[31:0] addr_646_6;

Selector_2 s646_6(wires_161_5[2], addr_161_5, wires_646_6,addr_646_6);

wire[3:0] wires_647_6;

wire[31:0] addr_647_6;

Selector_2 s647_6(wires_161_5[3], addr_161_5, wires_647_6,addr_647_6);

wire[3:0] wires_648_6;

wire[31:0] addr_648_6;

Selector_2 s648_6(wires_162_5[0], addr_162_5, wires_648_6,addr_648_6);

wire[3:0] wires_649_6;

wire[31:0] addr_649_6;

Selector_2 s649_6(wires_162_5[1], addr_162_5, wires_649_6,addr_649_6);

wire[3:0] wires_650_6;

wire[31:0] addr_650_6;

Selector_2 s650_6(wires_162_5[2], addr_162_5, wires_650_6,addr_650_6);

wire[3:0] wires_651_6;

wire[31:0] addr_651_6;

Selector_2 s651_6(wires_162_5[3], addr_162_5, wires_651_6,addr_651_6);

wire[3:0] wires_652_6;

wire[31:0] addr_652_6;

Selector_2 s652_6(wires_163_5[0], addr_163_5, wires_652_6,addr_652_6);

wire[3:0] wires_653_6;

wire[31:0] addr_653_6;

Selector_2 s653_6(wires_163_5[1], addr_163_5, wires_653_6,addr_653_6);

wire[3:0] wires_654_6;

wire[31:0] addr_654_6;

Selector_2 s654_6(wires_163_5[2], addr_163_5, wires_654_6,addr_654_6);

wire[3:0] wires_655_6;

wire[31:0] addr_655_6;

Selector_2 s655_6(wires_163_5[3], addr_163_5, wires_655_6,addr_655_6);

wire[3:0] wires_656_6;

wire[31:0] addr_656_6;

Selector_2 s656_6(wires_164_5[0], addr_164_5, wires_656_6,addr_656_6);

wire[3:0] wires_657_6;

wire[31:0] addr_657_6;

Selector_2 s657_6(wires_164_5[1], addr_164_5, wires_657_6,addr_657_6);

wire[3:0] wires_658_6;

wire[31:0] addr_658_6;

Selector_2 s658_6(wires_164_5[2], addr_164_5, wires_658_6,addr_658_6);

wire[3:0] wires_659_6;

wire[31:0] addr_659_6;

Selector_2 s659_6(wires_164_5[3], addr_164_5, wires_659_6,addr_659_6);

wire[3:0] wires_660_6;

wire[31:0] addr_660_6;

Selector_2 s660_6(wires_165_5[0], addr_165_5, wires_660_6,addr_660_6);

wire[3:0] wires_661_6;

wire[31:0] addr_661_6;

Selector_2 s661_6(wires_165_5[1], addr_165_5, wires_661_6,addr_661_6);

wire[3:0] wires_662_6;

wire[31:0] addr_662_6;

Selector_2 s662_6(wires_165_5[2], addr_165_5, wires_662_6,addr_662_6);

wire[3:0] wires_663_6;

wire[31:0] addr_663_6;

Selector_2 s663_6(wires_165_5[3], addr_165_5, wires_663_6,addr_663_6);

wire[3:0] wires_664_6;

wire[31:0] addr_664_6;

Selector_2 s664_6(wires_166_5[0], addr_166_5, wires_664_6,addr_664_6);

wire[3:0] wires_665_6;

wire[31:0] addr_665_6;

Selector_2 s665_6(wires_166_5[1], addr_166_5, wires_665_6,addr_665_6);

wire[3:0] wires_666_6;

wire[31:0] addr_666_6;

Selector_2 s666_6(wires_166_5[2], addr_166_5, wires_666_6,addr_666_6);

wire[3:0] wires_667_6;

wire[31:0] addr_667_6;

Selector_2 s667_6(wires_166_5[3], addr_166_5, wires_667_6,addr_667_6);

wire[3:0] wires_668_6;

wire[31:0] addr_668_6;

Selector_2 s668_6(wires_167_5[0], addr_167_5, wires_668_6,addr_668_6);

wire[3:0] wires_669_6;

wire[31:0] addr_669_6;

Selector_2 s669_6(wires_167_5[1], addr_167_5, wires_669_6,addr_669_6);

wire[3:0] wires_670_6;

wire[31:0] addr_670_6;

Selector_2 s670_6(wires_167_5[2], addr_167_5, wires_670_6,addr_670_6);

wire[3:0] wires_671_6;

wire[31:0] addr_671_6;

Selector_2 s671_6(wires_167_5[3], addr_167_5, wires_671_6,addr_671_6);

wire[3:0] wires_672_6;

wire[31:0] addr_672_6;

Selector_2 s672_6(wires_168_5[0], addr_168_5, wires_672_6,addr_672_6);

wire[3:0] wires_673_6;

wire[31:0] addr_673_6;

Selector_2 s673_6(wires_168_5[1], addr_168_5, wires_673_6,addr_673_6);

wire[3:0] wires_674_6;

wire[31:0] addr_674_6;

Selector_2 s674_6(wires_168_5[2], addr_168_5, wires_674_6,addr_674_6);

wire[3:0] wires_675_6;

wire[31:0] addr_675_6;

Selector_2 s675_6(wires_168_5[3], addr_168_5, wires_675_6,addr_675_6);

wire[3:0] wires_676_6;

wire[31:0] addr_676_6;

Selector_2 s676_6(wires_169_5[0], addr_169_5, wires_676_6,addr_676_6);

wire[3:0] wires_677_6;

wire[31:0] addr_677_6;

Selector_2 s677_6(wires_169_5[1], addr_169_5, wires_677_6,addr_677_6);

wire[3:0] wires_678_6;

wire[31:0] addr_678_6;

Selector_2 s678_6(wires_169_5[2], addr_169_5, wires_678_6,addr_678_6);

wire[3:0] wires_679_6;

wire[31:0] addr_679_6;

Selector_2 s679_6(wires_169_5[3], addr_169_5, wires_679_6,addr_679_6);

wire[3:0] wires_680_6;

wire[31:0] addr_680_6;

Selector_2 s680_6(wires_170_5[0], addr_170_5, wires_680_6,addr_680_6);

wire[3:0] wires_681_6;

wire[31:0] addr_681_6;

Selector_2 s681_6(wires_170_5[1], addr_170_5, wires_681_6,addr_681_6);

wire[3:0] wires_682_6;

wire[31:0] addr_682_6;

Selector_2 s682_6(wires_170_5[2], addr_170_5, wires_682_6,addr_682_6);

wire[3:0] wires_683_6;

wire[31:0] addr_683_6;

Selector_2 s683_6(wires_170_5[3], addr_170_5, wires_683_6,addr_683_6);

wire[3:0] wires_684_6;

wire[31:0] addr_684_6;

Selector_2 s684_6(wires_171_5[0], addr_171_5, wires_684_6,addr_684_6);

wire[3:0] wires_685_6;

wire[31:0] addr_685_6;

Selector_2 s685_6(wires_171_5[1], addr_171_5, wires_685_6,addr_685_6);

wire[3:0] wires_686_6;

wire[31:0] addr_686_6;

Selector_2 s686_6(wires_171_5[2], addr_171_5, wires_686_6,addr_686_6);

wire[3:0] wires_687_6;

wire[31:0] addr_687_6;

Selector_2 s687_6(wires_171_5[3], addr_171_5, wires_687_6,addr_687_6);

wire[3:0] wires_688_6;

wire[31:0] addr_688_6;

Selector_2 s688_6(wires_172_5[0], addr_172_5, wires_688_6,addr_688_6);

wire[3:0] wires_689_6;

wire[31:0] addr_689_6;

Selector_2 s689_6(wires_172_5[1], addr_172_5, wires_689_6,addr_689_6);

wire[3:0] wires_690_6;

wire[31:0] addr_690_6;

Selector_2 s690_6(wires_172_5[2], addr_172_5, wires_690_6,addr_690_6);

wire[3:0] wires_691_6;

wire[31:0] addr_691_6;

Selector_2 s691_6(wires_172_5[3], addr_172_5, wires_691_6,addr_691_6);

wire[3:0] wires_692_6;

wire[31:0] addr_692_6;

Selector_2 s692_6(wires_173_5[0], addr_173_5, wires_692_6,addr_692_6);

wire[3:0] wires_693_6;

wire[31:0] addr_693_6;

Selector_2 s693_6(wires_173_5[1], addr_173_5, wires_693_6,addr_693_6);

wire[3:0] wires_694_6;

wire[31:0] addr_694_6;

Selector_2 s694_6(wires_173_5[2], addr_173_5, wires_694_6,addr_694_6);

wire[3:0] wires_695_6;

wire[31:0] addr_695_6;

Selector_2 s695_6(wires_173_5[3], addr_173_5, wires_695_6,addr_695_6);

wire[3:0] wires_696_6;

wire[31:0] addr_696_6;

Selector_2 s696_6(wires_174_5[0], addr_174_5, wires_696_6,addr_696_6);

wire[3:0] wires_697_6;

wire[31:0] addr_697_6;

Selector_2 s697_6(wires_174_5[1], addr_174_5, wires_697_6,addr_697_6);

wire[3:0] wires_698_6;

wire[31:0] addr_698_6;

Selector_2 s698_6(wires_174_5[2], addr_174_5, wires_698_6,addr_698_6);

wire[3:0] wires_699_6;

wire[31:0] addr_699_6;

Selector_2 s699_6(wires_174_5[3], addr_174_5, wires_699_6,addr_699_6);

wire[3:0] wires_700_6;

wire[31:0] addr_700_6;

Selector_2 s700_6(wires_175_5[0], addr_175_5, wires_700_6,addr_700_6);

wire[3:0] wires_701_6;

wire[31:0] addr_701_6;

Selector_2 s701_6(wires_175_5[1], addr_175_5, wires_701_6,addr_701_6);

wire[3:0] wires_702_6;

wire[31:0] addr_702_6;

Selector_2 s702_6(wires_175_5[2], addr_175_5, wires_702_6,addr_702_6);

wire[3:0] wires_703_6;

wire[31:0] addr_703_6;

Selector_2 s703_6(wires_175_5[3], addr_175_5, wires_703_6,addr_703_6);

wire[3:0] wires_704_6;

wire[31:0] addr_704_6;

Selector_2 s704_6(wires_176_5[0], addr_176_5, wires_704_6,addr_704_6);

wire[3:0] wires_705_6;

wire[31:0] addr_705_6;

Selector_2 s705_6(wires_176_5[1], addr_176_5, wires_705_6,addr_705_6);

wire[3:0] wires_706_6;

wire[31:0] addr_706_6;

Selector_2 s706_6(wires_176_5[2], addr_176_5, wires_706_6,addr_706_6);

wire[3:0] wires_707_6;

wire[31:0] addr_707_6;

Selector_2 s707_6(wires_176_5[3], addr_176_5, wires_707_6,addr_707_6);

wire[3:0] wires_708_6;

wire[31:0] addr_708_6;

Selector_2 s708_6(wires_177_5[0], addr_177_5, wires_708_6,addr_708_6);

wire[3:0] wires_709_6;

wire[31:0] addr_709_6;

Selector_2 s709_6(wires_177_5[1], addr_177_5, wires_709_6,addr_709_6);

wire[3:0] wires_710_6;

wire[31:0] addr_710_6;

Selector_2 s710_6(wires_177_5[2], addr_177_5, wires_710_6,addr_710_6);

wire[3:0] wires_711_6;

wire[31:0] addr_711_6;

Selector_2 s711_6(wires_177_5[3], addr_177_5, wires_711_6,addr_711_6);

wire[3:0] wires_712_6;

wire[31:0] addr_712_6;

Selector_2 s712_6(wires_178_5[0], addr_178_5, wires_712_6,addr_712_6);

wire[3:0] wires_713_6;

wire[31:0] addr_713_6;

Selector_2 s713_6(wires_178_5[1], addr_178_5, wires_713_6,addr_713_6);

wire[3:0] wires_714_6;

wire[31:0] addr_714_6;

Selector_2 s714_6(wires_178_5[2], addr_178_5, wires_714_6,addr_714_6);

wire[3:0] wires_715_6;

wire[31:0] addr_715_6;

Selector_2 s715_6(wires_178_5[3], addr_178_5, wires_715_6,addr_715_6);

wire[3:0] wires_716_6;

wire[31:0] addr_716_6;

Selector_2 s716_6(wires_179_5[0], addr_179_5, wires_716_6,addr_716_6);

wire[3:0] wires_717_6;

wire[31:0] addr_717_6;

Selector_2 s717_6(wires_179_5[1], addr_179_5, wires_717_6,addr_717_6);

wire[3:0] wires_718_6;

wire[31:0] addr_718_6;

Selector_2 s718_6(wires_179_5[2], addr_179_5, wires_718_6,addr_718_6);

wire[3:0] wires_719_6;

wire[31:0] addr_719_6;

Selector_2 s719_6(wires_179_5[3], addr_179_5, wires_719_6,addr_719_6);

wire[3:0] wires_720_6;

wire[31:0] addr_720_6;

Selector_2 s720_6(wires_180_5[0], addr_180_5, wires_720_6,addr_720_6);

wire[3:0] wires_721_6;

wire[31:0] addr_721_6;

Selector_2 s721_6(wires_180_5[1], addr_180_5, wires_721_6,addr_721_6);

wire[3:0] wires_722_6;

wire[31:0] addr_722_6;

Selector_2 s722_6(wires_180_5[2], addr_180_5, wires_722_6,addr_722_6);

wire[3:0] wires_723_6;

wire[31:0] addr_723_6;

Selector_2 s723_6(wires_180_5[3], addr_180_5, wires_723_6,addr_723_6);

wire[3:0] wires_724_6;

wire[31:0] addr_724_6;

Selector_2 s724_6(wires_181_5[0], addr_181_5, wires_724_6,addr_724_6);

wire[3:0] wires_725_6;

wire[31:0] addr_725_6;

Selector_2 s725_6(wires_181_5[1], addr_181_5, wires_725_6,addr_725_6);

wire[3:0] wires_726_6;

wire[31:0] addr_726_6;

Selector_2 s726_6(wires_181_5[2], addr_181_5, wires_726_6,addr_726_6);

wire[3:0] wires_727_6;

wire[31:0] addr_727_6;

Selector_2 s727_6(wires_181_5[3], addr_181_5, wires_727_6,addr_727_6);

wire[3:0] wires_728_6;

wire[31:0] addr_728_6;

Selector_2 s728_6(wires_182_5[0], addr_182_5, wires_728_6,addr_728_6);

wire[3:0] wires_729_6;

wire[31:0] addr_729_6;

Selector_2 s729_6(wires_182_5[1], addr_182_5, wires_729_6,addr_729_6);

wire[3:0] wires_730_6;

wire[31:0] addr_730_6;

Selector_2 s730_6(wires_182_5[2], addr_182_5, wires_730_6,addr_730_6);

wire[3:0] wires_731_6;

wire[31:0] addr_731_6;

Selector_2 s731_6(wires_182_5[3], addr_182_5, wires_731_6,addr_731_6);

wire[3:0] wires_732_6;

wire[31:0] addr_732_6;

Selector_2 s732_6(wires_183_5[0], addr_183_5, wires_732_6,addr_732_6);

wire[3:0] wires_733_6;

wire[31:0] addr_733_6;

Selector_2 s733_6(wires_183_5[1], addr_183_5, wires_733_6,addr_733_6);

wire[3:0] wires_734_6;

wire[31:0] addr_734_6;

Selector_2 s734_6(wires_183_5[2], addr_183_5, wires_734_6,addr_734_6);

wire[3:0] wires_735_6;

wire[31:0] addr_735_6;

Selector_2 s735_6(wires_183_5[3], addr_183_5, wires_735_6,addr_735_6);

wire[3:0] wires_736_6;

wire[31:0] addr_736_6;

Selector_2 s736_6(wires_184_5[0], addr_184_5, wires_736_6,addr_736_6);

wire[3:0] wires_737_6;

wire[31:0] addr_737_6;

Selector_2 s737_6(wires_184_5[1], addr_184_5, wires_737_6,addr_737_6);

wire[3:0] wires_738_6;

wire[31:0] addr_738_6;

Selector_2 s738_6(wires_184_5[2], addr_184_5, wires_738_6,addr_738_6);

wire[3:0] wires_739_6;

wire[31:0] addr_739_6;

Selector_2 s739_6(wires_184_5[3], addr_184_5, wires_739_6,addr_739_6);

wire[3:0] wires_740_6;

wire[31:0] addr_740_6;

Selector_2 s740_6(wires_185_5[0], addr_185_5, wires_740_6,addr_740_6);

wire[3:0] wires_741_6;

wire[31:0] addr_741_6;

Selector_2 s741_6(wires_185_5[1], addr_185_5, wires_741_6,addr_741_6);

wire[3:0] wires_742_6;

wire[31:0] addr_742_6;

Selector_2 s742_6(wires_185_5[2], addr_185_5, wires_742_6,addr_742_6);

wire[3:0] wires_743_6;

wire[31:0] addr_743_6;

Selector_2 s743_6(wires_185_5[3], addr_185_5, wires_743_6,addr_743_6);

wire[3:0] wires_744_6;

wire[31:0] addr_744_6;

Selector_2 s744_6(wires_186_5[0], addr_186_5, wires_744_6,addr_744_6);

wire[3:0] wires_745_6;

wire[31:0] addr_745_6;

Selector_2 s745_6(wires_186_5[1], addr_186_5, wires_745_6,addr_745_6);

wire[3:0] wires_746_6;

wire[31:0] addr_746_6;

Selector_2 s746_6(wires_186_5[2], addr_186_5, wires_746_6,addr_746_6);

wire[3:0] wires_747_6;

wire[31:0] addr_747_6;

Selector_2 s747_6(wires_186_5[3], addr_186_5, wires_747_6,addr_747_6);

wire[3:0] wires_748_6;

wire[31:0] addr_748_6;

Selector_2 s748_6(wires_187_5[0], addr_187_5, wires_748_6,addr_748_6);

wire[3:0] wires_749_6;

wire[31:0] addr_749_6;

Selector_2 s749_6(wires_187_5[1], addr_187_5, wires_749_6,addr_749_6);

wire[3:0] wires_750_6;

wire[31:0] addr_750_6;

Selector_2 s750_6(wires_187_5[2], addr_187_5, wires_750_6,addr_750_6);

wire[3:0] wires_751_6;

wire[31:0] addr_751_6;

Selector_2 s751_6(wires_187_5[3], addr_187_5, wires_751_6,addr_751_6);

wire[3:0] wires_752_6;

wire[31:0] addr_752_6;

Selector_2 s752_6(wires_188_5[0], addr_188_5, wires_752_6,addr_752_6);

wire[3:0] wires_753_6;

wire[31:0] addr_753_6;

Selector_2 s753_6(wires_188_5[1], addr_188_5, wires_753_6,addr_753_6);

wire[3:0] wires_754_6;

wire[31:0] addr_754_6;

Selector_2 s754_6(wires_188_5[2], addr_188_5, wires_754_6,addr_754_6);

wire[3:0] wires_755_6;

wire[31:0] addr_755_6;

Selector_2 s755_6(wires_188_5[3], addr_188_5, wires_755_6,addr_755_6);

wire[3:0] wires_756_6;

wire[31:0] addr_756_6;

Selector_2 s756_6(wires_189_5[0], addr_189_5, wires_756_6,addr_756_6);

wire[3:0] wires_757_6;

wire[31:0] addr_757_6;

Selector_2 s757_6(wires_189_5[1], addr_189_5, wires_757_6,addr_757_6);

wire[3:0] wires_758_6;

wire[31:0] addr_758_6;

Selector_2 s758_6(wires_189_5[2], addr_189_5, wires_758_6,addr_758_6);

wire[3:0] wires_759_6;

wire[31:0] addr_759_6;

Selector_2 s759_6(wires_189_5[3], addr_189_5, wires_759_6,addr_759_6);

wire[3:0] wires_760_6;

wire[31:0] addr_760_6;

Selector_2 s760_6(wires_190_5[0], addr_190_5, wires_760_6,addr_760_6);

wire[3:0] wires_761_6;

wire[31:0] addr_761_6;

Selector_2 s761_6(wires_190_5[1], addr_190_5, wires_761_6,addr_761_6);

wire[3:0] wires_762_6;

wire[31:0] addr_762_6;

Selector_2 s762_6(wires_190_5[2], addr_190_5, wires_762_6,addr_762_6);

wire[3:0] wires_763_6;

wire[31:0] addr_763_6;

Selector_2 s763_6(wires_190_5[3], addr_190_5, wires_763_6,addr_763_6);

wire[3:0] wires_764_6;

wire[31:0] addr_764_6;

Selector_2 s764_6(wires_191_5[0], addr_191_5, wires_764_6,addr_764_6);

wire[3:0] wires_765_6;

wire[31:0] addr_765_6;

Selector_2 s765_6(wires_191_5[1], addr_191_5, wires_765_6,addr_765_6);

wire[3:0] wires_766_6;

wire[31:0] addr_766_6;

Selector_2 s766_6(wires_191_5[2], addr_191_5, wires_766_6,addr_766_6);

wire[3:0] wires_767_6;

wire[31:0] addr_767_6;

Selector_2 s767_6(wires_191_5[3], addr_191_5, wires_767_6,addr_767_6);

wire[3:0] wires_768_6;

wire[31:0] addr_768_6;

Selector_2 s768_6(wires_192_5[0], addr_192_5, wires_768_6,addr_768_6);

wire[3:0] wires_769_6;

wire[31:0] addr_769_6;

Selector_2 s769_6(wires_192_5[1], addr_192_5, wires_769_6,addr_769_6);

wire[3:0] wires_770_6;

wire[31:0] addr_770_6;

Selector_2 s770_6(wires_192_5[2], addr_192_5, wires_770_6,addr_770_6);

wire[3:0] wires_771_6;

wire[31:0] addr_771_6;

Selector_2 s771_6(wires_192_5[3], addr_192_5, wires_771_6,addr_771_6);

wire[3:0] wires_772_6;

wire[31:0] addr_772_6;

Selector_2 s772_6(wires_193_5[0], addr_193_5, wires_772_6,addr_772_6);

wire[3:0] wires_773_6;

wire[31:0] addr_773_6;

Selector_2 s773_6(wires_193_5[1], addr_193_5, wires_773_6,addr_773_6);

wire[3:0] wires_774_6;

wire[31:0] addr_774_6;

Selector_2 s774_6(wires_193_5[2], addr_193_5, wires_774_6,addr_774_6);

wire[3:0] wires_775_6;

wire[31:0] addr_775_6;

Selector_2 s775_6(wires_193_5[3], addr_193_5, wires_775_6,addr_775_6);

wire[3:0] wires_776_6;

wire[31:0] addr_776_6;

Selector_2 s776_6(wires_194_5[0], addr_194_5, wires_776_6,addr_776_6);

wire[3:0] wires_777_6;

wire[31:0] addr_777_6;

Selector_2 s777_6(wires_194_5[1], addr_194_5, wires_777_6,addr_777_6);

wire[3:0] wires_778_6;

wire[31:0] addr_778_6;

Selector_2 s778_6(wires_194_5[2], addr_194_5, wires_778_6,addr_778_6);

wire[3:0] wires_779_6;

wire[31:0] addr_779_6;

Selector_2 s779_6(wires_194_5[3], addr_194_5, wires_779_6,addr_779_6);

wire[3:0] wires_780_6;

wire[31:0] addr_780_6;

Selector_2 s780_6(wires_195_5[0], addr_195_5, wires_780_6,addr_780_6);

wire[3:0] wires_781_6;

wire[31:0] addr_781_6;

Selector_2 s781_6(wires_195_5[1], addr_195_5, wires_781_6,addr_781_6);

wire[3:0] wires_782_6;

wire[31:0] addr_782_6;

Selector_2 s782_6(wires_195_5[2], addr_195_5, wires_782_6,addr_782_6);

wire[3:0] wires_783_6;

wire[31:0] addr_783_6;

Selector_2 s783_6(wires_195_5[3], addr_195_5, wires_783_6,addr_783_6);

wire[3:0] wires_784_6;

wire[31:0] addr_784_6;

Selector_2 s784_6(wires_196_5[0], addr_196_5, wires_784_6,addr_784_6);

wire[3:0] wires_785_6;

wire[31:0] addr_785_6;

Selector_2 s785_6(wires_196_5[1], addr_196_5, wires_785_6,addr_785_6);

wire[3:0] wires_786_6;

wire[31:0] addr_786_6;

Selector_2 s786_6(wires_196_5[2], addr_196_5, wires_786_6,addr_786_6);

wire[3:0] wires_787_6;

wire[31:0] addr_787_6;

Selector_2 s787_6(wires_196_5[3], addr_196_5, wires_787_6,addr_787_6);

wire[3:0] wires_788_6;

wire[31:0] addr_788_6;

Selector_2 s788_6(wires_197_5[0], addr_197_5, wires_788_6,addr_788_6);

wire[3:0] wires_789_6;

wire[31:0] addr_789_6;

Selector_2 s789_6(wires_197_5[1], addr_197_5, wires_789_6,addr_789_6);

wire[3:0] wires_790_6;

wire[31:0] addr_790_6;

Selector_2 s790_6(wires_197_5[2], addr_197_5, wires_790_6,addr_790_6);

wire[3:0] wires_791_6;

wire[31:0] addr_791_6;

Selector_2 s791_6(wires_197_5[3], addr_197_5, wires_791_6,addr_791_6);

wire[3:0] wires_792_6;

wire[31:0] addr_792_6;

Selector_2 s792_6(wires_198_5[0], addr_198_5, wires_792_6,addr_792_6);

wire[3:0] wires_793_6;

wire[31:0] addr_793_6;

Selector_2 s793_6(wires_198_5[1], addr_198_5, wires_793_6,addr_793_6);

wire[3:0] wires_794_6;

wire[31:0] addr_794_6;

Selector_2 s794_6(wires_198_5[2], addr_198_5, wires_794_6,addr_794_6);

wire[3:0] wires_795_6;

wire[31:0] addr_795_6;

Selector_2 s795_6(wires_198_5[3], addr_198_5, wires_795_6,addr_795_6);

wire[3:0] wires_796_6;

wire[31:0] addr_796_6;

Selector_2 s796_6(wires_199_5[0], addr_199_5, wires_796_6,addr_796_6);

wire[3:0] wires_797_6;

wire[31:0] addr_797_6;

Selector_2 s797_6(wires_199_5[1], addr_199_5, wires_797_6,addr_797_6);

wire[3:0] wires_798_6;

wire[31:0] addr_798_6;

Selector_2 s798_6(wires_199_5[2], addr_199_5, wires_798_6,addr_798_6);

wire[3:0] wires_799_6;

wire[31:0] addr_799_6;

Selector_2 s799_6(wires_199_5[3], addr_199_5, wires_799_6,addr_799_6);

wire[3:0] wires_800_6;

wire[31:0] addr_800_6;

Selector_2 s800_6(wires_200_5[0], addr_200_5, wires_800_6,addr_800_6);

wire[3:0] wires_801_6;

wire[31:0] addr_801_6;

Selector_2 s801_6(wires_200_5[1], addr_200_5, wires_801_6,addr_801_6);

wire[3:0] wires_802_6;

wire[31:0] addr_802_6;

Selector_2 s802_6(wires_200_5[2], addr_200_5, wires_802_6,addr_802_6);

wire[3:0] wires_803_6;

wire[31:0] addr_803_6;

Selector_2 s803_6(wires_200_5[3], addr_200_5, wires_803_6,addr_803_6);

wire[3:0] wires_804_6;

wire[31:0] addr_804_6;

Selector_2 s804_6(wires_201_5[0], addr_201_5, wires_804_6,addr_804_6);

wire[3:0] wires_805_6;

wire[31:0] addr_805_6;

Selector_2 s805_6(wires_201_5[1], addr_201_5, wires_805_6,addr_805_6);

wire[3:0] wires_806_6;

wire[31:0] addr_806_6;

Selector_2 s806_6(wires_201_5[2], addr_201_5, wires_806_6,addr_806_6);

wire[3:0] wires_807_6;

wire[31:0] addr_807_6;

Selector_2 s807_6(wires_201_5[3], addr_201_5, wires_807_6,addr_807_6);

wire[3:0] wires_808_6;

wire[31:0] addr_808_6;

Selector_2 s808_6(wires_202_5[0], addr_202_5, wires_808_6,addr_808_6);

wire[3:0] wires_809_6;

wire[31:0] addr_809_6;

Selector_2 s809_6(wires_202_5[1], addr_202_5, wires_809_6,addr_809_6);

wire[3:0] wires_810_6;

wire[31:0] addr_810_6;

Selector_2 s810_6(wires_202_5[2], addr_202_5, wires_810_6,addr_810_6);

wire[3:0] wires_811_6;

wire[31:0] addr_811_6;

Selector_2 s811_6(wires_202_5[3], addr_202_5, wires_811_6,addr_811_6);

wire[3:0] wires_812_6;

wire[31:0] addr_812_6;

Selector_2 s812_6(wires_203_5[0], addr_203_5, wires_812_6,addr_812_6);

wire[3:0] wires_813_6;

wire[31:0] addr_813_6;

Selector_2 s813_6(wires_203_5[1], addr_203_5, wires_813_6,addr_813_6);

wire[3:0] wires_814_6;

wire[31:0] addr_814_6;

Selector_2 s814_6(wires_203_5[2], addr_203_5, wires_814_6,addr_814_6);

wire[3:0] wires_815_6;

wire[31:0] addr_815_6;

Selector_2 s815_6(wires_203_5[3], addr_203_5, wires_815_6,addr_815_6);

wire[3:0] wires_816_6;

wire[31:0] addr_816_6;

Selector_2 s816_6(wires_204_5[0], addr_204_5, wires_816_6,addr_816_6);

wire[3:0] wires_817_6;

wire[31:0] addr_817_6;

Selector_2 s817_6(wires_204_5[1], addr_204_5, wires_817_6,addr_817_6);

wire[3:0] wires_818_6;

wire[31:0] addr_818_6;

Selector_2 s818_6(wires_204_5[2], addr_204_5, wires_818_6,addr_818_6);

wire[3:0] wires_819_6;

wire[31:0] addr_819_6;

Selector_2 s819_6(wires_204_5[3], addr_204_5, wires_819_6,addr_819_6);

wire[3:0] wires_820_6;

wire[31:0] addr_820_6;

Selector_2 s820_6(wires_205_5[0], addr_205_5, wires_820_6,addr_820_6);

wire[3:0] wires_821_6;

wire[31:0] addr_821_6;

Selector_2 s821_6(wires_205_5[1], addr_205_5, wires_821_6,addr_821_6);

wire[3:0] wires_822_6;

wire[31:0] addr_822_6;

Selector_2 s822_6(wires_205_5[2], addr_205_5, wires_822_6,addr_822_6);

wire[3:0] wires_823_6;

wire[31:0] addr_823_6;

Selector_2 s823_6(wires_205_5[3], addr_205_5, wires_823_6,addr_823_6);

wire[3:0] wires_824_6;

wire[31:0] addr_824_6;

Selector_2 s824_6(wires_206_5[0], addr_206_5, wires_824_6,addr_824_6);

wire[3:0] wires_825_6;

wire[31:0] addr_825_6;

Selector_2 s825_6(wires_206_5[1], addr_206_5, wires_825_6,addr_825_6);

wire[3:0] wires_826_6;

wire[31:0] addr_826_6;

Selector_2 s826_6(wires_206_5[2], addr_206_5, wires_826_6,addr_826_6);

wire[3:0] wires_827_6;

wire[31:0] addr_827_6;

Selector_2 s827_6(wires_206_5[3], addr_206_5, wires_827_6,addr_827_6);

wire[3:0] wires_828_6;

wire[31:0] addr_828_6;

Selector_2 s828_6(wires_207_5[0], addr_207_5, wires_828_6,addr_828_6);

wire[3:0] wires_829_6;

wire[31:0] addr_829_6;

Selector_2 s829_6(wires_207_5[1], addr_207_5, wires_829_6,addr_829_6);

wire[3:0] wires_830_6;

wire[31:0] addr_830_6;

Selector_2 s830_6(wires_207_5[2], addr_207_5, wires_830_6,addr_830_6);

wire[3:0] wires_831_6;

wire[31:0] addr_831_6;

Selector_2 s831_6(wires_207_5[3], addr_207_5, wires_831_6,addr_831_6);

wire[3:0] wires_832_6;

wire[31:0] addr_832_6;

Selector_2 s832_6(wires_208_5[0], addr_208_5, wires_832_6,addr_832_6);

wire[3:0] wires_833_6;

wire[31:0] addr_833_6;

Selector_2 s833_6(wires_208_5[1], addr_208_5, wires_833_6,addr_833_6);

wire[3:0] wires_834_6;

wire[31:0] addr_834_6;

Selector_2 s834_6(wires_208_5[2], addr_208_5, wires_834_6,addr_834_6);

wire[3:0] wires_835_6;

wire[31:0] addr_835_6;

Selector_2 s835_6(wires_208_5[3], addr_208_5, wires_835_6,addr_835_6);

wire[3:0] wires_836_6;

wire[31:0] addr_836_6;

Selector_2 s836_6(wires_209_5[0], addr_209_5, wires_836_6,addr_836_6);

wire[3:0] wires_837_6;

wire[31:0] addr_837_6;

Selector_2 s837_6(wires_209_5[1], addr_209_5, wires_837_6,addr_837_6);

wire[3:0] wires_838_6;

wire[31:0] addr_838_6;

Selector_2 s838_6(wires_209_5[2], addr_209_5, wires_838_6,addr_838_6);

wire[3:0] wires_839_6;

wire[31:0] addr_839_6;

Selector_2 s839_6(wires_209_5[3], addr_209_5, wires_839_6,addr_839_6);

wire[3:0] wires_840_6;

wire[31:0] addr_840_6;

Selector_2 s840_6(wires_210_5[0], addr_210_5, wires_840_6,addr_840_6);

wire[3:0] wires_841_6;

wire[31:0] addr_841_6;

Selector_2 s841_6(wires_210_5[1], addr_210_5, wires_841_6,addr_841_6);

wire[3:0] wires_842_6;

wire[31:0] addr_842_6;

Selector_2 s842_6(wires_210_5[2], addr_210_5, wires_842_6,addr_842_6);

wire[3:0] wires_843_6;

wire[31:0] addr_843_6;

Selector_2 s843_6(wires_210_5[3], addr_210_5, wires_843_6,addr_843_6);

wire[3:0] wires_844_6;

wire[31:0] addr_844_6;

Selector_2 s844_6(wires_211_5[0], addr_211_5, wires_844_6,addr_844_6);

wire[3:0] wires_845_6;

wire[31:0] addr_845_6;

Selector_2 s845_6(wires_211_5[1], addr_211_5, wires_845_6,addr_845_6);

wire[3:0] wires_846_6;

wire[31:0] addr_846_6;

Selector_2 s846_6(wires_211_5[2], addr_211_5, wires_846_6,addr_846_6);

wire[3:0] wires_847_6;

wire[31:0] addr_847_6;

Selector_2 s847_6(wires_211_5[3], addr_211_5, wires_847_6,addr_847_6);

wire[3:0] wires_848_6;

wire[31:0] addr_848_6;

Selector_2 s848_6(wires_212_5[0], addr_212_5, wires_848_6,addr_848_6);

wire[3:0] wires_849_6;

wire[31:0] addr_849_6;

Selector_2 s849_6(wires_212_5[1], addr_212_5, wires_849_6,addr_849_6);

wire[3:0] wires_850_6;

wire[31:0] addr_850_6;

Selector_2 s850_6(wires_212_5[2], addr_212_5, wires_850_6,addr_850_6);

wire[3:0] wires_851_6;

wire[31:0] addr_851_6;

Selector_2 s851_6(wires_212_5[3], addr_212_5, wires_851_6,addr_851_6);

wire[3:0] wires_852_6;

wire[31:0] addr_852_6;

Selector_2 s852_6(wires_213_5[0], addr_213_5, wires_852_6,addr_852_6);

wire[3:0] wires_853_6;

wire[31:0] addr_853_6;

Selector_2 s853_6(wires_213_5[1], addr_213_5, wires_853_6,addr_853_6);

wire[3:0] wires_854_6;

wire[31:0] addr_854_6;

Selector_2 s854_6(wires_213_5[2], addr_213_5, wires_854_6,addr_854_6);

wire[3:0] wires_855_6;

wire[31:0] addr_855_6;

Selector_2 s855_6(wires_213_5[3], addr_213_5, wires_855_6,addr_855_6);

wire[3:0] wires_856_6;

wire[31:0] addr_856_6;

Selector_2 s856_6(wires_214_5[0], addr_214_5, wires_856_6,addr_856_6);

wire[3:0] wires_857_6;

wire[31:0] addr_857_6;

Selector_2 s857_6(wires_214_5[1], addr_214_5, wires_857_6,addr_857_6);

wire[3:0] wires_858_6;

wire[31:0] addr_858_6;

Selector_2 s858_6(wires_214_5[2], addr_214_5, wires_858_6,addr_858_6);

wire[3:0] wires_859_6;

wire[31:0] addr_859_6;

Selector_2 s859_6(wires_214_5[3], addr_214_5, wires_859_6,addr_859_6);

wire[3:0] wires_860_6;

wire[31:0] addr_860_6;

Selector_2 s860_6(wires_215_5[0], addr_215_5, wires_860_6,addr_860_6);

wire[3:0] wires_861_6;

wire[31:0] addr_861_6;

Selector_2 s861_6(wires_215_5[1], addr_215_5, wires_861_6,addr_861_6);

wire[3:0] wires_862_6;

wire[31:0] addr_862_6;

Selector_2 s862_6(wires_215_5[2], addr_215_5, wires_862_6,addr_862_6);

wire[3:0] wires_863_6;

wire[31:0] addr_863_6;

Selector_2 s863_6(wires_215_5[3], addr_215_5, wires_863_6,addr_863_6);

wire[3:0] wires_864_6;

wire[31:0] addr_864_6;

Selector_2 s864_6(wires_216_5[0], addr_216_5, wires_864_6,addr_864_6);

wire[3:0] wires_865_6;

wire[31:0] addr_865_6;

Selector_2 s865_6(wires_216_5[1], addr_216_5, wires_865_6,addr_865_6);

wire[3:0] wires_866_6;

wire[31:0] addr_866_6;

Selector_2 s866_6(wires_216_5[2], addr_216_5, wires_866_6,addr_866_6);

wire[3:0] wires_867_6;

wire[31:0] addr_867_6;

Selector_2 s867_6(wires_216_5[3], addr_216_5, wires_867_6,addr_867_6);

wire[3:0] wires_868_6;

wire[31:0] addr_868_6;

Selector_2 s868_6(wires_217_5[0], addr_217_5, wires_868_6,addr_868_6);

wire[3:0] wires_869_6;

wire[31:0] addr_869_6;

Selector_2 s869_6(wires_217_5[1], addr_217_5, wires_869_6,addr_869_6);

wire[3:0] wires_870_6;

wire[31:0] addr_870_6;

Selector_2 s870_6(wires_217_5[2], addr_217_5, wires_870_6,addr_870_6);

wire[3:0] wires_871_6;

wire[31:0] addr_871_6;

Selector_2 s871_6(wires_217_5[3], addr_217_5, wires_871_6,addr_871_6);

wire[3:0] wires_872_6;

wire[31:0] addr_872_6;

Selector_2 s872_6(wires_218_5[0], addr_218_5, wires_872_6,addr_872_6);

wire[3:0] wires_873_6;

wire[31:0] addr_873_6;

Selector_2 s873_6(wires_218_5[1], addr_218_5, wires_873_6,addr_873_6);

wire[3:0] wires_874_6;

wire[31:0] addr_874_6;

Selector_2 s874_6(wires_218_5[2], addr_218_5, wires_874_6,addr_874_6);

wire[3:0] wires_875_6;

wire[31:0] addr_875_6;

Selector_2 s875_6(wires_218_5[3], addr_218_5, wires_875_6,addr_875_6);

wire[3:0] wires_876_6;

wire[31:0] addr_876_6;

Selector_2 s876_6(wires_219_5[0], addr_219_5, wires_876_6,addr_876_6);

wire[3:0] wires_877_6;

wire[31:0] addr_877_6;

Selector_2 s877_6(wires_219_5[1], addr_219_5, wires_877_6,addr_877_6);

wire[3:0] wires_878_6;

wire[31:0] addr_878_6;

Selector_2 s878_6(wires_219_5[2], addr_219_5, wires_878_6,addr_878_6);

wire[3:0] wires_879_6;

wire[31:0] addr_879_6;

Selector_2 s879_6(wires_219_5[3], addr_219_5, wires_879_6,addr_879_6);

wire[3:0] wires_880_6;

wire[31:0] addr_880_6;

Selector_2 s880_6(wires_220_5[0], addr_220_5, wires_880_6,addr_880_6);

wire[3:0] wires_881_6;

wire[31:0] addr_881_6;

Selector_2 s881_6(wires_220_5[1], addr_220_5, wires_881_6,addr_881_6);

wire[3:0] wires_882_6;

wire[31:0] addr_882_6;

Selector_2 s882_6(wires_220_5[2], addr_220_5, wires_882_6,addr_882_6);

wire[3:0] wires_883_6;

wire[31:0] addr_883_6;

Selector_2 s883_6(wires_220_5[3], addr_220_5, wires_883_6,addr_883_6);

wire[3:0] wires_884_6;

wire[31:0] addr_884_6;

Selector_2 s884_6(wires_221_5[0], addr_221_5, wires_884_6,addr_884_6);

wire[3:0] wires_885_6;

wire[31:0] addr_885_6;

Selector_2 s885_6(wires_221_5[1], addr_221_5, wires_885_6,addr_885_6);

wire[3:0] wires_886_6;

wire[31:0] addr_886_6;

Selector_2 s886_6(wires_221_5[2], addr_221_5, wires_886_6,addr_886_6);

wire[3:0] wires_887_6;

wire[31:0] addr_887_6;

Selector_2 s887_6(wires_221_5[3], addr_221_5, wires_887_6,addr_887_6);

wire[3:0] wires_888_6;

wire[31:0] addr_888_6;

Selector_2 s888_6(wires_222_5[0], addr_222_5, wires_888_6,addr_888_6);

wire[3:0] wires_889_6;

wire[31:0] addr_889_6;

Selector_2 s889_6(wires_222_5[1], addr_222_5, wires_889_6,addr_889_6);

wire[3:0] wires_890_6;

wire[31:0] addr_890_6;

Selector_2 s890_6(wires_222_5[2], addr_222_5, wires_890_6,addr_890_6);

wire[3:0] wires_891_6;

wire[31:0] addr_891_6;

Selector_2 s891_6(wires_222_5[3], addr_222_5, wires_891_6,addr_891_6);

wire[3:0] wires_892_6;

wire[31:0] addr_892_6;

Selector_2 s892_6(wires_223_5[0], addr_223_5, wires_892_6,addr_892_6);

wire[3:0] wires_893_6;

wire[31:0] addr_893_6;

Selector_2 s893_6(wires_223_5[1], addr_223_5, wires_893_6,addr_893_6);

wire[3:0] wires_894_6;

wire[31:0] addr_894_6;

Selector_2 s894_6(wires_223_5[2], addr_223_5, wires_894_6,addr_894_6);

wire[3:0] wires_895_6;

wire[31:0] addr_895_6;

Selector_2 s895_6(wires_223_5[3], addr_223_5, wires_895_6,addr_895_6);

wire[3:0] wires_896_6;

wire[31:0] addr_896_6;

Selector_2 s896_6(wires_224_5[0], addr_224_5, wires_896_6,addr_896_6);

wire[3:0] wires_897_6;

wire[31:0] addr_897_6;

Selector_2 s897_6(wires_224_5[1], addr_224_5, wires_897_6,addr_897_6);

wire[3:0] wires_898_6;

wire[31:0] addr_898_6;

Selector_2 s898_6(wires_224_5[2], addr_224_5, wires_898_6,addr_898_6);

wire[3:0] wires_899_6;

wire[31:0] addr_899_6;

Selector_2 s899_6(wires_224_5[3], addr_224_5, wires_899_6,addr_899_6);

wire[3:0] wires_900_6;

wire[31:0] addr_900_6;

Selector_2 s900_6(wires_225_5[0], addr_225_5, wires_900_6,addr_900_6);

wire[3:0] wires_901_6;

wire[31:0] addr_901_6;

Selector_2 s901_6(wires_225_5[1], addr_225_5, wires_901_6,addr_901_6);

wire[3:0] wires_902_6;

wire[31:0] addr_902_6;

Selector_2 s902_6(wires_225_5[2], addr_225_5, wires_902_6,addr_902_6);

wire[3:0] wires_903_6;

wire[31:0] addr_903_6;

Selector_2 s903_6(wires_225_5[3], addr_225_5, wires_903_6,addr_903_6);

wire[3:0] wires_904_6;

wire[31:0] addr_904_6;

Selector_2 s904_6(wires_226_5[0], addr_226_5, wires_904_6,addr_904_6);

wire[3:0] wires_905_6;

wire[31:0] addr_905_6;

Selector_2 s905_6(wires_226_5[1], addr_226_5, wires_905_6,addr_905_6);

wire[3:0] wires_906_6;

wire[31:0] addr_906_6;

Selector_2 s906_6(wires_226_5[2], addr_226_5, wires_906_6,addr_906_6);

wire[3:0] wires_907_6;

wire[31:0] addr_907_6;

Selector_2 s907_6(wires_226_5[3], addr_226_5, wires_907_6,addr_907_6);

wire[3:0] wires_908_6;

wire[31:0] addr_908_6;

Selector_2 s908_6(wires_227_5[0], addr_227_5, wires_908_6,addr_908_6);

wire[3:0] wires_909_6;

wire[31:0] addr_909_6;

Selector_2 s909_6(wires_227_5[1], addr_227_5, wires_909_6,addr_909_6);

wire[3:0] wires_910_6;

wire[31:0] addr_910_6;

Selector_2 s910_6(wires_227_5[2], addr_227_5, wires_910_6,addr_910_6);

wire[3:0] wires_911_6;

wire[31:0] addr_911_6;

Selector_2 s911_6(wires_227_5[3], addr_227_5, wires_911_6,addr_911_6);

wire[3:0] wires_912_6;

wire[31:0] addr_912_6;

Selector_2 s912_6(wires_228_5[0], addr_228_5, wires_912_6,addr_912_6);

wire[3:0] wires_913_6;

wire[31:0] addr_913_6;

Selector_2 s913_6(wires_228_5[1], addr_228_5, wires_913_6,addr_913_6);

wire[3:0] wires_914_6;

wire[31:0] addr_914_6;

Selector_2 s914_6(wires_228_5[2], addr_228_5, wires_914_6,addr_914_6);

wire[3:0] wires_915_6;

wire[31:0] addr_915_6;

Selector_2 s915_6(wires_228_5[3], addr_228_5, wires_915_6,addr_915_6);

wire[3:0] wires_916_6;

wire[31:0] addr_916_6;

Selector_2 s916_6(wires_229_5[0], addr_229_5, wires_916_6,addr_916_6);

wire[3:0] wires_917_6;

wire[31:0] addr_917_6;

Selector_2 s917_6(wires_229_5[1], addr_229_5, wires_917_6,addr_917_6);

wire[3:0] wires_918_6;

wire[31:0] addr_918_6;

Selector_2 s918_6(wires_229_5[2], addr_229_5, wires_918_6,addr_918_6);

wire[3:0] wires_919_6;

wire[31:0] addr_919_6;

Selector_2 s919_6(wires_229_5[3], addr_229_5, wires_919_6,addr_919_6);

wire[3:0] wires_920_6;

wire[31:0] addr_920_6;

Selector_2 s920_6(wires_230_5[0], addr_230_5, wires_920_6,addr_920_6);

wire[3:0] wires_921_6;

wire[31:0] addr_921_6;

Selector_2 s921_6(wires_230_5[1], addr_230_5, wires_921_6,addr_921_6);

wire[3:0] wires_922_6;

wire[31:0] addr_922_6;

Selector_2 s922_6(wires_230_5[2], addr_230_5, wires_922_6,addr_922_6);

wire[3:0] wires_923_6;

wire[31:0] addr_923_6;

Selector_2 s923_6(wires_230_5[3], addr_230_5, wires_923_6,addr_923_6);

wire[3:0] wires_924_6;

wire[31:0] addr_924_6;

Selector_2 s924_6(wires_231_5[0], addr_231_5, wires_924_6,addr_924_6);

wire[3:0] wires_925_6;

wire[31:0] addr_925_6;

Selector_2 s925_6(wires_231_5[1], addr_231_5, wires_925_6,addr_925_6);

wire[3:0] wires_926_6;

wire[31:0] addr_926_6;

Selector_2 s926_6(wires_231_5[2], addr_231_5, wires_926_6,addr_926_6);

wire[3:0] wires_927_6;

wire[31:0] addr_927_6;

Selector_2 s927_6(wires_231_5[3], addr_231_5, wires_927_6,addr_927_6);

wire[3:0] wires_928_6;

wire[31:0] addr_928_6;

Selector_2 s928_6(wires_232_5[0], addr_232_5, wires_928_6,addr_928_6);

wire[3:0] wires_929_6;

wire[31:0] addr_929_6;

Selector_2 s929_6(wires_232_5[1], addr_232_5, wires_929_6,addr_929_6);

wire[3:0] wires_930_6;

wire[31:0] addr_930_6;

Selector_2 s930_6(wires_232_5[2], addr_232_5, wires_930_6,addr_930_6);

wire[3:0] wires_931_6;

wire[31:0] addr_931_6;

Selector_2 s931_6(wires_232_5[3], addr_232_5, wires_931_6,addr_931_6);

wire[3:0] wires_932_6;

wire[31:0] addr_932_6;

Selector_2 s932_6(wires_233_5[0], addr_233_5, wires_932_6,addr_932_6);

wire[3:0] wires_933_6;

wire[31:0] addr_933_6;

Selector_2 s933_6(wires_233_5[1], addr_233_5, wires_933_6,addr_933_6);

wire[3:0] wires_934_6;

wire[31:0] addr_934_6;

Selector_2 s934_6(wires_233_5[2], addr_233_5, wires_934_6,addr_934_6);

wire[3:0] wires_935_6;

wire[31:0] addr_935_6;

Selector_2 s935_6(wires_233_5[3], addr_233_5, wires_935_6,addr_935_6);

wire[3:0] wires_936_6;

wire[31:0] addr_936_6;

Selector_2 s936_6(wires_234_5[0], addr_234_5, wires_936_6,addr_936_6);

wire[3:0] wires_937_6;

wire[31:0] addr_937_6;

Selector_2 s937_6(wires_234_5[1], addr_234_5, wires_937_6,addr_937_6);

wire[3:0] wires_938_6;

wire[31:0] addr_938_6;

Selector_2 s938_6(wires_234_5[2], addr_234_5, wires_938_6,addr_938_6);

wire[3:0] wires_939_6;

wire[31:0] addr_939_6;

Selector_2 s939_6(wires_234_5[3], addr_234_5, wires_939_6,addr_939_6);

wire[3:0] wires_940_6;

wire[31:0] addr_940_6;

Selector_2 s940_6(wires_235_5[0], addr_235_5, wires_940_6,addr_940_6);

wire[3:0] wires_941_6;

wire[31:0] addr_941_6;

Selector_2 s941_6(wires_235_5[1], addr_235_5, wires_941_6,addr_941_6);

wire[3:0] wires_942_6;

wire[31:0] addr_942_6;

Selector_2 s942_6(wires_235_5[2], addr_235_5, wires_942_6,addr_942_6);

wire[3:0] wires_943_6;

wire[31:0] addr_943_6;

Selector_2 s943_6(wires_235_5[3], addr_235_5, wires_943_6,addr_943_6);

wire[3:0] wires_944_6;

wire[31:0] addr_944_6;

Selector_2 s944_6(wires_236_5[0], addr_236_5, wires_944_6,addr_944_6);

wire[3:0] wires_945_6;

wire[31:0] addr_945_6;

Selector_2 s945_6(wires_236_5[1], addr_236_5, wires_945_6,addr_945_6);

wire[3:0] wires_946_6;

wire[31:0] addr_946_6;

Selector_2 s946_6(wires_236_5[2], addr_236_5, wires_946_6,addr_946_6);

wire[3:0] wires_947_6;

wire[31:0] addr_947_6;

Selector_2 s947_6(wires_236_5[3], addr_236_5, wires_947_6,addr_947_6);

wire[3:0] wires_948_6;

wire[31:0] addr_948_6;

Selector_2 s948_6(wires_237_5[0], addr_237_5, wires_948_6,addr_948_6);

wire[3:0] wires_949_6;

wire[31:0] addr_949_6;

Selector_2 s949_6(wires_237_5[1], addr_237_5, wires_949_6,addr_949_6);

wire[3:0] wires_950_6;

wire[31:0] addr_950_6;

Selector_2 s950_6(wires_237_5[2], addr_237_5, wires_950_6,addr_950_6);

wire[3:0] wires_951_6;

wire[31:0] addr_951_6;

Selector_2 s951_6(wires_237_5[3], addr_237_5, wires_951_6,addr_951_6);

wire[3:0] wires_952_6;

wire[31:0] addr_952_6;

Selector_2 s952_6(wires_238_5[0], addr_238_5, wires_952_6,addr_952_6);

wire[3:0] wires_953_6;

wire[31:0] addr_953_6;

Selector_2 s953_6(wires_238_5[1], addr_238_5, wires_953_6,addr_953_6);

wire[3:0] wires_954_6;

wire[31:0] addr_954_6;

Selector_2 s954_6(wires_238_5[2], addr_238_5, wires_954_6,addr_954_6);

wire[3:0] wires_955_6;

wire[31:0] addr_955_6;

Selector_2 s955_6(wires_238_5[3], addr_238_5, wires_955_6,addr_955_6);

wire[3:0] wires_956_6;

wire[31:0] addr_956_6;

Selector_2 s956_6(wires_239_5[0], addr_239_5, wires_956_6,addr_956_6);

wire[3:0] wires_957_6;

wire[31:0] addr_957_6;

Selector_2 s957_6(wires_239_5[1], addr_239_5, wires_957_6,addr_957_6);

wire[3:0] wires_958_6;

wire[31:0] addr_958_6;

Selector_2 s958_6(wires_239_5[2], addr_239_5, wires_958_6,addr_958_6);

wire[3:0] wires_959_6;

wire[31:0] addr_959_6;

Selector_2 s959_6(wires_239_5[3], addr_239_5, wires_959_6,addr_959_6);

wire[3:0] wires_960_6;

wire[31:0] addr_960_6;

Selector_2 s960_6(wires_240_5[0], addr_240_5, wires_960_6,addr_960_6);

wire[3:0] wires_961_6;

wire[31:0] addr_961_6;

Selector_2 s961_6(wires_240_5[1], addr_240_5, wires_961_6,addr_961_6);

wire[3:0] wires_962_6;

wire[31:0] addr_962_6;

Selector_2 s962_6(wires_240_5[2], addr_240_5, wires_962_6,addr_962_6);

wire[3:0] wires_963_6;

wire[31:0] addr_963_6;

Selector_2 s963_6(wires_240_5[3], addr_240_5, wires_963_6,addr_963_6);

wire[3:0] wires_964_6;

wire[31:0] addr_964_6;

Selector_2 s964_6(wires_241_5[0], addr_241_5, wires_964_6,addr_964_6);

wire[3:0] wires_965_6;

wire[31:0] addr_965_6;

Selector_2 s965_6(wires_241_5[1], addr_241_5, wires_965_6,addr_965_6);

wire[3:0] wires_966_6;

wire[31:0] addr_966_6;

Selector_2 s966_6(wires_241_5[2], addr_241_5, wires_966_6,addr_966_6);

wire[3:0] wires_967_6;

wire[31:0] addr_967_6;

Selector_2 s967_6(wires_241_5[3], addr_241_5, wires_967_6,addr_967_6);

wire[3:0] wires_968_6;

wire[31:0] addr_968_6;

Selector_2 s968_6(wires_242_5[0], addr_242_5, wires_968_6,addr_968_6);

wire[3:0] wires_969_6;

wire[31:0] addr_969_6;

Selector_2 s969_6(wires_242_5[1], addr_242_5, wires_969_6,addr_969_6);

wire[3:0] wires_970_6;

wire[31:0] addr_970_6;

Selector_2 s970_6(wires_242_5[2], addr_242_5, wires_970_6,addr_970_6);

wire[3:0] wires_971_6;

wire[31:0] addr_971_6;

Selector_2 s971_6(wires_242_5[3], addr_242_5, wires_971_6,addr_971_6);

wire[3:0] wires_972_6;

wire[31:0] addr_972_6;

Selector_2 s972_6(wires_243_5[0], addr_243_5, wires_972_6,addr_972_6);

wire[3:0] wires_973_6;

wire[31:0] addr_973_6;

Selector_2 s973_6(wires_243_5[1], addr_243_5, wires_973_6,addr_973_6);

wire[3:0] wires_974_6;

wire[31:0] addr_974_6;

Selector_2 s974_6(wires_243_5[2], addr_243_5, wires_974_6,addr_974_6);

wire[3:0] wires_975_6;

wire[31:0] addr_975_6;

Selector_2 s975_6(wires_243_5[3], addr_243_5, wires_975_6,addr_975_6);

wire[3:0] wires_976_6;

wire[31:0] addr_976_6;

Selector_2 s976_6(wires_244_5[0], addr_244_5, wires_976_6,addr_976_6);

wire[3:0] wires_977_6;

wire[31:0] addr_977_6;

Selector_2 s977_6(wires_244_5[1], addr_244_5, wires_977_6,addr_977_6);

wire[3:0] wires_978_6;

wire[31:0] addr_978_6;

Selector_2 s978_6(wires_244_5[2], addr_244_5, wires_978_6,addr_978_6);

wire[3:0] wires_979_6;

wire[31:0] addr_979_6;

Selector_2 s979_6(wires_244_5[3], addr_244_5, wires_979_6,addr_979_6);

wire[3:0] wires_980_6;

wire[31:0] addr_980_6;

Selector_2 s980_6(wires_245_5[0], addr_245_5, wires_980_6,addr_980_6);

wire[3:0] wires_981_6;

wire[31:0] addr_981_6;

Selector_2 s981_6(wires_245_5[1], addr_245_5, wires_981_6,addr_981_6);

wire[3:0] wires_982_6;

wire[31:0] addr_982_6;

Selector_2 s982_6(wires_245_5[2], addr_245_5, wires_982_6,addr_982_6);

wire[3:0] wires_983_6;

wire[31:0] addr_983_6;

Selector_2 s983_6(wires_245_5[3], addr_245_5, wires_983_6,addr_983_6);

wire[3:0] wires_984_6;

wire[31:0] addr_984_6;

Selector_2 s984_6(wires_246_5[0], addr_246_5, wires_984_6,addr_984_6);

wire[3:0] wires_985_6;

wire[31:0] addr_985_6;

Selector_2 s985_6(wires_246_5[1], addr_246_5, wires_985_6,addr_985_6);

wire[3:0] wires_986_6;

wire[31:0] addr_986_6;

Selector_2 s986_6(wires_246_5[2], addr_246_5, wires_986_6,addr_986_6);

wire[3:0] wires_987_6;

wire[31:0] addr_987_6;

Selector_2 s987_6(wires_246_5[3], addr_246_5, wires_987_6,addr_987_6);

wire[3:0] wires_988_6;

wire[31:0] addr_988_6;

Selector_2 s988_6(wires_247_5[0], addr_247_5, wires_988_6,addr_988_6);

wire[3:0] wires_989_6;

wire[31:0] addr_989_6;

Selector_2 s989_6(wires_247_5[1], addr_247_5, wires_989_6,addr_989_6);

wire[3:0] wires_990_6;

wire[31:0] addr_990_6;

Selector_2 s990_6(wires_247_5[2], addr_247_5, wires_990_6,addr_990_6);

wire[3:0] wires_991_6;

wire[31:0] addr_991_6;

Selector_2 s991_6(wires_247_5[3], addr_247_5, wires_991_6,addr_991_6);

wire[3:0] wires_992_6;

wire[31:0] addr_992_6;

Selector_2 s992_6(wires_248_5[0], addr_248_5, wires_992_6,addr_992_6);

wire[3:0] wires_993_6;

wire[31:0] addr_993_6;

Selector_2 s993_6(wires_248_5[1], addr_248_5, wires_993_6,addr_993_6);

wire[3:0] wires_994_6;

wire[31:0] addr_994_6;

Selector_2 s994_6(wires_248_5[2], addr_248_5, wires_994_6,addr_994_6);

wire[3:0] wires_995_6;

wire[31:0] addr_995_6;

Selector_2 s995_6(wires_248_5[3], addr_248_5, wires_995_6,addr_995_6);

wire[3:0] wires_996_6;

wire[31:0] addr_996_6;

Selector_2 s996_6(wires_249_5[0], addr_249_5, wires_996_6,addr_996_6);

wire[3:0] wires_997_6;

wire[31:0] addr_997_6;

Selector_2 s997_6(wires_249_5[1], addr_249_5, wires_997_6,addr_997_6);

wire[3:0] wires_998_6;

wire[31:0] addr_998_6;

Selector_2 s998_6(wires_249_5[2], addr_249_5, wires_998_6,addr_998_6);

wire[3:0] wires_999_6;

wire[31:0] addr_999_6;

Selector_2 s999_6(wires_249_5[3], addr_249_5, wires_999_6,addr_999_6);

wire[3:0] wires_1000_6;

wire[31:0] addr_1000_6;

Selector_2 s1000_6(wires_250_5[0], addr_250_5, wires_1000_6,addr_1000_6);

wire[3:0] wires_1001_6;

wire[31:0] addr_1001_6;

Selector_2 s1001_6(wires_250_5[1], addr_250_5, wires_1001_6,addr_1001_6);

wire[3:0] wires_1002_6;

wire[31:0] addr_1002_6;

Selector_2 s1002_6(wires_250_5[2], addr_250_5, wires_1002_6,addr_1002_6);

wire[3:0] wires_1003_6;

wire[31:0] addr_1003_6;

Selector_2 s1003_6(wires_250_5[3], addr_250_5, wires_1003_6,addr_1003_6);

wire[3:0] wires_1004_6;

wire[31:0] addr_1004_6;

Selector_2 s1004_6(wires_251_5[0], addr_251_5, wires_1004_6,addr_1004_6);

wire[3:0] wires_1005_6;

wire[31:0] addr_1005_6;

Selector_2 s1005_6(wires_251_5[1], addr_251_5, wires_1005_6,addr_1005_6);

wire[3:0] wires_1006_6;

wire[31:0] addr_1006_6;

Selector_2 s1006_6(wires_251_5[2], addr_251_5, wires_1006_6,addr_1006_6);

wire[3:0] wires_1007_6;

wire[31:0] addr_1007_6;

Selector_2 s1007_6(wires_251_5[3], addr_251_5, wires_1007_6,addr_1007_6);

wire[3:0] wires_1008_6;

wire[31:0] addr_1008_6;

Selector_2 s1008_6(wires_252_5[0], addr_252_5, wires_1008_6,addr_1008_6);

wire[3:0] wires_1009_6;

wire[31:0] addr_1009_6;

Selector_2 s1009_6(wires_252_5[1], addr_252_5, wires_1009_6,addr_1009_6);

wire[3:0] wires_1010_6;

wire[31:0] addr_1010_6;

Selector_2 s1010_6(wires_252_5[2], addr_252_5, wires_1010_6,addr_1010_6);

wire[3:0] wires_1011_6;

wire[31:0] addr_1011_6;

Selector_2 s1011_6(wires_252_5[3], addr_252_5, wires_1011_6,addr_1011_6);

wire[3:0] wires_1012_6;

wire[31:0] addr_1012_6;

Selector_2 s1012_6(wires_253_5[0], addr_253_5, wires_1012_6,addr_1012_6);

wire[3:0] wires_1013_6;

wire[31:0] addr_1013_6;

Selector_2 s1013_6(wires_253_5[1], addr_253_5, wires_1013_6,addr_1013_6);

wire[3:0] wires_1014_6;

wire[31:0] addr_1014_6;

Selector_2 s1014_6(wires_253_5[2], addr_253_5, wires_1014_6,addr_1014_6);

wire[3:0] wires_1015_6;

wire[31:0] addr_1015_6;

Selector_2 s1015_6(wires_253_5[3], addr_253_5, wires_1015_6,addr_1015_6);

wire[3:0] wires_1016_6;

wire[31:0] addr_1016_6;

Selector_2 s1016_6(wires_254_5[0], addr_254_5, wires_1016_6,addr_1016_6);

wire[3:0] wires_1017_6;

wire[31:0] addr_1017_6;

Selector_2 s1017_6(wires_254_5[1], addr_254_5, wires_1017_6,addr_1017_6);

wire[3:0] wires_1018_6;

wire[31:0] addr_1018_6;

Selector_2 s1018_6(wires_254_5[2], addr_254_5, wires_1018_6,addr_1018_6);

wire[3:0] wires_1019_6;

wire[31:0] addr_1019_6;

Selector_2 s1019_6(wires_254_5[3], addr_254_5, wires_1019_6,addr_1019_6);

wire[3:0] wires_1020_6;

wire[31:0] addr_1020_6;

Selector_2 s1020_6(wires_255_5[0], addr_255_5, wires_1020_6,addr_1020_6);

wire[3:0] wires_1021_6;

wire[31:0] addr_1021_6;

Selector_2 s1021_6(wires_255_5[1], addr_255_5, wires_1021_6,addr_1021_6);

wire[3:0] wires_1022_6;

wire[31:0] addr_1022_6;

Selector_2 s1022_6(wires_255_5[2], addr_255_5, wires_1022_6,addr_1022_6);

wire[3:0] wires_1023_6;

wire[31:0] addr_1023_6;

Selector_2 s1023_6(wires_255_5[3], addr_255_5, wires_1023_6,addr_1023_6);

wire[3:0] wires_1024_6;

wire[31:0] addr_1024_6;

Selector_2 s1024_6(wires_256_5[0], addr_256_5, wires_1024_6,addr_1024_6);

wire[3:0] wires_1025_6;

wire[31:0] addr_1025_6;

Selector_2 s1025_6(wires_256_5[1], addr_256_5, wires_1025_6,addr_1025_6);

wire[3:0] wires_1026_6;

wire[31:0] addr_1026_6;

Selector_2 s1026_6(wires_256_5[2], addr_256_5, wires_1026_6,addr_1026_6);

wire[3:0] wires_1027_6;

wire[31:0] addr_1027_6;

Selector_2 s1027_6(wires_256_5[3], addr_256_5, wires_1027_6,addr_1027_6);

wire[3:0] wires_1028_6;

wire[31:0] addr_1028_6;

Selector_2 s1028_6(wires_257_5[0], addr_257_5, wires_1028_6,addr_1028_6);

wire[3:0] wires_1029_6;

wire[31:0] addr_1029_6;

Selector_2 s1029_6(wires_257_5[1], addr_257_5, wires_1029_6,addr_1029_6);

wire[3:0] wires_1030_6;

wire[31:0] addr_1030_6;

Selector_2 s1030_6(wires_257_5[2], addr_257_5, wires_1030_6,addr_1030_6);

wire[3:0] wires_1031_6;

wire[31:0] addr_1031_6;

Selector_2 s1031_6(wires_257_5[3], addr_257_5, wires_1031_6,addr_1031_6);

wire[3:0] wires_1032_6;

wire[31:0] addr_1032_6;

Selector_2 s1032_6(wires_258_5[0], addr_258_5, wires_1032_6,addr_1032_6);

wire[3:0] wires_1033_6;

wire[31:0] addr_1033_6;

Selector_2 s1033_6(wires_258_5[1], addr_258_5, wires_1033_6,addr_1033_6);

wire[3:0] wires_1034_6;

wire[31:0] addr_1034_6;

Selector_2 s1034_6(wires_258_5[2], addr_258_5, wires_1034_6,addr_1034_6);

wire[3:0] wires_1035_6;

wire[31:0] addr_1035_6;

Selector_2 s1035_6(wires_258_5[3], addr_258_5, wires_1035_6,addr_1035_6);

wire[3:0] wires_1036_6;

wire[31:0] addr_1036_6;

Selector_2 s1036_6(wires_259_5[0], addr_259_5, wires_1036_6,addr_1036_6);

wire[3:0] wires_1037_6;

wire[31:0] addr_1037_6;

Selector_2 s1037_6(wires_259_5[1], addr_259_5, wires_1037_6,addr_1037_6);

wire[3:0] wires_1038_6;

wire[31:0] addr_1038_6;

Selector_2 s1038_6(wires_259_5[2], addr_259_5, wires_1038_6,addr_1038_6);

wire[3:0] wires_1039_6;

wire[31:0] addr_1039_6;

Selector_2 s1039_6(wires_259_5[3], addr_259_5, wires_1039_6,addr_1039_6);

wire[3:0] wires_1040_6;

wire[31:0] addr_1040_6;

Selector_2 s1040_6(wires_260_5[0], addr_260_5, wires_1040_6,addr_1040_6);

wire[3:0] wires_1041_6;

wire[31:0] addr_1041_6;

Selector_2 s1041_6(wires_260_5[1], addr_260_5, wires_1041_6,addr_1041_6);

wire[3:0] wires_1042_6;

wire[31:0] addr_1042_6;

Selector_2 s1042_6(wires_260_5[2], addr_260_5, wires_1042_6,addr_1042_6);

wire[3:0] wires_1043_6;

wire[31:0] addr_1043_6;

Selector_2 s1043_6(wires_260_5[3], addr_260_5, wires_1043_6,addr_1043_6);

wire[3:0] wires_1044_6;

wire[31:0] addr_1044_6;

Selector_2 s1044_6(wires_261_5[0], addr_261_5, wires_1044_6,addr_1044_6);

wire[3:0] wires_1045_6;

wire[31:0] addr_1045_6;

Selector_2 s1045_6(wires_261_5[1], addr_261_5, wires_1045_6,addr_1045_6);

wire[3:0] wires_1046_6;

wire[31:0] addr_1046_6;

Selector_2 s1046_6(wires_261_5[2], addr_261_5, wires_1046_6,addr_1046_6);

wire[3:0] wires_1047_6;

wire[31:0] addr_1047_6;

Selector_2 s1047_6(wires_261_5[3], addr_261_5, wires_1047_6,addr_1047_6);

wire[3:0] wires_1048_6;

wire[31:0] addr_1048_6;

Selector_2 s1048_6(wires_262_5[0], addr_262_5, wires_1048_6,addr_1048_6);

wire[3:0] wires_1049_6;

wire[31:0] addr_1049_6;

Selector_2 s1049_6(wires_262_5[1], addr_262_5, wires_1049_6,addr_1049_6);

wire[3:0] wires_1050_6;

wire[31:0] addr_1050_6;

Selector_2 s1050_6(wires_262_5[2], addr_262_5, wires_1050_6,addr_1050_6);

wire[3:0] wires_1051_6;

wire[31:0] addr_1051_6;

Selector_2 s1051_6(wires_262_5[3], addr_262_5, wires_1051_6,addr_1051_6);

wire[3:0] wires_1052_6;

wire[31:0] addr_1052_6;

Selector_2 s1052_6(wires_263_5[0], addr_263_5, wires_1052_6,addr_1052_6);

wire[3:0] wires_1053_6;

wire[31:0] addr_1053_6;

Selector_2 s1053_6(wires_263_5[1], addr_263_5, wires_1053_6,addr_1053_6);

wire[3:0] wires_1054_6;

wire[31:0] addr_1054_6;

Selector_2 s1054_6(wires_263_5[2], addr_263_5, wires_1054_6,addr_1054_6);

wire[3:0] wires_1055_6;

wire[31:0] addr_1055_6;

Selector_2 s1055_6(wires_263_5[3], addr_263_5, wires_1055_6,addr_1055_6);

wire[3:0] wires_1056_6;

wire[31:0] addr_1056_6;

Selector_2 s1056_6(wires_264_5[0], addr_264_5, wires_1056_6,addr_1056_6);

wire[3:0] wires_1057_6;

wire[31:0] addr_1057_6;

Selector_2 s1057_6(wires_264_5[1], addr_264_5, wires_1057_6,addr_1057_6);

wire[3:0] wires_1058_6;

wire[31:0] addr_1058_6;

Selector_2 s1058_6(wires_264_5[2], addr_264_5, wires_1058_6,addr_1058_6);

wire[3:0] wires_1059_6;

wire[31:0] addr_1059_6;

Selector_2 s1059_6(wires_264_5[3], addr_264_5, wires_1059_6,addr_1059_6);

wire[3:0] wires_1060_6;

wire[31:0] addr_1060_6;

Selector_2 s1060_6(wires_265_5[0], addr_265_5, wires_1060_6,addr_1060_6);

wire[3:0] wires_1061_6;

wire[31:0] addr_1061_6;

Selector_2 s1061_6(wires_265_5[1], addr_265_5, wires_1061_6,addr_1061_6);

wire[3:0] wires_1062_6;

wire[31:0] addr_1062_6;

Selector_2 s1062_6(wires_265_5[2], addr_265_5, wires_1062_6,addr_1062_6);

wire[3:0] wires_1063_6;

wire[31:0] addr_1063_6;

Selector_2 s1063_6(wires_265_5[3], addr_265_5, wires_1063_6,addr_1063_6);

wire[3:0] wires_1064_6;

wire[31:0] addr_1064_6;

Selector_2 s1064_6(wires_266_5[0], addr_266_5, wires_1064_6,addr_1064_6);

wire[3:0] wires_1065_6;

wire[31:0] addr_1065_6;

Selector_2 s1065_6(wires_266_5[1], addr_266_5, wires_1065_6,addr_1065_6);

wire[3:0] wires_1066_6;

wire[31:0] addr_1066_6;

Selector_2 s1066_6(wires_266_5[2], addr_266_5, wires_1066_6,addr_1066_6);

wire[3:0] wires_1067_6;

wire[31:0] addr_1067_6;

Selector_2 s1067_6(wires_266_5[3], addr_266_5, wires_1067_6,addr_1067_6);

wire[3:0] wires_1068_6;

wire[31:0] addr_1068_6;

Selector_2 s1068_6(wires_267_5[0], addr_267_5, wires_1068_6,addr_1068_6);

wire[3:0] wires_1069_6;

wire[31:0] addr_1069_6;

Selector_2 s1069_6(wires_267_5[1], addr_267_5, wires_1069_6,addr_1069_6);

wire[3:0] wires_1070_6;

wire[31:0] addr_1070_6;

Selector_2 s1070_6(wires_267_5[2], addr_267_5, wires_1070_6,addr_1070_6);

wire[3:0] wires_1071_6;

wire[31:0] addr_1071_6;

Selector_2 s1071_6(wires_267_5[3], addr_267_5, wires_1071_6,addr_1071_6);

wire[3:0] wires_1072_6;

wire[31:0] addr_1072_6;

Selector_2 s1072_6(wires_268_5[0], addr_268_5, wires_1072_6,addr_1072_6);

wire[3:0] wires_1073_6;

wire[31:0] addr_1073_6;

Selector_2 s1073_6(wires_268_5[1], addr_268_5, wires_1073_6,addr_1073_6);

wire[3:0] wires_1074_6;

wire[31:0] addr_1074_6;

Selector_2 s1074_6(wires_268_5[2], addr_268_5, wires_1074_6,addr_1074_6);

wire[3:0] wires_1075_6;

wire[31:0] addr_1075_6;

Selector_2 s1075_6(wires_268_5[3], addr_268_5, wires_1075_6,addr_1075_6);

wire[3:0] wires_1076_6;

wire[31:0] addr_1076_6;

Selector_2 s1076_6(wires_269_5[0], addr_269_5, wires_1076_6,addr_1076_6);

wire[3:0] wires_1077_6;

wire[31:0] addr_1077_6;

Selector_2 s1077_6(wires_269_5[1], addr_269_5, wires_1077_6,addr_1077_6);

wire[3:0] wires_1078_6;

wire[31:0] addr_1078_6;

Selector_2 s1078_6(wires_269_5[2], addr_269_5, wires_1078_6,addr_1078_6);

wire[3:0] wires_1079_6;

wire[31:0] addr_1079_6;

Selector_2 s1079_6(wires_269_5[3], addr_269_5, wires_1079_6,addr_1079_6);

wire[3:0] wires_1080_6;

wire[31:0] addr_1080_6;

Selector_2 s1080_6(wires_270_5[0], addr_270_5, wires_1080_6,addr_1080_6);

wire[3:0] wires_1081_6;

wire[31:0] addr_1081_6;

Selector_2 s1081_6(wires_270_5[1], addr_270_5, wires_1081_6,addr_1081_6);

wire[3:0] wires_1082_6;

wire[31:0] addr_1082_6;

Selector_2 s1082_6(wires_270_5[2], addr_270_5, wires_1082_6,addr_1082_6);

wire[3:0] wires_1083_6;

wire[31:0] addr_1083_6;

Selector_2 s1083_6(wires_270_5[3], addr_270_5, wires_1083_6,addr_1083_6);

wire[3:0] wires_1084_6;

wire[31:0] addr_1084_6;

Selector_2 s1084_6(wires_271_5[0], addr_271_5, wires_1084_6,addr_1084_6);

wire[3:0] wires_1085_6;

wire[31:0] addr_1085_6;

Selector_2 s1085_6(wires_271_5[1], addr_271_5, wires_1085_6,addr_1085_6);

wire[3:0] wires_1086_6;

wire[31:0] addr_1086_6;

Selector_2 s1086_6(wires_271_5[2], addr_271_5, wires_1086_6,addr_1086_6);

wire[3:0] wires_1087_6;

wire[31:0] addr_1087_6;

Selector_2 s1087_6(wires_271_5[3], addr_271_5, wires_1087_6,addr_1087_6);

wire[3:0] wires_1088_6;

wire[31:0] addr_1088_6;

Selector_2 s1088_6(wires_272_5[0], addr_272_5, wires_1088_6,addr_1088_6);

wire[3:0] wires_1089_6;

wire[31:0] addr_1089_6;

Selector_2 s1089_6(wires_272_5[1], addr_272_5, wires_1089_6,addr_1089_6);

wire[3:0] wires_1090_6;

wire[31:0] addr_1090_6;

Selector_2 s1090_6(wires_272_5[2], addr_272_5, wires_1090_6,addr_1090_6);

wire[3:0] wires_1091_6;

wire[31:0] addr_1091_6;

Selector_2 s1091_6(wires_272_5[3], addr_272_5, wires_1091_6,addr_1091_6);

wire[3:0] wires_1092_6;

wire[31:0] addr_1092_6;

Selector_2 s1092_6(wires_273_5[0], addr_273_5, wires_1092_6,addr_1092_6);

wire[3:0] wires_1093_6;

wire[31:0] addr_1093_6;

Selector_2 s1093_6(wires_273_5[1], addr_273_5, wires_1093_6,addr_1093_6);

wire[3:0] wires_1094_6;

wire[31:0] addr_1094_6;

Selector_2 s1094_6(wires_273_5[2], addr_273_5, wires_1094_6,addr_1094_6);

wire[3:0] wires_1095_6;

wire[31:0] addr_1095_6;

Selector_2 s1095_6(wires_273_5[3], addr_273_5, wires_1095_6,addr_1095_6);

wire[3:0] wires_1096_6;

wire[31:0] addr_1096_6;

Selector_2 s1096_6(wires_274_5[0], addr_274_5, wires_1096_6,addr_1096_6);

wire[3:0] wires_1097_6;

wire[31:0] addr_1097_6;

Selector_2 s1097_6(wires_274_5[1], addr_274_5, wires_1097_6,addr_1097_6);

wire[3:0] wires_1098_6;

wire[31:0] addr_1098_6;

Selector_2 s1098_6(wires_274_5[2], addr_274_5, wires_1098_6,addr_1098_6);

wire[3:0] wires_1099_6;

wire[31:0] addr_1099_6;

Selector_2 s1099_6(wires_274_5[3], addr_274_5, wires_1099_6,addr_1099_6);

wire[3:0] wires_1100_6;

wire[31:0] addr_1100_6;

Selector_2 s1100_6(wires_275_5[0], addr_275_5, wires_1100_6,addr_1100_6);

wire[3:0] wires_1101_6;

wire[31:0] addr_1101_6;

Selector_2 s1101_6(wires_275_5[1], addr_275_5, wires_1101_6,addr_1101_6);

wire[3:0] wires_1102_6;

wire[31:0] addr_1102_6;

Selector_2 s1102_6(wires_275_5[2], addr_275_5, wires_1102_6,addr_1102_6);

wire[3:0] wires_1103_6;

wire[31:0] addr_1103_6;

Selector_2 s1103_6(wires_275_5[3], addr_275_5, wires_1103_6,addr_1103_6);

wire[3:0] wires_1104_6;

wire[31:0] addr_1104_6;

Selector_2 s1104_6(wires_276_5[0], addr_276_5, wires_1104_6,addr_1104_6);

wire[3:0] wires_1105_6;

wire[31:0] addr_1105_6;

Selector_2 s1105_6(wires_276_5[1], addr_276_5, wires_1105_6,addr_1105_6);

wire[3:0] wires_1106_6;

wire[31:0] addr_1106_6;

Selector_2 s1106_6(wires_276_5[2], addr_276_5, wires_1106_6,addr_1106_6);

wire[3:0] wires_1107_6;

wire[31:0] addr_1107_6;

Selector_2 s1107_6(wires_276_5[3], addr_276_5, wires_1107_6,addr_1107_6);

wire[3:0] wires_1108_6;

wire[31:0] addr_1108_6;

Selector_2 s1108_6(wires_277_5[0], addr_277_5, wires_1108_6,addr_1108_6);

wire[3:0] wires_1109_6;

wire[31:0] addr_1109_6;

Selector_2 s1109_6(wires_277_5[1], addr_277_5, wires_1109_6,addr_1109_6);

wire[3:0] wires_1110_6;

wire[31:0] addr_1110_6;

Selector_2 s1110_6(wires_277_5[2], addr_277_5, wires_1110_6,addr_1110_6);

wire[3:0] wires_1111_6;

wire[31:0] addr_1111_6;

Selector_2 s1111_6(wires_277_5[3], addr_277_5, wires_1111_6,addr_1111_6);

wire[3:0] wires_1112_6;

wire[31:0] addr_1112_6;

Selector_2 s1112_6(wires_278_5[0], addr_278_5, wires_1112_6,addr_1112_6);

wire[3:0] wires_1113_6;

wire[31:0] addr_1113_6;

Selector_2 s1113_6(wires_278_5[1], addr_278_5, wires_1113_6,addr_1113_6);

wire[3:0] wires_1114_6;

wire[31:0] addr_1114_6;

Selector_2 s1114_6(wires_278_5[2], addr_278_5, wires_1114_6,addr_1114_6);

wire[3:0] wires_1115_6;

wire[31:0] addr_1115_6;

Selector_2 s1115_6(wires_278_5[3], addr_278_5, wires_1115_6,addr_1115_6);

wire[3:0] wires_1116_6;

wire[31:0] addr_1116_6;

Selector_2 s1116_6(wires_279_5[0], addr_279_5, wires_1116_6,addr_1116_6);

wire[3:0] wires_1117_6;

wire[31:0] addr_1117_6;

Selector_2 s1117_6(wires_279_5[1], addr_279_5, wires_1117_6,addr_1117_6);

wire[3:0] wires_1118_6;

wire[31:0] addr_1118_6;

Selector_2 s1118_6(wires_279_5[2], addr_279_5, wires_1118_6,addr_1118_6);

wire[3:0] wires_1119_6;

wire[31:0] addr_1119_6;

Selector_2 s1119_6(wires_279_5[3], addr_279_5, wires_1119_6,addr_1119_6);

wire[3:0] wires_1120_6;

wire[31:0] addr_1120_6;

Selector_2 s1120_6(wires_280_5[0], addr_280_5, wires_1120_6,addr_1120_6);

wire[3:0] wires_1121_6;

wire[31:0] addr_1121_6;

Selector_2 s1121_6(wires_280_5[1], addr_280_5, wires_1121_6,addr_1121_6);

wire[3:0] wires_1122_6;

wire[31:0] addr_1122_6;

Selector_2 s1122_6(wires_280_5[2], addr_280_5, wires_1122_6,addr_1122_6);

wire[3:0] wires_1123_6;

wire[31:0] addr_1123_6;

Selector_2 s1123_6(wires_280_5[3], addr_280_5, wires_1123_6,addr_1123_6);

wire[3:0] wires_1124_6;

wire[31:0] addr_1124_6;

Selector_2 s1124_6(wires_281_5[0], addr_281_5, wires_1124_6,addr_1124_6);

wire[3:0] wires_1125_6;

wire[31:0] addr_1125_6;

Selector_2 s1125_6(wires_281_5[1], addr_281_5, wires_1125_6,addr_1125_6);

wire[3:0] wires_1126_6;

wire[31:0] addr_1126_6;

Selector_2 s1126_6(wires_281_5[2], addr_281_5, wires_1126_6,addr_1126_6);

wire[3:0] wires_1127_6;

wire[31:0] addr_1127_6;

Selector_2 s1127_6(wires_281_5[3], addr_281_5, wires_1127_6,addr_1127_6);

wire[3:0] wires_1128_6;

wire[31:0] addr_1128_6;

Selector_2 s1128_6(wires_282_5[0], addr_282_5, wires_1128_6,addr_1128_6);

wire[3:0] wires_1129_6;

wire[31:0] addr_1129_6;

Selector_2 s1129_6(wires_282_5[1], addr_282_5, wires_1129_6,addr_1129_6);

wire[3:0] wires_1130_6;

wire[31:0] addr_1130_6;

Selector_2 s1130_6(wires_282_5[2], addr_282_5, wires_1130_6,addr_1130_6);

wire[3:0] wires_1131_6;

wire[31:0] addr_1131_6;

Selector_2 s1131_6(wires_282_5[3], addr_282_5, wires_1131_6,addr_1131_6);

wire[3:0] wires_1132_6;

wire[31:0] addr_1132_6;

Selector_2 s1132_6(wires_283_5[0], addr_283_5, wires_1132_6,addr_1132_6);

wire[3:0] wires_1133_6;

wire[31:0] addr_1133_6;

Selector_2 s1133_6(wires_283_5[1], addr_283_5, wires_1133_6,addr_1133_6);

wire[3:0] wires_1134_6;

wire[31:0] addr_1134_6;

Selector_2 s1134_6(wires_283_5[2], addr_283_5, wires_1134_6,addr_1134_6);

wire[3:0] wires_1135_6;

wire[31:0] addr_1135_6;

Selector_2 s1135_6(wires_283_5[3], addr_283_5, wires_1135_6,addr_1135_6);

wire[3:0] wires_1136_6;

wire[31:0] addr_1136_6;

Selector_2 s1136_6(wires_284_5[0], addr_284_5, wires_1136_6,addr_1136_6);

wire[3:0] wires_1137_6;

wire[31:0] addr_1137_6;

Selector_2 s1137_6(wires_284_5[1], addr_284_5, wires_1137_6,addr_1137_6);

wire[3:0] wires_1138_6;

wire[31:0] addr_1138_6;

Selector_2 s1138_6(wires_284_5[2], addr_284_5, wires_1138_6,addr_1138_6);

wire[3:0] wires_1139_6;

wire[31:0] addr_1139_6;

Selector_2 s1139_6(wires_284_5[3], addr_284_5, wires_1139_6,addr_1139_6);

wire[3:0] wires_1140_6;

wire[31:0] addr_1140_6;

Selector_2 s1140_6(wires_285_5[0], addr_285_5, wires_1140_6,addr_1140_6);

wire[3:0] wires_1141_6;

wire[31:0] addr_1141_6;

Selector_2 s1141_6(wires_285_5[1], addr_285_5, wires_1141_6,addr_1141_6);

wire[3:0] wires_1142_6;

wire[31:0] addr_1142_6;

Selector_2 s1142_6(wires_285_5[2], addr_285_5, wires_1142_6,addr_1142_6);

wire[3:0] wires_1143_6;

wire[31:0] addr_1143_6;

Selector_2 s1143_6(wires_285_5[3], addr_285_5, wires_1143_6,addr_1143_6);

wire[3:0] wires_1144_6;

wire[31:0] addr_1144_6;

Selector_2 s1144_6(wires_286_5[0], addr_286_5, wires_1144_6,addr_1144_6);

wire[3:0] wires_1145_6;

wire[31:0] addr_1145_6;

Selector_2 s1145_6(wires_286_5[1], addr_286_5, wires_1145_6,addr_1145_6);

wire[3:0] wires_1146_6;

wire[31:0] addr_1146_6;

Selector_2 s1146_6(wires_286_5[2], addr_286_5, wires_1146_6,addr_1146_6);

wire[3:0] wires_1147_6;

wire[31:0] addr_1147_6;

Selector_2 s1147_6(wires_286_5[3], addr_286_5, wires_1147_6,addr_1147_6);

wire[3:0] wires_1148_6;

wire[31:0] addr_1148_6;

Selector_2 s1148_6(wires_287_5[0], addr_287_5, wires_1148_6,addr_1148_6);

wire[3:0] wires_1149_6;

wire[31:0] addr_1149_6;

Selector_2 s1149_6(wires_287_5[1], addr_287_5, wires_1149_6,addr_1149_6);

wire[3:0] wires_1150_6;

wire[31:0] addr_1150_6;

Selector_2 s1150_6(wires_287_5[2], addr_287_5, wires_1150_6,addr_1150_6);

wire[3:0] wires_1151_6;

wire[31:0] addr_1151_6;

Selector_2 s1151_6(wires_287_5[3], addr_287_5, wires_1151_6,addr_1151_6);

wire[3:0] wires_1152_6;

wire[31:0] addr_1152_6;

Selector_2 s1152_6(wires_288_5[0], addr_288_5, wires_1152_6,addr_1152_6);

wire[3:0] wires_1153_6;

wire[31:0] addr_1153_6;

Selector_2 s1153_6(wires_288_5[1], addr_288_5, wires_1153_6,addr_1153_6);

wire[3:0] wires_1154_6;

wire[31:0] addr_1154_6;

Selector_2 s1154_6(wires_288_5[2], addr_288_5, wires_1154_6,addr_1154_6);

wire[3:0] wires_1155_6;

wire[31:0] addr_1155_6;

Selector_2 s1155_6(wires_288_5[3], addr_288_5, wires_1155_6,addr_1155_6);

wire[3:0] wires_1156_6;

wire[31:0] addr_1156_6;

Selector_2 s1156_6(wires_289_5[0], addr_289_5, wires_1156_6,addr_1156_6);

wire[3:0] wires_1157_6;

wire[31:0] addr_1157_6;

Selector_2 s1157_6(wires_289_5[1], addr_289_5, wires_1157_6,addr_1157_6);

wire[3:0] wires_1158_6;

wire[31:0] addr_1158_6;

Selector_2 s1158_6(wires_289_5[2], addr_289_5, wires_1158_6,addr_1158_6);

wire[3:0] wires_1159_6;

wire[31:0] addr_1159_6;

Selector_2 s1159_6(wires_289_5[3], addr_289_5, wires_1159_6,addr_1159_6);

wire[3:0] wires_1160_6;

wire[31:0] addr_1160_6;

Selector_2 s1160_6(wires_290_5[0], addr_290_5, wires_1160_6,addr_1160_6);

wire[3:0] wires_1161_6;

wire[31:0] addr_1161_6;

Selector_2 s1161_6(wires_290_5[1], addr_290_5, wires_1161_6,addr_1161_6);

wire[3:0] wires_1162_6;

wire[31:0] addr_1162_6;

Selector_2 s1162_6(wires_290_5[2], addr_290_5, wires_1162_6,addr_1162_6);

wire[3:0] wires_1163_6;

wire[31:0] addr_1163_6;

Selector_2 s1163_6(wires_290_5[3], addr_290_5, wires_1163_6,addr_1163_6);

wire[3:0] wires_1164_6;

wire[31:0] addr_1164_6;

Selector_2 s1164_6(wires_291_5[0], addr_291_5, wires_1164_6,addr_1164_6);

wire[3:0] wires_1165_6;

wire[31:0] addr_1165_6;

Selector_2 s1165_6(wires_291_5[1], addr_291_5, wires_1165_6,addr_1165_6);

wire[3:0] wires_1166_6;

wire[31:0] addr_1166_6;

Selector_2 s1166_6(wires_291_5[2], addr_291_5, wires_1166_6,addr_1166_6);

wire[3:0] wires_1167_6;

wire[31:0] addr_1167_6;

Selector_2 s1167_6(wires_291_5[3], addr_291_5, wires_1167_6,addr_1167_6);

wire[3:0] wires_1168_6;

wire[31:0] addr_1168_6;

Selector_2 s1168_6(wires_292_5[0], addr_292_5, wires_1168_6,addr_1168_6);

wire[3:0] wires_1169_6;

wire[31:0] addr_1169_6;

Selector_2 s1169_6(wires_292_5[1], addr_292_5, wires_1169_6,addr_1169_6);

wire[3:0] wires_1170_6;

wire[31:0] addr_1170_6;

Selector_2 s1170_6(wires_292_5[2], addr_292_5, wires_1170_6,addr_1170_6);

wire[3:0] wires_1171_6;

wire[31:0] addr_1171_6;

Selector_2 s1171_6(wires_292_5[3], addr_292_5, wires_1171_6,addr_1171_6);

wire[3:0] wires_1172_6;

wire[31:0] addr_1172_6;

Selector_2 s1172_6(wires_293_5[0], addr_293_5, wires_1172_6,addr_1172_6);

wire[3:0] wires_1173_6;

wire[31:0] addr_1173_6;

Selector_2 s1173_6(wires_293_5[1], addr_293_5, wires_1173_6,addr_1173_6);

wire[3:0] wires_1174_6;

wire[31:0] addr_1174_6;

Selector_2 s1174_6(wires_293_5[2], addr_293_5, wires_1174_6,addr_1174_6);

wire[3:0] wires_1175_6;

wire[31:0] addr_1175_6;

Selector_2 s1175_6(wires_293_5[3], addr_293_5, wires_1175_6,addr_1175_6);

wire[3:0] wires_1176_6;

wire[31:0] addr_1176_6;

Selector_2 s1176_6(wires_294_5[0], addr_294_5, wires_1176_6,addr_1176_6);

wire[3:0] wires_1177_6;

wire[31:0] addr_1177_6;

Selector_2 s1177_6(wires_294_5[1], addr_294_5, wires_1177_6,addr_1177_6);

wire[3:0] wires_1178_6;

wire[31:0] addr_1178_6;

Selector_2 s1178_6(wires_294_5[2], addr_294_5, wires_1178_6,addr_1178_6);

wire[3:0] wires_1179_6;

wire[31:0] addr_1179_6;

Selector_2 s1179_6(wires_294_5[3], addr_294_5, wires_1179_6,addr_1179_6);

wire[3:0] wires_1180_6;

wire[31:0] addr_1180_6;

Selector_2 s1180_6(wires_295_5[0], addr_295_5, wires_1180_6,addr_1180_6);

wire[3:0] wires_1181_6;

wire[31:0] addr_1181_6;

Selector_2 s1181_6(wires_295_5[1], addr_295_5, wires_1181_6,addr_1181_6);

wire[3:0] wires_1182_6;

wire[31:0] addr_1182_6;

Selector_2 s1182_6(wires_295_5[2], addr_295_5, wires_1182_6,addr_1182_6);

wire[3:0] wires_1183_6;

wire[31:0] addr_1183_6;

Selector_2 s1183_6(wires_295_5[3], addr_295_5, wires_1183_6,addr_1183_6);

wire[3:0] wires_1184_6;

wire[31:0] addr_1184_6;

Selector_2 s1184_6(wires_296_5[0], addr_296_5, wires_1184_6,addr_1184_6);

wire[3:0] wires_1185_6;

wire[31:0] addr_1185_6;

Selector_2 s1185_6(wires_296_5[1], addr_296_5, wires_1185_6,addr_1185_6);

wire[3:0] wires_1186_6;

wire[31:0] addr_1186_6;

Selector_2 s1186_6(wires_296_5[2], addr_296_5, wires_1186_6,addr_1186_6);

wire[3:0] wires_1187_6;

wire[31:0] addr_1187_6;

Selector_2 s1187_6(wires_296_5[3], addr_296_5, wires_1187_6,addr_1187_6);

wire[3:0] wires_1188_6;

wire[31:0] addr_1188_6;

Selector_2 s1188_6(wires_297_5[0], addr_297_5, wires_1188_6,addr_1188_6);

wire[3:0] wires_1189_6;

wire[31:0] addr_1189_6;

Selector_2 s1189_6(wires_297_5[1], addr_297_5, wires_1189_6,addr_1189_6);

wire[3:0] wires_1190_6;

wire[31:0] addr_1190_6;

Selector_2 s1190_6(wires_297_5[2], addr_297_5, wires_1190_6,addr_1190_6);

wire[3:0] wires_1191_6;

wire[31:0] addr_1191_6;

Selector_2 s1191_6(wires_297_5[3], addr_297_5, wires_1191_6,addr_1191_6);

wire[3:0] wires_1192_6;

wire[31:0] addr_1192_6;

Selector_2 s1192_6(wires_298_5[0], addr_298_5, wires_1192_6,addr_1192_6);

wire[3:0] wires_1193_6;

wire[31:0] addr_1193_6;

Selector_2 s1193_6(wires_298_5[1], addr_298_5, wires_1193_6,addr_1193_6);

wire[3:0] wires_1194_6;

wire[31:0] addr_1194_6;

Selector_2 s1194_6(wires_298_5[2], addr_298_5, wires_1194_6,addr_1194_6);

wire[3:0] wires_1195_6;

wire[31:0] addr_1195_6;

Selector_2 s1195_6(wires_298_5[3], addr_298_5, wires_1195_6,addr_1195_6);

wire[3:0] wires_1196_6;

wire[31:0] addr_1196_6;

Selector_2 s1196_6(wires_299_5[0], addr_299_5, wires_1196_6,addr_1196_6);

wire[3:0] wires_1197_6;

wire[31:0] addr_1197_6;

Selector_2 s1197_6(wires_299_5[1], addr_299_5, wires_1197_6,addr_1197_6);

wire[3:0] wires_1198_6;

wire[31:0] addr_1198_6;

Selector_2 s1198_6(wires_299_5[2], addr_299_5, wires_1198_6,addr_1198_6);

wire[3:0] wires_1199_6;

wire[31:0] addr_1199_6;

Selector_2 s1199_6(wires_299_5[3], addr_299_5, wires_1199_6,addr_1199_6);

wire[3:0] wires_1200_6;

wire[31:0] addr_1200_6;

Selector_2 s1200_6(wires_300_5[0], addr_300_5, wires_1200_6,addr_1200_6);

wire[3:0] wires_1201_6;

wire[31:0] addr_1201_6;

Selector_2 s1201_6(wires_300_5[1], addr_300_5, wires_1201_6,addr_1201_6);

wire[3:0] wires_1202_6;

wire[31:0] addr_1202_6;

Selector_2 s1202_6(wires_300_5[2], addr_300_5, wires_1202_6,addr_1202_6);

wire[3:0] wires_1203_6;

wire[31:0] addr_1203_6;

Selector_2 s1203_6(wires_300_5[3], addr_300_5, wires_1203_6,addr_1203_6);

wire[3:0] wires_1204_6;

wire[31:0] addr_1204_6;

Selector_2 s1204_6(wires_301_5[0], addr_301_5, wires_1204_6,addr_1204_6);

wire[3:0] wires_1205_6;

wire[31:0] addr_1205_6;

Selector_2 s1205_6(wires_301_5[1], addr_301_5, wires_1205_6,addr_1205_6);

wire[3:0] wires_1206_6;

wire[31:0] addr_1206_6;

Selector_2 s1206_6(wires_301_5[2], addr_301_5, wires_1206_6,addr_1206_6);

wire[3:0] wires_1207_6;

wire[31:0] addr_1207_6;

Selector_2 s1207_6(wires_301_5[3], addr_301_5, wires_1207_6,addr_1207_6);

wire[3:0] wires_1208_6;

wire[31:0] addr_1208_6;

Selector_2 s1208_6(wires_302_5[0], addr_302_5, wires_1208_6,addr_1208_6);

wire[3:0] wires_1209_6;

wire[31:0] addr_1209_6;

Selector_2 s1209_6(wires_302_5[1], addr_302_5, wires_1209_6,addr_1209_6);

wire[3:0] wires_1210_6;

wire[31:0] addr_1210_6;

Selector_2 s1210_6(wires_302_5[2], addr_302_5, wires_1210_6,addr_1210_6);

wire[3:0] wires_1211_6;

wire[31:0] addr_1211_6;

Selector_2 s1211_6(wires_302_5[3], addr_302_5, wires_1211_6,addr_1211_6);

wire[3:0] wires_1212_6;

wire[31:0] addr_1212_6;

Selector_2 s1212_6(wires_303_5[0], addr_303_5, wires_1212_6,addr_1212_6);

wire[3:0] wires_1213_6;

wire[31:0] addr_1213_6;

Selector_2 s1213_6(wires_303_5[1], addr_303_5, wires_1213_6,addr_1213_6);

wire[3:0] wires_1214_6;

wire[31:0] addr_1214_6;

Selector_2 s1214_6(wires_303_5[2], addr_303_5, wires_1214_6,addr_1214_6);

wire[3:0] wires_1215_6;

wire[31:0] addr_1215_6;

Selector_2 s1215_6(wires_303_5[3], addr_303_5, wires_1215_6,addr_1215_6);

wire[3:0] wires_1216_6;

wire[31:0] addr_1216_6;

Selector_2 s1216_6(wires_304_5[0], addr_304_5, wires_1216_6,addr_1216_6);

wire[3:0] wires_1217_6;

wire[31:0] addr_1217_6;

Selector_2 s1217_6(wires_304_5[1], addr_304_5, wires_1217_6,addr_1217_6);

wire[3:0] wires_1218_6;

wire[31:0] addr_1218_6;

Selector_2 s1218_6(wires_304_5[2], addr_304_5, wires_1218_6,addr_1218_6);

wire[3:0] wires_1219_6;

wire[31:0] addr_1219_6;

Selector_2 s1219_6(wires_304_5[3], addr_304_5, wires_1219_6,addr_1219_6);

wire[3:0] wires_1220_6;

wire[31:0] addr_1220_6;

Selector_2 s1220_6(wires_305_5[0], addr_305_5, wires_1220_6,addr_1220_6);

wire[3:0] wires_1221_6;

wire[31:0] addr_1221_6;

Selector_2 s1221_6(wires_305_5[1], addr_305_5, wires_1221_6,addr_1221_6);

wire[3:0] wires_1222_6;

wire[31:0] addr_1222_6;

Selector_2 s1222_6(wires_305_5[2], addr_305_5, wires_1222_6,addr_1222_6);

wire[3:0] wires_1223_6;

wire[31:0] addr_1223_6;

Selector_2 s1223_6(wires_305_5[3], addr_305_5, wires_1223_6,addr_1223_6);

wire[3:0] wires_1224_6;

wire[31:0] addr_1224_6;

Selector_2 s1224_6(wires_306_5[0], addr_306_5, wires_1224_6,addr_1224_6);

wire[3:0] wires_1225_6;

wire[31:0] addr_1225_6;

Selector_2 s1225_6(wires_306_5[1], addr_306_5, wires_1225_6,addr_1225_6);

wire[3:0] wires_1226_6;

wire[31:0] addr_1226_6;

Selector_2 s1226_6(wires_306_5[2], addr_306_5, wires_1226_6,addr_1226_6);

wire[3:0] wires_1227_6;

wire[31:0] addr_1227_6;

Selector_2 s1227_6(wires_306_5[3], addr_306_5, wires_1227_6,addr_1227_6);

wire[3:0] wires_1228_6;

wire[31:0] addr_1228_6;

Selector_2 s1228_6(wires_307_5[0], addr_307_5, wires_1228_6,addr_1228_6);

wire[3:0] wires_1229_6;

wire[31:0] addr_1229_6;

Selector_2 s1229_6(wires_307_5[1], addr_307_5, wires_1229_6,addr_1229_6);

wire[3:0] wires_1230_6;

wire[31:0] addr_1230_6;

Selector_2 s1230_6(wires_307_5[2], addr_307_5, wires_1230_6,addr_1230_6);

wire[3:0] wires_1231_6;

wire[31:0] addr_1231_6;

Selector_2 s1231_6(wires_307_5[3], addr_307_5, wires_1231_6,addr_1231_6);

wire[3:0] wires_1232_6;

wire[31:0] addr_1232_6;

Selector_2 s1232_6(wires_308_5[0], addr_308_5, wires_1232_6,addr_1232_6);

wire[3:0] wires_1233_6;

wire[31:0] addr_1233_6;

Selector_2 s1233_6(wires_308_5[1], addr_308_5, wires_1233_6,addr_1233_6);

wire[3:0] wires_1234_6;

wire[31:0] addr_1234_6;

Selector_2 s1234_6(wires_308_5[2], addr_308_5, wires_1234_6,addr_1234_6);

wire[3:0] wires_1235_6;

wire[31:0] addr_1235_6;

Selector_2 s1235_6(wires_308_5[3], addr_308_5, wires_1235_6,addr_1235_6);

wire[3:0] wires_1236_6;

wire[31:0] addr_1236_6;

Selector_2 s1236_6(wires_309_5[0], addr_309_5, wires_1236_6,addr_1236_6);

wire[3:0] wires_1237_6;

wire[31:0] addr_1237_6;

Selector_2 s1237_6(wires_309_5[1], addr_309_5, wires_1237_6,addr_1237_6);

wire[3:0] wires_1238_6;

wire[31:0] addr_1238_6;

Selector_2 s1238_6(wires_309_5[2], addr_309_5, wires_1238_6,addr_1238_6);

wire[3:0] wires_1239_6;

wire[31:0] addr_1239_6;

Selector_2 s1239_6(wires_309_5[3], addr_309_5, wires_1239_6,addr_1239_6);

wire[3:0] wires_1240_6;

wire[31:0] addr_1240_6;

Selector_2 s1240_6(wires_310_5[0], addr_310_5, wires_1240_6,addr_1240_6);

wire[3:0] wires_1241_6;

wire[31:0] addr_1241_6;

Selector_2 s1241_6(wires_310_5[1], addr_310_5, wires_1241_6,addr_1241_6);

wire[3:0] wires_1242_6;

wire[31:0] addr_1242_6;

Selector_2 s1242_6(wires_310_5[2], addr_310_5, wires_1242_6,addr_1242_6);

wire[3:0] wires_1243_6;

wire[31:0] addr_1243_6;

Selector_2 s1243_6(wires_310_5[3], addr_310_5, wires_1243_6,addr_1243_6);

wire[3:0] wires_1244_6;

wire[31:0] addr_1244_6;

Selector_2 s1244_6(wires_311_5[0], addr_311_5, wires_1244_6,addr_1244_6);

wire[3:0] wires_1245_6;

wire[31:0] addr_1245_6;

Selector_2 s1245_6(wires_311_5[1], addr_311_5, wires_1245_6,addr_1245_6);

wire[3:0] wires_1246_6;

wire[31:0] addr_1246_6;

Selector_2 s1246_6(wires_311_5[2], addr_311_5, wires_1246_6,addr_1246_6);

wire[3:0] wires_1247_6;

wire[31:0] addr_1247_6;

Selector_2 s1247_6(wires_311_5[3], addr_311_5, wires_1247_6,addr_1247_6);

wire[3:0] wires_1248_6;

wire[31:0] addr_1248_6;

Selector_2 s1248_6(wires_312_5[0], addr_312_5, wires_1248_6,addr_1248_6);

wire[3:0] wires_1249_6;

wire[31:0] addr_1249_6;

Selector_2 s1249_6(wires_312_5[1], addr_312_5, wires_1249_6,addr_1249_6);

wire[3:0] wires_1250_6;

wire[31:0] addr_1250_6;

Selector_2 s1250_6(wires_312_5[2], addr_312_5, wires_1250_6,addr_1250_6);

wire[3:0] wires_1251_6;

wire[31:0] addr_1251_6;

Selector_2 s1251_6(wires_312_5[3], addr_312_5, wires_1251_6,addr_1251_6);

wire[3:0] wires_1252_6;

wire[31:0] addr_1252_6;

Selector_2 s1252_6(wires_313_5[0], addr_313_5, wires_1252_6,addr_1252_6);

wire[3:0] wires_1253_6;

wire[31:0] addr_1253_6;

Selector_2 s1253_6(wires_313_5[1], addr_313_5, wires_1253_6,addr_1253_6);

wire[3:0] wires_1254_6;

wire[31:0] addr_1254_6;

Selector_2 s1254_6(wires_313_5[2], addr_313_5, wires_1254_6,addr_1254_6);

wire[3:0] wires_1255_6;

wire[31:0] addr_1255_6;

Selector_2 s1255_6(wires_313_5[3], addr_313_5, wires_1255_6,addr_1255_6);

wire[3:0] wires_1256_6;

wire[31:0] addr_1256_6;

Selector_2 s1256_6(wires_314_5[0], addr_314_5, wires_1256_6,addr_1256_6);

wire[3:0] wires_1257_6;

wire[31:0] addr_1257_6;

Selector_2 s1257_6(wires_314_5[1], addr_314_5, wires_1257_6,addr_1257_6);

wire[3:0] wires_1258_6;

wire[31:0] addr_1258_6;

Selector_2 s1258_6(wires_314_5[2], addr_314_5, wires_1258_6,addr_1258_6);

wire[3:0] wires_1259_6;

wire[31:0] addr_1259_6;

Selector_2 s1259_6(wires_314_5[3], addr_314_5, wires_1259_6,addr_1259_6);

wire[3:0] wires_1260_6;

wire[31:0] addr_1260_6;

Selector_2 s1260_6(wires_315_5[0], addr_315_5, wires_1260_6,addr_1260_6);

wire[3:0] wires_1261_6;

wire[31:0] addr_1261_6;

Selector_2 s1261_6(wires_315_5[1], addr_315_5, wires_1261_6,addr_1261_6);

wire[3:0] wires_1262_6;

wire[31:0] addr_1262_6;

Selector_2 s1262_6(wires_315_5[2], addr_315_5, wires_1262_6,addr_1262_6);

wire[3:0] wires_1263_6;

wire[31:0] addr_1263_6;

Selector_2 s1263_6(wires_315_5[3], addr_315_5, wires_1263_6,addr_1263_6);

wire[3:0] wires_1264_6;

wire[31:0] addr_1264_6;

Selector_2 s1264_6(wires_316_5[0], addr_316_5, wires_1264_6,addr_1264_6);

wire[3:0] wires_1265_6;

wire[31:0] addr_1265_6;

Selector_2 s1265_6(wires_316_5[1], addr_316_5, wires_1265_6,addr_1265_6);

wire[3:0] wires_1266_6;

wire[31:0] addr_1266_6;

Selector_2 s1266_6(wires_316_5[2], addr_316_5, wires_1266_6,addr_1266_6);

wire[3:0] wires_1267_6;

wire[31:0] addr_1267_6;

Selector_2 s1267_6(wires_316_5[3], addr_316_5, wires_1267_6,addr_1267_6);

wire[3:0] wires_1268_6;

wire[31:0] addr_1268_6;

Selector_2 s1268_6(wires_317_5[0], addr_317_5, wires_1268_6,addr_1268_6);

wire[3:0] wires_1269_6;

wire[31:0] addr_1269_6;

Selector_2 s1269_6(wires_317_5[1], addr_317_5, wires_1269_6,addr_1269_6);

wire[3:0] wires_1270_6;

wire[31:0] addr_1270_6;

Selector_2 s1270_6(wires_317_5[2], addr_317_5, wires_1270_6,addr_1270_6);

wire[3:0] wires_1271_6;

wire[31:0] addr_1271_6;

Selector_2 s1271_6(wires_317_5[3], addr_317_5, wires_1271_6,addr_1271_6);

wire[3:0] wires_1272_6;

wire[31:0] addr_1272_6;

Selector_2 s1272_6(wires_318_5[0], addr_318_5, wires_1272_6,addr_1272_6);

wire[3:0] wires_1273_6;

wire[31:0] addr_1273_6;

Selector_2 s1273_6(wires_318_5[1], addr_318_5, wires_1273_6,addr_1273_6);

wire[3:0] wires_1274_6;

wire[31:0] addr_1274_6;

Selector_2 s1274_6(wires_318_5[2], addr_318_5, wires_1274_6,addr_1274_6);

wire[3:0] wires_1275_6;

wire[31:0] addr_1275_6;

Selector_2 s1275_6(wires_318_5[3], addr_318_5, wires_1275_6,addr_1275_6);

wire[3:0] wires_1276_6;

wire[31:0] addr_1276_6;

Selector_2 s1276_6(wires_319_5[0], addr_319_5, wires_1276_6,addr_1276_6);

wire[3:0] wires_1277_6;

wire[31:0] addr_1277_6;

Selector_2 s1277_6(wires_319_5[1], addr_319_5, wires_1277_6,addr_1277_6);

wire[3:0] wires_1278_6;

wire[31:0] addr_1278_6;

Selector_2 s1278_6(wires_319_5[2], addr_319_5, wires_1278_6,addr_1278_6);

wire[3:0] wires_1279_6;

wire[31:0] addr_1279_6;

Selector_2 s1279_6(wires_319_5[3], addr_319_5, wires_1279_6,addr_1279_6);

wire[3:0] wires_1280_6;

wire[31:0] addr_1280_6;

Selector_2 s1280_6(wires_320_5[0], addr_320_5, wires_1280_6,addr_1280_6);

wire[3:0] wires_1281_6;

wire[31:0] addr_1281_6;

Selector_2 s1281_6(wires_320_5[1], addr_320_5, wires_1281_6,addr_1281_6);

wire[3:0] wires_1282_6;

wire[31:0] addr_1282_6;

Selector_2 s1282_6(wires_320_5[2], addr_320_5, wires_1282_6,addr_1282_6);

wire[3:0] wires_1283_6;

wire[31:0] addr_1283_6;

Selector_2 s1283_6(wires_320_5[3], addr_320_5, wires_1283_6,addr_1283_6);

wire[3:0] wires_1284_6;

wire[31:0] addr_1284_6;

Selector_2 s1284_6(wires_321_5[0], addr_321_5, wires_1284_6,addr_1284_6);

wire[3:0] wires_1285_6;

wire[31:0] addr_1285_6;

Selector_2 s1285_6(wires_321_5[1], addr_321_5, wires_1285_6,addr_1285_6);

wire[3:0] wires_1286_6;

wire[31:0] addr_1286_6;

Selector_2 s1286_6(wires_321_5[2], addr_321_5, wires_1286_6,addr_1286_6);

wire[3:0] wires_1287_6;

wire[31:0] addr_1287_6;

Selector_2 s1287_6(wires_321_5[3], addr_321_5, wires_1287_6,addr_1287_6);

wire[3:0] wires_1288_6;

wire[31:0] addr_1288_6;

Selector_2 s1288_6(wires_322_5[0], addr_322_5, wires_1288_6,addr_1288_6);

wire[3:0] wires_1289_6;

wire[31:0] addr_1289_6;

Selector_2 s1289_6(wires_322_5[1], addr_322_5, wires_1289_6,addr_1289_6);

wire[3:0] wires_1290_6;

wire[31:0] addr_1290_6;

Selector_2 s1290_6(wires_322_5[2], addr_322_5, wires_1290_6,addr_1290_6);

wire[3:0] wires_1291_6;

wire[31:0] addr_1291_6;

Selector_2 s1291_6(wires_322_5[3], addr_322_5, wires_1291_6,addr_1291_6);

wire[3:0] wires_1292_6;

wire[31:0] addr_1292_6;

Selector_2 s1292_6(wires_323_5[0], addr_323_5, wires_1292_6,addr_1292_6);

wire[3:0] wires_1293_6;

wire[31:0] addr_1293_6;

Selector_2 s1293_6(wires_323_5[1], addr_323_5, wires_1293_6,addr_1293_6);

wire[3:0] wires_1294_6;

wire[31:0] addr_1294_6;

Selector_2 s1294_6(wires_323_5[2], addr_323_5, wires_1294_6,addr_1294_6);

wire[3:0] wires_1295_6;

wire[31:0] addr_1295_6;

Selector_2 s1295_6(wires_323_5[3], addr_323_5, wires_1295_6,addr_1295_6);

wire[3:0] wires_1296_6;

wire[31:0] addr_1296_6;

Selector_2 s1296_6(wires_324_5[0], addr_324_5, wires_1296_6,addr_1296_6);

wire[3:0] wires_1297_6;

wire[31:0] addr_1297_6;

Selector_2 s1297_6(wires_324_5[1], addr_324_5, wires_1297_6,addr_1297_6);

wire[3:0] wires_1298_6;

wire[31:0] addr_1298_6;

Selector_2 s1298_6(wires_324_5[2], addr_324_5, wires_1298_6,addr_1298_6);

wire[3:0] wires_1299_6;

wire[31:0] addr_1299_6;

Selector_2 s1299_6(wires_324_5[3], addr_324_5, wires_1299_6,addr_1299_6);

wire[3:0] wires_1300_6;

wire[31:0] addr_1300_6;

Selector_2 s1300_6(wires_325_5[0], addr_325_5, wires_1300_6,addr_1300_6);

wire[3:0] wires_1301_6;

wire[31:0] addr_1301_6;

Selector_2 s1301_6(wires_325_5[1], addr_325_5, wires_1301_6,addr_1301_6);

wire[3:0] wires_1302_6;

wire[31:0] addr_1302_6;

Selector_2 s1302_6(wires_325_5[2], addr_325_5, wires_1302_6,addr_1302_6);

wire[3:0] wires_1303_6;

wire[31:0] addr_1303_6;

Selector_2 s1303_6(wires_325_5[3], addr_325_5, wires_1303_6,addr_1303_6);

wire[3:0] wires_1304_6;

wire[31:0] addr_1304_6;

Selector_2 s1304_6(wires_326_5[0], addr_326_5, wires_1304_6,addr_1304_6);

wire[3:0] wires_1305_6;

wire[31:0] addr_1305_6;

Selector_2 s1305_6(wires_326_5[1], addr_326_5, wires_1305_6,addr_1305_6);

wire[3:0] wires_1306_6;

wire[31:0] addr_1306_6;

Selector_2 s1306_6(wires_326_5[2], addr_326_5, wires_1306_6,addr_1306_6);

wire[3:0] wires_1307_6;

wire[31:0] addr_1307_6;

Selector_2 s1307_6(wires_326_5[3], addr_326_5, wires_1307_6,addr_1307_6);

wire[3:0] wires_1308_6;

wire[31:0] addr_1308_6;

Selector_2 s1308_6(wires_327_5[0], addr_327_5, wires_1308_6,addr_1308_6);

wire[3:0] wires_1309_6;

wire[31:0] addr_1309_6;

Selector_2 s1309_6(wires_327_5[1], addr_327_5, wires_1309_6,addr_1309_6);

wire[3:0] wires_1310_6;

wire[31:0] addr_1310_6;

Selector_2 s1310_6(wires_327_5[2], addr_327_5, wires_1310_6,addr_1310_6);

wire[3:0] wires_1311_6;

wire[31:0] addr_1311_6;

Selector_2 s1311_6(wires_327_5[3], addr_327_5, wires_1311_6,addr_1311_6);

wire[3:0] wires_1312_6;

wire[31:0] addr_1312_6;

Selector_2 s1312_6(wires_328_5[0], addr_328_5, wires_1312_6,addr_1312_6);

wire[3:0] wires_1313_6;

wire[31:0] addr_1313_6;

Selector_2 s1313_6(wires_328_5[1], addr_328_5, wires_1313_6,addr_1313_6);

wire[3:0] wires_1314_6;

wire[31:0] addr_1314_6;

Selector_2 s1314_6(wires_328_5[2], addr_328_5, wires_1314_6,addr_1314_6);

wire[3:0] wires_1315_6;

wire[31:0] addr_1315_6;

Selector_2 s1315_6(wires_328_5[3], addr_328_5, wires_1315_6,addr_1315_6);

wire[3:0] wires_1316_6;

wire[31:0] addr_1316_6;

Selector_2 s1316_6(wires_329_5[0], addr_329_5, wires_1316_6,addr_1316_6);

wire[3:0] wires_1317_6;

wire[31:0] addr_1317_6;

Selector_2 s1317_6(wires_329_5[1], addr_329_5, wires_1317_6,addr_1317_6);

wire[3:0] wires_1318_6;

wire[31:0] addr_1318_6;

Selector_2 s1318_6(wires_329_5[2], addr_329_5, wires_1318_6,addr_1318_6);

wire[3:0] wires_1319_6;

wire[31:0] addr_1319_6;

Selector_2 s1319_6(wires_329_5[3], addr_329_5, wires_1319_6,addr_1319_6);

wire[3:0] wires_1320_6;

wire[31:0] addr_1320_6;

Selector_2 s1320_6(wires_330_5[0], addr_330_5, wires_1320_6,addr_1320_6);

wire[3:0] wires_1321_6;

wire[31:0] addr_1321_6;

Selector_2 s1321_6(wires_330_5[1], addr_330_5, wires_1321_6,addr_1321_6);

wire[3:0] wires_1322_6;

wire[31:0] addr_1322_6;

Selector_2 s1322_6(wires_330_5[2], addr_330_5, wires_1322_6,addr_1322_6);

wire[3:0] wires_1323_6;

wire[31:0] addr_1323_6;

Selector_2 s1323_6(wires_330_5[3], addr_330_5, wires_1323_6,addr_1323_6);

wire[3:0] wires_1324_6;

wire[31:0] addr_1324_6;

Selector_2 s1324_6(wires_331_5[0], addr_331_5, wires_1324_6,addr_1324_6);

wire[3:0] wires_1325_6;

wire[31:0] addr_1325_6;

Selector_2 s1325_6(wires_331_5[1], addr_331_5, wires_1325_6,addr_1325_6);

wire[3:0] wires_1326_6;

wire[31:0] addr_1326_6;

Selector_2 s1326_6(wires_331_5[2], addr_331_5, wires_1326_6,addr_1326_6);

wire[3:0] wires_1327_6;

wire[31:0] addr_1327_6;

Selector_2 s1327_6(wires_331_5[3], addr_331_5, wires_1327_6,addr_1327_6);

wire[3:0] wires_1328_6;

wire[31:0] addr_1328_6;

Selector_2 s1328_6(wires_332_5[0], addr_332_5, wires_1328_6,addr_1328_6);

wire[3:0] wires_1329_6;

wire[31:0] addr_1329_6;

Selector_2 s1329_6(wires_332_5[1], addr_332_5, wires_1329_6,addr_1329_6);

wire[3:0] wires_1330_6;

wire[31:0] addr_1330_6;

Selector_2 s1330_6(wires_332_5[2], addr_332_5, wires_1330_6,addr_1330_6);

wire[3:0] wires_1331_6;

wire[31:0] addr_1331_6;

Selector_2 s1331_6(wires_332_5[3], addr_332_5, wires_1331_6,addr_1331_6);

wire[3:0] wires_1332_6;

wire[31:0] addr_1332_6;

Selector_2 s1332_6(wires_333_5[0], addr_333_5, wires_1332_6,addr_1332_6);

wire[3:0] wires_1333_6;

wire[31:0] addr_1333_6;

Selector_2 s1333_6(wires_333_5[1], addr_333_5, wires_1333_6,addr_1333_6);

wire[3:0] wires_1334_6;

wire[31:0] addr_1334_6;

Selector_2 s1334_6(wires_333_5[2], addr_333_5, wires_1334_6,addr_1334_6);

wire[3:0] wires_1335_6;

wire[31:0] addr_1335_6;

Selector_2 s1335_6(wires_333_5[3], addr_333_5, wires_1335_6,addr_1335_6);

wire[3:0] wires_1336_6;

wire[31:0] addr_1336_6;

Selector_2 s1336_6(wires_334_5[0], addr_334_5, wires_1336_6,addr_1336_6);

wire[3:0] wires_1337_6;

wire[31:0] addr_1337_6;

Selector_2 s1337_6(wires_334_5[1], addr_334_5, wires_1337_6,addr_1337_6);

wire[3:0] wires_1338_6;

wire[31:0] addr_1338_6;

Selector_2 s1338_6(wires_334_5[2], addr_334_5, wires_1338_6,addr_1338_6);

wire[3:0] wires_1339_6;

wire[31:0] addr_1339_6;

Selector_2 s1339_6(wires_334_5[3], addr_334_5, wires_1339_6,addr_1339_6);

wire[3:0] wires_1340_6;

wire[31:0] addr_1340_6;

Selector_2 s1340_6(wires_335_5[0], addr_335_5, wires_1340_6,addr_1340_6);

wire[3:0] wires_1341_6;

wire[31:0] addr_1341_6;

Selector_2 s1341_6(wires_335_5[1], addr_335_5, wires_1341_6,addr_1341_6);

wire[3:0] wires_1342_6;

wire[31:0] addr_1342_6;

Selector_2 s1342_6(wires_335_5[2], addr_335_5, wires_1342_6,addr_1342_6);

wire[3:0] wires_1343_6;

wire[31:0] addr_1343_6;

Selector_2 s1343_6(wires_335_5[3], addr_335_5, wires_1343_6,addr_1343_6);

wire[3:0] wires_1344_6;

wire[31:0] addr_1344_6;

Selector_2 s1344_6(wires_336_5[0], addr_336_5, wires_1344_6,addr_1344_6);

wire[3:0] wires_1345_6;

wire[31:0] addr_1345_6;

Selector_2 s1345_6(wires_336_5[1], addr_336_5, wires_1345_6,addr_1345_6);

wire[3:0] wires_1346_6;

wire[31:0] addr_1346_6;

Selector_2 s1346_6(wires_336_5[2], addr_336_5, wires_1346_6,addr_1346_6);

wire[3:0] wires_1347_6;

wire[31:0] addr_1347_6;

Selector_2 s1347_6(wires_336_5[3], addr_336_5, wires_1347_6,addr_1347_6);

wire[3:0] wires_1348_6;

wire[31:0] addr_1348_6;

Selector_2 s1348_6(wires_337_5[0], addr_337_5, wires_1348_6,addr_1348_6);

wire[3:0] wires_1349_6;

wire[31:0] addr_1349_6;

Selector_2 s1349_6(wires_337_5[1], addr_337_5, wires_1349_6,addr_1349_6);

wire[3:0] wires_1350_6;

wire[31:0] addr_1350_6;

Selector_2 s1350_6(wires_337_5[2], addr_337_5, wires_1350_6,addr_1350_6);

wire[3:0] wires_1351_6;

wire[31:0] addr_1351_6;

Selector_2 s1351_6(wires_337_5[3], addr_337_5, wires_1351_6,addr_1351_6);

wire[3:0] wires_1352_6;

wire[31:0] addr_1352_6;

Selector_2 s1352_6(wires_338_5[0], addr_338_5, wires_1352_6,addr_1352_6);

wire[3:0] wires_1353_6;

wire[31:0] addr_1353_6;

Selector_2 s1353_6(wires_338_5[1], addr_338_5, wires_1353_6,addr_1353_6);

wire[3:0] wires_1354_6;

wire[31:0] addr_1354_6;

Selector_2 s1354_6(wires_338_5[2], addr_338_5, wires_1354_6,addr_1354_6);

wire[3:0] wires_1355_6;

wire[31:0] addr_1355_6;

Selector_2 s1355_6(wires_338_5[3], addr_338_5, wires_1355_6,addr_1355_6);

wire[3:0] wires_1356_6;

wire[31:0] addr_1356_6;

Selector_2 s1356_6(wires_339_5[0], addr_339_5, wires_1356_6,addr_1356_6);

wire[3:0] wires_1357_6;

wire[31:0] addr_1357_6;

Selector_2 s1357_6(wires_339_5[1], addr_339_5, wires_1357_6,addr_1357_6);

wire[3:0] wires_1358_6;

wire[31:0] addr_1358_6;

Selector_2 s1358_6(wires_339_5[2], addr_339_5, wires_1358_6,addr_1358_6);

wire[3:0] wires_1359_6;

wire[31:0] addr_1359_6;

Selector_2 s1359_6(wires_339_5[3], addr_339_5, wires_1359_6,addr_1359_6);

wire[3:0] wires_1360_6;

wire[31:0] addr_1360_6;

Selector_2 s1360_6(wires_340_5[0], addr_340_5, wires_1360_6,addr_1360_6);

wire[3:0] wires_1361_6;

wire[31:0] addr_1361_6;

Selector_2 s1361_6(wires_340_5[1], addr_340_5, wires_1361_6,addr_1361_6);

wire[3:0] wires_1362_6;

wire[31:0] addr_1362_6;

Selector_2 s1362_6(wires_340_5[2], addr_340_5, wires_1362_6,addr_1362_6);

wire[3:0] wires_1363_6;

wire[31:0] addr_1363_6;

Selector_2 s1363_6(wires_340_5[3], addr_340_5, wires_1363_6,addr_1363_6);

wire[3:0] wires_1364_6;

wire[31:0] addr_1364_6;

Selector_2 s1364_6(wires_341_5[0], addr_341_5, wires_1364_6,addr_1364_6);

wire[3:0] wires_1365_6;

wire[31:0] addr_1365_6;

Selector_2 s1365_6(wires_341_5[1], addr_341_5, wires_1365_6,addr_1365_6);

wire[3:0] wires_1366_6;

wire[31:0] addr_1366_6;

Selector_2 s1366_6(wires_341_5[2], addr_341_5, wires_1366_6,addr_1366_6);

wire[3:0] wires_1367_6;

wire[31:0] addr_1367_6;

Selector_2 s1367_6(wires_341_5[3], addr_341_5, wires_1367_6,addr_1367_6);

wire[3:0] wires_1368_6;

wire[31:0] addr_1368_6;

Selector_2 s1368_6(wires_342_5[0], addr_342_5, wires_1368_6,addr_1368_6);

wire[3:0] wires_1369_6;

wire[31:0] addr_1369_6;

Selector_2 s1369_6(wires_342_5[1], addr_342_5, wires_1369_6,addr_1369_6);

wire[3:0] wires_1370_6;

wire[31:0] addr_1370_6;

Selector_2 s1370_6(wires_342_5[2], addr_342_5, wires_1370_6,addr_1370_6);

wire[3:0] wires_1371_6;

wire[31:0] addr_1371_6;

Selector_2 s1371_6(wires_342_5[3], addr_342_5, wires_1371_6,addr_1371_6);

wire[3:0] wires_1372_6;

wire[31:0] addr_1372_6;

Selector_2 s1372_6(wires_343_5[0], addr_343_5, wires_1372_6,addr_1372_6);

wire[3:0] wires_1373_6;

wire[31:0] addr_1373_6;

Selector_2 s1373_6(wires_343_5[1], addr_343_5, wires_1373_6,addr_1373_6);

wire[3:0] wires_1374_6;

wire[31:0] addr_1374_6;

Selector_2 s1374_6(wires_343_5[2], addr_343_5, wires_1374_6,addr_1374_6);

wire[3:0] wires_1375_6;

wire[31:0] addr_1375_6;

Selector_2 s1375_6(wires_343_5[3], addr_343_5, wires_1375_6,addr_1375_6);

wire[3:0] wires_1376_6;

wire[31:0] addr_1376_6;

Selector_2 s1376_6(wires_344_5[0], addr_344_5, wires_1376_6,addr_1376_6);

wire[3:0] wires_1377_6;

wire[31:0] addr_1377_6;

Selector_2 s1377_6(wires_344_5[1], addr_344_5, wires_1377_6,addr_1377_6);

wire[3:0] wires_1378_6;

wire[31:0] addr_1378_6;

Selector_2 s1378_6(wires_344_5[2], addr_344_5, wires_1378_6,addr_1378_6);

wire[3:0] wires_1379_6;

wire[31:0] addr_1379_6;

Selector_2 s1379_6(wires_344_5[3], addr_344_5, wires_1379_6,addr_1379_6);

wire[3:0] wires_1380_6;

wire[31:0] addr_1380_6;

Selector_2 s1380_6(wires_345_5[0], addr_345_5, wires_1380_6,addr_1380_6);

wire[3:0] wires_1381_6;

wire[31:0] addr_1381_6;

Selector_2 s1381_6(wires_345_5[1], addr_345_5, wires_1381_6,addr_1381_6);

wire[3:0] wires_1382_6;

wire[31:0] addr_1382_6;

Selector_2 s1382_6(wires_345_5[2], addr_345_5, wires_1382_6,addr_1382_6);

wire[3:0] wires_1383_6;

wire[31:0] addr_1383_6;

Selector_2 s1383_6(wires_345_5[3], addr_345_5, wires_1383_6,addr_1383_6);

wire[3:0] wires_1384_6;

wire[31:0] addr_1384_6;

Selector_2 s1384_6(wires_346_5[0], addr_346_5, wires_1384_6,addr_1384_6);

wire[3:0] wires_1385_6;

wire[31:0] addr_1385_6;

Selector_2 s1385_6(wires_346_5[1], addr_346_5, wires_1385_6,addr_1385_6);

wire[3:0] wires_1386_6;

wire[31:0] addr_1386_6;

Selector_2 s1386_6(wires_346_5[2], addr_346_5, wires_1386_6,addr_1386_6);

wire[3:0] wires_1387_6;

wire[31:0] addr_1387_6;

Selector_2 s1387_6(wires_346_5[3], addr_346_5, wires_1387_6,addr_1387_6);

wire[3:0] wires_1388_6;

wire[31:0] addr_1388_6;

Selector_2 s1388_6(wires_347_5[0], addr_347_5, wires_1388_6,addr_1388_6);

wire[3:0] wires_1389_6;

wire[31:0] addr_1389_6;

Selector_2 s1389_6(wires_347_5[1], addr_347_5, wires_1389_6,addr_1389_6);

wire[3:0] wires_1390_6;

wire[31:0] addr_1390_6;

Selector_2 s1390_6(wires_347_5[2], addr_347_5, wires_1390_6,addr_1390_6);

wire[3:0] wires_1391_6;

wire[31:0] addr_1391_6;

Selector_2 s1391_6(wires_347_5[3], addr_347_5, wires_1391_6,addr_1391_6);

wire[3:0] wires_1392_6;

wire[31:0] addr_1392_6;

Selector_2 s1392_6(wires_348_5[0], addr_348_5, wires_1392_6,addr_1392_6);

wire[3:0] wires_1393_6;

wire[31:0] addr_1393_6;

Selector_2 s1393_6(wires_348_5[1], addr_348_5, wires_1393_6,addr_1393_6);

wire[3:0] wires_1394_6;

wire[31:0] addr_1394_6;

Selector_2 s1394_6(wires_348_5[2], addr_348_5, wires_1394_6,addr_1394_6);

wire[3:0] wires_1395_6;

wire[31:0] addr_1395_6;

Selector_2 s1395_6(wires_348_5[3], addr_348_5, wires_1395_6,addr_1395_6);

wire[3:0] wires_1396_6;

wire[31:0] addr_1396_6;

Selector_2 s1396_6(wires_349_5[0], addr_349_5, wires_1396_6,addr_1396_6);

wire[3:0] wires_1397_6;

wire[31:0] addr_1397_6;

Selector_2 s1397_6(wires_349_5[1], addr_349_5, wires_1397_6,addr_1397_6);

wire[3:0] wires_1398_6;

wire[31:0] addr_1398_6;

Selector_2 s1398_6(wires_349_5[2], addr_349_5, wires_1398_6,addr_1398_6);

wire[3:0] wires_1399_6;

wire[31:0] addr_1399_6;

Selector_2 s1399_6(wires_349_5[3], addr_349_5, wires_1399_6,addr_1399_6);

wire[3:0] wires_1400_6;

wire[31:0] addr_1400_6;

Selector_2 s1400_6(wires_350_5[0], addr_350_5, wires_1400_6,addr_1400_6);

wire[3:0] wires_1401_6;

wire[31:0] addr_1401_6;

Selector_2 s1401_6(wires_350_5[1], addr_350_5, wires_1401_6,addr_1401_6);

wire[3:0] wires_1402_6;

wire[31:0] addr_1402_6;

Selector_2 s1402_6(wires_350_5[2], addr_350_5, wires_1402_6,addr_1402_6);

wire[3:0] wires_1403_6;

wire[31:0] addr_1403_6;

Selector_2 s1403_6(wires_350_5[3], addr_350_5, wires_1403_6,addr_1403_6);

wire[3:0] wires_1404_6;

wire[31:0] addr_1404_6;

Selector_2 s1404_6(wires_351_5[0], addr_351_5, wires_1404_6,addr_1404_6);

wire[3:0] wires_1405_6;

wire[31:0] addr_1405_6;

Selector_2 s1405_6(wires_351_5[1], addr_351_5, wires_1405_6,addr_1405_6);

wire[3:0] wires_1406_6;

wire[31:0] addr_1406_6;

Selector_2 s1406_6(wires_351_5[2], addr_351_5, wires_1406_6,addr_1406_6);

wire[3:0] wires_1407_6;

wire[31:0] addr_1407_6;

Selector_2 s1407_6(wires_351_5[3], addr_351_5, wires_1407_6,addr_1407_6);

wire[3:0] wires_1408_6;

wire[31:0] addr_1408_6;

Selector_2 s1408_6(wires_352_5[0], addr_352_5, wires_1408_6,addr_1408_6);

wire[3:0] wires_1409_6;

wire[31:0] addr_1409_6;

Selector_2 s1409_6(wires_352_5[1], addr_352_5, wires_1409_6,addr_1409_6);

wire[3:0] wires_1410_6;

wire[31:0] addr_1410_6;

Selector_2 s1410_6(wires_352_5[2], addr_352_5, wires_1410_6,addr_1410_6);

wire[3:0] wires_1411_6;

wire[31:0] addr_1411_6;

Selector_2 s1411_6(wires_352_5[3], addr_352_5, wires_1411_6,addr_1411_6);

wire[3:0] wires_1412_6;

wire[31:0] addr_1412_6;

Selector_2 s1412_6(wires_353_5[0], addr_353_5, wires_1412_6,addr_1412_6);

wire[3:0] wires_1413_6;

wire[31:0] addr_1413_6;

Selector_2 s1413_6(wires_353_5[1], addr_353_5, wires_1413_6,addr_1413_6);

wire[3:0] wires_1414_6;

wire[31:0] addr_1414_6;

Selector_2 s1414_6(wires_353_5[2], addr_353_5, wires_1414_6,addr_1414_6);

wire[3:0] wires_1415_6;

wire[31:0] addr_1415_6;

Selector_2 s1415_6(wires_353_5[3], addr_353_5, wires_1415_6,addr_1415_6);

wire[3:0] wires_1416_6;

wire[31:0] addr_1416_6;

Selector_2 s1416_6(wires_354_5[0], addr_354_5, wires_1416_6,addr_1416_6);

wire[3:0] wires_1417_6;

wire[31:0] addr_1417_6;

Selector_2 s1417_6(wires_354_5[1], addr_354_5, wires_1417_6,addr_1417_6);

wire[3:0] wires_1418_6;

wire[31:0] addr_1418_6;

Selector_2 s1418_6(wires_354_5[2], addr_354_5, wires_1418_6,addr_1418_6);

wire[3:0] wires_1419_6;

wire[31:0] addr_1419_6;

Selector_2 s1419_6(wires_354_5[3], addr_354_5, wires_1419_6,addr_1419_6);

wire[3:0] wires_1420_6;

wire[31:0] addr_1420_6;

Selector_2 s1420_6(wires_355_5[0], addr_355_5, wires_1420_6,addr_1420_6);

wire[3:0] wires_1421_6;

wire[31:0] addr_1421_6;

Selector_2 s1421_6(wires_355_5[1], addr_355_5, wires_1421_6,addr_1421_6);

wire[3:0] wires_1422_6;

wire[31:0] addr_1422_6;

Selector_2 s1422_6(wires_355_5[2], addr_355_5, wires_1422_6,addr_1422_6);

wire[3:0] wires_1423_6;

wire[31:0] addr_1423_6;

Selector_2 s1423_6(wires_355_5[3], addr_355_5, wires_1423_6,addr_1423_6);

wire[3:0] wires_1424_6;

wire[31:0] addr_1424_6;

Selector_2 s1424_6(wires_356_5[0], addr_356_5, wires_1424_6,addr_1424_6);

wire[3:0] wires_1425_6;

wire[31:0] addr_1425_6;

Selector_2 s1425_6(wires_356_5[1], addr_356_5, wires_1425_6,addr_1425_6);

wire[3:0] wires_1426_6;

wire[31:0] addr_1426_6;

Selector_2 s1426_6(wires_356_5[2], addr_356_5, wires_1426_6,addr_1426_6);

wire[3:0] wires_1427_6;

wire[31:0] addr_1427_6;

Selector_2 s1427_6(wires_356_5[3], addr_356_5, wires_1427_6,addr_1427_6);

wire[3:0] wires_1428_6;

wire[31:0] addr_1428_6;

Selector_2 s1428_6(wires_357_5[0], addr_357_5, wires_1428_6,addr_1428_6);

wire[3:0] wires_1429_6;

wire[31:0] addr_1429_6;

Selector_2 s1429_6(wires_357_5[1], addr_357_5, wires_1429_6,addr_1429_6);

wire[3:0] wires_1430_6;

wire[31:0] addr_1430_6;

Selector_2 s1430_6(wires_357_5[2], addr_357_5, wires_1430_6,addr_1430_6);

wire[3:0] wires_1431_6;

wire[31:0] addr_1431_6;

Selector_2 s1431_6(wires_357_5[3], addr_357_5, wires_1431_6,addr_1431_6);

wire[3:0] wires_1432_6;

wire[31:0] addr_1432_6;

Selector_2 s1432_6(wires_358_5[0], addr_358_5, wires_1432_6,addr_1432_6);

wire[3:0] wires_1433_6;

wire[31:0] addr_1433_6;

Selector_2 s1433_6(wires_358_5[1], addr_358_5, wires_1433_6,addr_1433_6);

wire[3:0] wires_1434_6;

wire[31:0] addr_1434_6;

Selector_2 s1434_6(wires_358_5[2], addr_358_5, wires_1434_6,addr_1434_6);

wire[3:0] wires_1435_6;

wire[31:0] addr_1435_6;

Selector_2 s1435_6(wires_358_5[3], addr_358_5, wires_1435_6,addr_1435_6);

wire[3:0] wires_1436_6;

wire[31:0] addr_1436_6;

Selector_2 s1436_6(wires_359_5[0], addr_359_5, wires_1436_6,addr_1436_6);

wire[3:0] wires_1437_6;

wire[31:0] addr_1437_6;

Selector_2 s1437_6(wires_359_5[1], addr_359_5, wires_1437_6,addr_1437_6);

wire[3:0] wires_1438_6;

wire[31:0] addr_1438_6;

Selector_2 s1438_6(wires_359_5[2], addr_359_5, wires_1438_6,addr_1438_6);

wire[3:0] wires_1439_6;

wire[31:0] addr_1439_6;

Selector_2 s1439_6(wires_359_5[3], addr_359_5, wires_1439_6,addr_1439_6);

wire[3:0] wires_1440_6;

wire[31:0] addr_1440_6;

Selector_2 s1440_6(wires_360_5[0], addr_360_5, wires_1440_6,addr_1440_6);

wire[3:0] wires_1441_6;

wire[31:0] addr_1441_6;

Selector_2 s1441_6(wires_360_5[1], addr_360_5, wires_1441_6,addr_1441_6);

wire[3:0] wires_1442_6;

wire[31:0] addr_1442_6;

Selector_2 s1442_6(wires_360_5[2], addr_360_5, wires_1442_6,addr_1442_6);

wire[3:0] wires_1443_6;

wire[31:0] addr_1443_6;

Selector_2 s1443_6(wires_360_5[3], addr_360_5, wires_1443_6,addr_1443_6);

wire[3:0] wires_1444_6;

wire[31:0] addr_1444_6;

Selector_2 s1444_6(wires_361_5[0], addr_361_5, wires_1444_6,addr_1444_6);

wire[3:0] wires_1445_6;

wire[31:0] addr_1445_6;

Selector_2 s1445_6(wires_361_5[1], addr_361_5, wires_1445_6,addr_1445_6);

wire[3:0] wires_1446_6;

wire[31:0] addr_1446_6;

Selector_2 s1446_6(wires_361_5[2], addr_361_5, wires_1446_6,addr_1446_6);

wire[3:0] wires_1447_6;

wire[31:0] addr_1447_6;

Selector_2 s1447_6(wires_361_5[3], addr_361_5, wires_1447_6,addr_1447_6);

wire[3:0] wires_1448_6;

wire[31:0] addr_1448_6;

Selector_2 s1448_6(wires_362_5[0], addr_362_5, wires_1448_6,addr_1448_6);

wire[3:0] wires_1449_6;

wire[31:0] addr_1449_6;

Selector_2 s1449_6(wires_362_5[1], addr_362_5, wires_1449_6,addr_1449_6);

wire[3:0] wires_1450_6;

wire[31:0] addr_1450_6;

Selector_2 s1450_6(wires_362_5[2], addr_362_5, wires_1450_6,addr_1450_6);

wire[3:0] wires_1451_6;

wire[31:0] addr_1451_6;

Selector_2 s1451_6(wires_362_5[3], addr_362_5, wires_1451_6,addr_1451_6);

wire[3:0] wires_1452_6;

wire[31:0] addr_1452_6;

Selector_2 s1452_6(wires_363_5[0], addr_363_5, wires_1452_6,addr_1452_6);

wire[3:0] wires_1453_6;

wire[31:0] addr_1453_6;

Selector_2 s1453_6(wires_363_5[1], addr_363_5, wires_1453_6,addr_1453_6);

wire[3:0] wires_1454_6;

wire[31:0] addr_1454_6;

Selector_2 s1454_6(wires_363_5[2], addr_363_5, wires_1454_6,addr_1454_6);

wire[3:0] wires_1455_6;

wire[31:0] addr_1455_6;

Selector_2 s1455_6(wires_363_5[3], addr_363_5, wires_1455_6,addr_1455_6);

wire[3:0] wires_1456_6;

wire[31:0] addr_1456_6;

Selector_2 s1456_6(wires_364_5[0], addr_364_5, wires_1456_6,addr_1456_6);

wire[3:0] wires_1457_6;

wire[31:0] addr_1457_6;

Selector_2 s1457_6(wires_364_5[1], addr_364_5, wires_1457_6,addr_1457_6);

wire[3:0] wires_1458_6;

wire[31:0] addr_1458_6;

Selector_2 s1458_6(wires_364_5[2], addr_364_5, wires_1458_6,addr_1458_6);

wire[3:0] wires_1459_6;

wire[31:0] addr_1459_6;

Selector_2 s1459_6(wires_364_5[3], addr_364_5, wires_1459_6,addr_1459_6);

wire[3:0] wires_1460_6;

wire[31:0] addr_1460_6;

Selector_2 s1460_6(wires_365_5[0], addr_365_5, wires_1460_6,addr_1460_6);

wire[3:0] wires_1461_6;

wire[31:0] addr_1461_6;

Selector_2 s1461_6(wires_365_5[1], addr_365_5, wires_1461_6,addr_1461_6);

wire[3:0] wires_1462_6;

wire[31:0] addr_1462_6;

Selector_2 s1462_6(wires_365_5[2], addr_365_5, wires_1462_6,addr_1462_6);

wire[3:0] wires_1463_6;

wire[31:0] addr_1463_6;

Selector_2 s1463_6(wires_365_5[3], addr_365_5, wires_1463_6,addr_1463_6);

wire[3:0] wires_1464_6;

wire[31:0] addr_1464_6;

Selector_2 s1464_6(wires_366_5[0], addr_366_5, wires_1464_6,addr_1464_6);

wire[3:0] wires_1465_6;

wire[31:0] addr_1465_6;

Selector_2 s1465_6(wires_366_5[1], addr_366_5, wires_1465_6,addr_1465_6);

wire[3:0] wires_1466_6;

wire[31:0] addr_1466_6;

Selector_2 s1466_6(wires_366_5[2], addr_366_5, wires_1466_6,addr_1466_6);

wire[3:0] wires_1467_6;

wire[31:0] addr_1467_6;

Selector_2 s1467_6(wires_366_5[3], addr_366_5, wires_1467_6,addr_1467_6);

wire[3:0] wires_1468_6;

wire[31:0] addr_1468_6;

Selector_2 s1468_6(wires_367_5[0], addr_367_5, wires_1468_6,addr_1468_6);

wire[3:0] wires_1469_6;

wire[31:0] addr_1469_6;

Selector_2 s1469_6(wires_367_5[1], addr_367_5, wires_1469_6,addr_1469_6);

wire[3:0] wires_1470_6;

wire[31:0] addr_1470_6;

Selector_2 s1470_6(wires_367_5[2], addr_367_5, wires_1470_6,addr_1470_6);

wire[3:0] wires_1471_6;

wire[31:0] addr_1471_6;

Selector_2 s1471_6(wires_367_5[3], addr_367_5, wires_1471_6,addr_1471_6);

wire[3:0] wires_1472_6;

wire[31:0] addr_1472_6;

Selector_2 s1472_6(wires_368_5[0], addr_368_5, wires_1472_6,addr_1472_6);

wire[3:0] wires_1473_6;

wire[31:0] addr_1473_6;

Selector_2 s1473_6(wires_368_5[1], addr_368_5, wires_1473_6,addr_1473_6);

wire[3:0] wires_1474_6;

wire[31:0] addr_1474_6;

Selector_2 s1474_6(wires_368_5[2], addr_368_5, wires_1474_6,addr_1474_6);

wire[3:0] wires_1475_6;

wire[31:0] addr_1475_6;

Selector_2 s1475_6(wires_368_5[3], addr_368_5, wires_1475_6,addr_1475_6);

wire[3:0] wires_1476_6;

wire[31:0] addr_1476_6;

Selector_2 s1476_6(wires_369_5[0], addr_369_5, wires_1476_6,addr_1476_6);

wire[3:0] wires_1477_6;

wire[31:0] addr_1477_6;

Selector_2 s1477_6(wires_369_5[1], addr_369_5, wires_1477_6,addr_1477_6);

wire[3:0] wires_1478_6;

wire[31:0] addr_1478_6;

Selector_2 s1478_6(wires_369_5[2], addr_369_5, wires_1478_6,addr_1478_6);

wire[3:0] wires_1479_6;

wire[31:0] addr_1479_6;

Selector_2 s1479_6(wires_369_5[3], addr_369_5, wires_1479_6,addr_1479_6);

wire[3:0] wires_1480_6;

wire[31:0] addr_1480_6;

Selector_2 s1480_6(wires_370_5[0], addr_370_5, wires_1480_6,addr_1480_6);

wire[3:0] wires_1481_6;

wire[31:0] addr_1481_6;

Selector_2 s1481_6(wires_370_5[1], addr_370_5, wires_1481_6,addr_1481_6);

wire[3:0] wires_1482_6;

wire[31:0] addr_1482_6;

Selector_2 s1482_6(wires_370_5[2], addr_370_5, wires_1482_6,addr_1482_6);

wire[3:0] wires_1483_6;

wire[31:0] addr_1483_6;

Selector_2 s1483_6(wires_370_5[3], addr_370_5, wires_1483_6,addr_1483_6);

wire[3:0] wires_1484_6;

wire[31:0] addr_1484_6;

Selector_2 s1484_6(wires_371_5[0], addr_371_5, wires_1484_6,addr_1484_6);

wire[3:0] wires_1485_6;

wire[31:0] addr_1485_6;

Selector_2 s1485_6(wires_371_5[1], addr_371_5, wires_1485_6,addr_1485_6);

wire[3:0] wires_1486_6;

wire[31:0] addr_1486_6;

Selector_2 s1486_6(wires_371_5[2], addr_371_5, wires_1486_6,addr_1486_6);

wire[3:0] wires_1487_6;

wire[31:0] addr_1487_6;

Selector_2 s1487_6(wires_371_5[3], addr_371_5, wires_1487_6,addr_1487_6);

wire[3:0] wires_1488_6;

wire[31:0] addr_1488_6;

Selector_2 s1488_6(wires_372_5[0], addr_372_5, wires_1488_6,addr_1488_6);

wire[3:0] wires_1489_6;

wire[31:0] addr_1489_6;

Selector_2 s1489_6(wires_372_5[1], addr_372_5, wires_1489_6,addr_1489_6);

wire[3:0] wires_1490_6;

wire[31:0] addr_1490_6;

Selector_2 s1490_6(wires_372_5[2], addr_372_5, wires_1490_6,addr_1490_6);

wire[3:0] wires_1491_6;

wire[31:0] addr_1491_6;

Selector_2 s1491_6(wires_372_5[3], addr_372_5, wires_1491_6,addr_1491_6);

wire[3:0] wires_1492_6;

wire[31:0] addr_1492_6;

Selector_2 s1492_6(wires_373_5[0], addr_373_5, wires_1492_6,addr_1492_6);

wire[3:0] wires_1493_6;

wire[31:0] addr_1493_6;

Selector_2 s1493_6(wires_373_5[1], addr_373_5, wires_1493_6,addr_1493_6);

wire[3:0] wires_1494_6;

wire[31:0] addr_1494_6;

Selector_2 s1494_6(wires_373_5[2], addr_373_5, wires_1494_6,addr_1494_6);

wire[3:0] wires_1495_6;

wire[31:0] addr_1495_6;

Selector_2 s1495_6(wires_373_5[3], addr_373_5, wires_1495_6,addr_1495_6);

wire[3:0] wires_1496_6;

wire[31:0] addr_1496_6;

Selector_2 s1496_6(wires_374_5[0], addr_374_5, wires_1496_6,addr_1496_6);

wire[3:0] wires_1497_6;

wire[31:0] addr_1497_6;

Selector_2 s1497_6(wires_374_5[1], addr_374_5, wires_1497_6,addr_1497_6);

wire[3:0] wires_1498_6;

wire[31:0] addr_1498_6;

Selector_2 s1498_6(wires_374_5[2], addr_374_5, wires_1498_6,addr_1498_6);

wire[3:0] wires_1499_6;

wire[31:0] addr_1499_6;

Selector_2 s1499_6(wires_374_5[3], addr_374_5, wires_1499_6,addr_1499_6);

wire[3:0] wires_1500_6;

wire[31:0] addr_1500_6;

Selector_2 s1500_6(wires_375_5[0], addr_375_5, wires_1500_6,addr_1500_6);

wire[3:0] wires_1501_6;

wire[31:0] addr_1501_6;

Selector_2 s1501_6(wires_375_5[1], addr_375_5, wires_1501_6,addr_1501_6);

wire[3:0] wires_1502_6;

wire[31:0] addr_1502_6;

Selector_2 s1502_6(wires_375_5[2], addr_375_5, wires_1502_6,addr_1502_6);

wire[3:0] wires_1503_6;

wire[31:0] addr_1503_6;

Selector_2 s1503_6(wires_375_5[3], addr_375_5, wires_1503_6,addr_1503_6);

wire[3:0] wires_1504_6;

wire[31:0] addr_1504_6;

Selector_2 s1504_6(wires_376_5[0], addr_376_5, wires_1504_6,addr_1504_6);

wire[3:0] wires_1505_6;

wire[31:0] addr_1505_6;

Selector_2 s1505_6(wires_376_5[1], addr_376_5, wires_1505_6,addr_1505_6);

wire[3:0] wires_1506_6;

wire[31:0] addr_1506_6;

Selector_2 s1506_6(wires_376_5[2], addr_376_5, wires_1506_6,addr_1506_6);

wire[3:0] wires_1507_6;

wire[31:0] addr_1507_6;

Selector_2 s1507_6(wires_376_5[3], addr_376_5, wires_1507_6,addr_1507_6);

wire[3:0] wires_1508_6;

wire[31:0] addr_1508_6;

Selector_2 s1508_6(wires_377_5[0], addr_377_5, wires_1508_6,addr_1508_6);

wire[3:0] wires_1509_6;

wire[31:0] addr_1509_6;

Selector_2 s1509_6(wires_377_5[1], addr_377_5, wires_1509_6,addr_1509_6);

wire[3:0] wires_1510_6;

wire[31:0] addr_1510_6;

Selector_2 s1510_6(wires_377_5[2], addr_377_5, wires_1510_6,addr_1510_6);

wire[3:0] wires_1511_6;

wire[31:0] addr_1511_6;

Selector_2 s1511_6(wires_377_5[3], addr_377_5, wires_1511_6,addr_1511_6);

wire[3:0] wires_1512_6;

wire[31:0] addr_1512_6;

Selector_2 s1512_6(wires_378_5[0], addr_378_5, wires_1512_6,addr_1512_6);

wire[3:0] wires_1513_6;

wire[31:0] addr_1513_6;

Selector_2 s1513_6(wires_378_5[1], addr_378_5, wires_1513_6,addr_1513_6);

wire[3:0] wires_1514_6;

wire[31:0] addr_1514_6;

Selector_2 s1514_6(wires_378_5[2], addr_378_5, wires_1514_6,addr_1514_6);

wire[3:0] wires_1515_6;

wire[31:0] addr_1515_6;

Selector_2 s1515_6(wires_378_5[3], addr_378_5, wires_1515_6,addr_1515_6);

wire[3:0] wires_1516_6;

wire[31:0] addr_1516_6;

Selector_2 s1516_6(wires_379_5[0], addr_379_5, wires_1516_6,addr_1516_6);

wire[3:0] wires_1517_6;

wire[31:0] addr_1517_6;

Selector_2 s1517_6(wires_379_5[1], addr_379_5, wires_1517_6,addr_1517_6);

wire[3:0] wires_1518_6;

wire[31:0] addr_1518_6;

Selector_2 s1518_6(wires_379_5[2], addr_379_5, wires_1518_6,addr_1518_6);

wire[3:0] wires_1519_6;

wire[31:0] addr_1519_6;

Selector_2 s1519_6(wires_379_5[3], addr_379_5, wires_1519_6,addr_1519_6);

wire[3:0] wires_1520_6;

wire[31:0] addr_1520_6;

Selector_2 s1520_6(wires_380_5[0], addr_380_5, wires_1520_6,addr_1520_6);

wire[3:0] wires_1521_6;

wire[31:0] addr_1521_6;

Selector_2 s1521_6(wires_380_5[1], addr_380_5, wires_1521_6,addr_1521_6);

wire[3:0] wires_1522_6;

wire[31:0] addr_1522_6;

Selector_2 s1522_6(wires_380_5[2], addr_380_5, wires_1522_6,addr_1522_6);

wire[3:0] wires_1523_6;

wire[31:0] addr_1523_6;

Selector_2 s1523_6(wires_380_5[3], addr_380_5, wires_1523_6,addr_1523_6);

wire[3:0] wires_1524_6;

wire[31:0] addr_1524_6;

Selector_2 s1524_6(wires_381_5[0], addr_381_5, wires_1524_6,addr_1524_6);

wire[3:0] wires_1525_6;

wire[31:0] addr_1525_6;

Selector_2 s1525_6(wires_381_5[1], addr_381_5, wires_1525_6,addr_1525_6);

wire[3:0] wires_1526_6;

wire[31:0] addr_1526_6;

Selector_2 s1526_6(wires_381_5[2], addr_381_5, wires_1526_6,addr_1526_6);

wire[3:0] wires_1527_6;

wire[31:0] addr_1527_6;

Selector_2 s1527_6(wires_381_5[3], addr_381_5, wires_1527_6,addr_1527_6);

wire[3:0] wires_1528_6;

wire[31:0] addr_1528_6;

Selector_2 s1528_6(wires_382_5[0], addr_382_5, wires_1528_6,addr_1528_6);

wire[3:0] wires_1529_6;

wire[31:0] addr_1529_6;

Selector_2 s1529_6(wires_382_5[1], addr_382_5, wires_1529_6,addr_1529_6);

wire[3:0] wires_1530_6;

wire[31:0] addr_1530_6;

Selector_2 s1530_6(wires_382_5[2], addr_382_5, wires_1530_6,addr_1530_6);

wire[3:0] wires_1531_6;

wire[31:0] addr_1531_6;

Selector_2 s1531_6(wires_382_5[3], addr_382_5, wires_1531_6,addr_1531_6);

wire[3:0] wires_1532_6;

wire[31:0] addr_1532_6;

Selector_2 s1532_6(wires_383_5[0], addr_383_5, wires_1532_6,addr_1532_6);

wire[3:0] wires_1533_6;

wire[31:0] addr_1533_6;

Selector_2 s1533_6(wires_383_5[1], addr_383_5, wires_1533_6,addr_1533_6);

wire[3:0] wires_1534_6;

wire[31:0] addr_1534_6;

Selector_2 s1534_6(wires_383_5[2], addr_383_5, wires_1534_6,addr_1534_6);

wire[3:0] wires_1535_6;

wire[31:0] addr_1535_6;

Selector_2 s1535_6(wires_383_5[3], addr_383_5, wires_1535_6,addr_1535_6);

wire[3:0] wires_1536_6;

wire[31:0] addr_1536_6;

Selector_2 s1536_6(wires_384_5[0], addr_384_5, wires_1536_6,addr_1536_6);

wire[3:0] wires_1537_6;

wire[31:0] addr_1537_6;

Selector_2 s1537_6(wires_384_5[1], addr_384_5, wires_1537_6,addr_1537_6);

wire[3:0] wires_1538_6;

wire[31:0] addr_1538_6;

Selector_2 s1538_6(wires_384_5[2], addr_384_5, wires_1538_6,addr_1538_6);

wire[3:0] wires_1539_6;

wire[31:0] addr_1539_6;

Selector_2 s1539_6(wires_384_5[3], addr_384_5, wires_1539_6,addr_1539_6);

wire[3:0] wires_1540_6;

wire[31:0] addr_1540_6;

Selector_2 s1540_6(wires_385_5[0], addr_385_5, wires_1540_6,addr_1540_6);

wire[3:0] wires_1541_6;

wire[31:0] addr_1541_6;

Selector_2 s1541_6(wires_385_5[1], addr_385_5, wires_1541_6,addr_1541_6);

wire[3:0] wires_1542_6;

wire[31:0] addr_1542_6;

Selector_2 s1542_6(wires_385_5[2], addr_385_5, wires_1542_6,addr_1542_6);

wire[3:0] wires_1543_6;

wire[31:0] addr_1543_6;

Selector_2 s1543_6(wires_385_5[3], addr_385_5, wires_1543_6,addr_1543_6);

wire[3:0] wires_1544_6;

wire[31:0] addr_1544_6;

Selector_2 s1544_6(wires_386_5[0], addr_386_5, wires_1544_6,addr_1544_6);

wire[3:0] wires_1545_6;

wire[31:0] addr_1545_6;

Selector_2 s1545_6(wires_386_5[1], addr_386_5, wires_1545_6,addr_1545_6);

wire[3:0] wires_1546_6;

wire[31:0] addr_1546_6;

Selector_2 s1546_6(wires_386_5[2], addr_386_5, wires_1546_6,addr_1546_6);

wire[3:0] wires_1547_6;

wire[31:0] addr_1547_6;

Selector_2 s1547_6(wires_386_5[3], addr_386_5, wires_1547_6,addr_1547_6);

wire[3:0] wires_1548_6;

wire[31:0] addr_1548_6;

Selector_2 s1548_6(wires_387_5[0], addr_387_5, wires_1548_6,addr_1548_6);

wire[3:0] wires_1549_6;

wire[31:0] addr_1549_6;

Selector_2 s1549_6(wires_387_5[1], addr_387_5, wires_1549_6,addr_1549_6);

wire[3:0] wires_1550_6;

wire[31:0] addr_1550_6;

Selector_2 s1550_6(wires_387_5[2], addr_387_5, wires_1550_6,addr_1550_6);

wire[3:0] wires_1551_6;

wire[31:0] addr_1551_6;

Selector_2 s1551_6(wires_387_5[3], addr_387_5, wires_1551_6,addr_1551_6);

wire[3:0] wires_1552_6;

wire[31:0] addr_1552_6;

Selector_2 s1552_6(wires_388_5[0], addr_388_5, wires_1552_6,addr_1552_6);

wire[3:0] wires_1553_6;

wire[31:0] addr_1553_6;

Selector_2 s1553_6(wires_388_5[1], addr_388_5, wires_1553_6,addr_1553_6);

wire[3:0] wires_1554_6;

wire[31:0] addr_1554_6;

Selector_2 s1554_6(wires_388_5[2], addr_388_5, wires_1554_6,addr_1554_6);

wire[3:0] wires_1555_6;

wire[31:0] addr_1555_6;

Selector_2 s1555_6(wires_388_5[3], addr_388_5, wires_1555_6,addr_1555_6);

wire[3:0] wires_1556_6;

wire[31:0] addr_1556_6;

Selector_2 s1556_6(wires_389_5[0], addr_389_5, wires_1556_6,addr_1556_6);

wire[3:0] wires_1557_6;

wire[31:0] addr_1557_6;

Selector_2 s1557_6(wires_389_5[1], addr_389_5, wires_1557_6,addr_1557_6);

wire[3:0] wires_1558_6;

wire[31:0] addr_1558_6;

Selector_2 s1558_6(wires_389_5[2], addr_389_5, wires_1558_6,addr_1558_6);

wire[3:0] wires_1559_6;

wire[31:0] addr_1559_6;

Selector_2 s1559_6(wires_389_5[3], addr_389_5, wires_1559_6,addr_1559_6);

wire[3:0] wires_1560_6;

wire[31:0] addr_1560_6;

Selector_2 s1560_6(wires_390_5[0], addr_390_5, wires_1560_6,addr_1560_6);

wire[3:0] wires_1561_6;

wire[31:0] addr_1561_6;

Selector_2 s1561_6(wires_390_5[1], addr_390_5, wires_1561_6,addr_1561_6);

wire[3:0] wires_1562_6;

wire[31:0] addr_1562_6;

Selector_2 s1562_6(wires_390_5[2], addr_390_5, wires_1562_6,addr_1562_6);

wire[3:0] wires_1563_6;

wire[31:0] addr_1563_6;

Selector_2 s1563_6(wires_390_5[3], addr_390_5, wires_1563_6,addr_1563_6);

wire[3:0] wires_1564_6;

wire[31:0] addr_1564_6;

Selector_2 s1564_6(wires_391_5[0], addr_391_5, wires_1564_6,addr_1564_6);

wire[3:0] wires_1565_6;

wire[31:0] addr_1565_6;

Selector_2 s1565_6(wires_391_5[1], addr_391_5, wires_1565_6,addr_1565_6);

wire[3:0] wires_1566_6;

wire[31:0] addr_1566_6;

Selector_2 s1566_6(wires_391_5[2], addr_391_5, wires_1566_6,addr_1566_6);

wire[3:0] wires_1567_6;

wire[31:0] addr_1567_6;

Selector_2 s1567_6(wires_391_5[3], addr_391_5, wires_1567_6,addr_1567_6);

wire[3:0] wires_1568_6;

wire[31:0] addr_1568_6;

Selector_2 s1568_6(wires_392_5[0], addr_392_5, wires_1568_6,addr_1568_6);

wire[3:0] wires_1569_6;

wire[31:0] addr_1569_6;

Selector_2 s1569_6(wires_392_5[1], addr_392_5, wires_1569_6,addr_1569_6);

wire[3:0] wires_1570_6;

wire[31:0] addr_1570_6;

Selector_2 s1570_6(wires_392_5[2], addr_392_5, wires_1570_6,addr_1570_6);

wire[3:0] wires_1571_6;

wire[31:0] addr_1571_6;

Selector_2 s1571_6(wires_392_5[3], addr_392_5, wires_1571_6,addr_1571_6);

wire[3:0] wires_1572_6;

wire[31:0] addr_1572_6;

Selector_2 s1572_6(wires_393_5[0], addr_393_5, wires_1572_6,addr_1572_6);

wire[3:0] wires_1573_6;

wire[31:0] addr_1573_6;

Selector_2 s1573_6(wires_393_5[1], addr_393_5, wires_1573_6,addr_1573_6);

wire[3:0] wires_1574_6;

wire[31:0] addr_1574_6;

Selector_2 s1574_6(wires_393_5[2], addr_393_5, wires_1574_6,addr_1574_6);

wire[3:0] wires_1575_6;

wire[31:0] addr_1575_6;

Selector_2 s1575_6(wires_393_5[3], addr_393_5, wires_1575_6,addr_1575_6);

wire[3:0] wires_1576_6;

wire[31:0] addr_1576_6;

Selector_2 s1576_6(wires_394_5[0], addr_394_5, wires_1576_6,addr_1576_6);

wire[3:0] wires_1577_6;

wire[31:0] addr_1577_6;

Selector_2 s1577_6(wires_394_5[1], addr_394_5, wires_1577_6,addr_1577_6);

wire[3:0] wires_1578_6;

wire[31:0] addr_1578_6;

Selector_2 s1578_6(wires_394_5[2], addr_394_5, wires_1578_6,addr_1578_6);

wire[3:0] wires_1579_6;

wire[31:0] addr_1579_6;

Selector_2 s1579_6(wires_394_5[3], addr_394_5, wires_1579_6,addr_1579_6);

wire[3:0] wires_1580_6;

wire[31:0] addr_1580_6;

Selector_2 s1580_6(wires_395_5[0], addr_395_5, wires_1580_6,addr_1580_6);

wire[3:0] wires_1581_6;

wire[31:0] addr_1581_6;

Selector_2 s1581_6(wires_395_5[1], addr_395_5, wires_1581_6,addr_1581_6);

wire[3:0] wires_1582_6;

wire[31:0] addr_1582_6;

Selector_2 s1582_6(wires_395_5[2], addr_395_5, wires_1582_6,addr_1582_6);

wire[3:0] wires_1583_6;

wire[31:0] addr_1583_6;

Selector_2 s1583_6(wires_395_5[3], addr_395_5, wires_1583_6,addr_1583_6);

wire[3:0] wires_1584_6;

wire[31:0] addr_1584_6;

Selector_2 s1584_6(wires_396_5[0], addr_396_5, wires_1584_6,addr_1584_6);

wire[3:0] wires_1585_6;

wire[31:0] addr_1585_6;

Selector_2 s1585_6(wires_396_5[1], addr_396_5, wires_1585_6,addr_1585_6);

wire[3:0] wires_1586_6;

wire[31:0] addr_1586_6;

Selector_2 s1586_6(wires_396_5[2], addr_396_5, wires_1586_6,addr_1586_6);

wire[3:0] wires_1587_6;

wire[31:0] addr_1587_6;

Selector_2 s1587_6(wires_396_5[3], addr_396_5, wires_1587_6,addr_1587_6);

wire[3:0] wires_1588_6;

wire[31:0] addr_1588_6;

Selector_2 s1588_6(wires_397_5[0], addr_397_5, wires_1588_6,addr_1588_6);

wire[3:0] wires_1589_6;

wire[31:0] addr_1589_6;

Selector_2 s1589_6(wires_397_5[1], addr_397_5, wires_1589_6,addr_1589_6);

wire[3:0] wires_1590_6;

wire[31:0] addr_1590_6;

Selector_2 s1590_6(wires_397_5[2], addr_397_5, wires_1590_6,addr_1590_6);

wire[3:0] wires_1591_6;

wire[31:0] addr_1591_6;

Selector_2 s1591_6(wires_397_5[3], addr_397_5, wires_1591_6,addr_1591_6);

wire[3:0] wires_1592_6;

wire[31:0] addr_1592_6;

Selector_2 s1592_6(wires_398_5[0], addr_398_5, wires_1592_6,addr_1592_6);

wire[3:0] wires_1593_6;

wire[31:0] addr_1593_6;

Selector_2 s1593_6(wires_398_5[1], addr_398_5, wires_1593_6,addr_1593_6);

wire[3:0] wires_1594_6;

wire[31:0] addr_1594_6;

Selector_2 s1594_6(wires_398_5[2], addr_398_5, wires_1594_6,addr_1594_6);

wire[3:0] wires_1595_6;

wire[31:0] addr_1595_6;

Selector_2 s1595_6(wires_398_5[3], addr_398_5, wires_1595_6,addr_1595_6);

wire[3:0] wires_1596_6;

wire[31:0] addr_1596_6;

Selector_2 s1596_6(wires_399_5[0], addr_399_5, wires_1596_6,addr_1596_6);

wire[3:0] wires_1597_6;

wire[31:0] addr_1597_6;

Selector_2 s1597_6(wires_399_5[1], addr_399_5, wires_1597_6,addr_1597_6);

wire[3:0] wires_1598_6;

wire[31:0] addr_1598_6;

Selector_2 s1598_6(wires_399_5[2], addr_399_5, wires_1598_6,addr_1598_6);

wire[3:0] wires_1599_6;

wire[31:0] addr_1599_6;

Selector_2 s1599_6(wires_399_5[3], addr_399_5, wires_1599_6,addr_1599_6);

wire[3:0] wires_1600_6;

wire[31:0] addr_1600_6;

Selector_2 s1600_6(wires_400_5[0], addr_400_5, wires_1600_6,addr_1600_6);

wire[3:0] wires_1601_6;

wire[31:0] addr_1601_6;

Selector_2 s1601_6(wires_400_5[1], addr_400_5, wires_1601_6,addr_1601_6);

wire[3:0] wires_1602_6;

wire[31:0] addr_1602_6;

Selector_2 s1602_6(wires_400_5[2], addr_400_5, wires_1602_6,addr_1602_6);

wire[3:0] wires_1603_6;

wire[31:0] addr_1603_6;

Selector_2 s1603_6(wires_400_5[3], addr_400_5, wires_1603_6,addr_1603_6);

wire[3:0] wires_1604_6;

wire[31:0] addr_1604_6;

Selector_2 s1604_6(wires_401_5[0], addr_401_5, wires_1604_6,addr_1604_6);

wire[3:0] wires_1605_6;

wire[31:0] addr_1605_6;

Selector_2 s1605_6(wires_401_5[1], addr_401_5, wires_1605_6,addr_1605_6);

wire[3:0] wires_1606_6;

wire[31:0] addr_1606_6;

Selector_2 s1606_6(wires_401_5[2], addr_401_5, wires_1606_6,addr_1606_6);

wire[3:0] wires_1607_6;

wire[31:0] addr_1607_6;

Selector_2 s1607_6(wires_401_5[3], addr_401_5, wires_1607_6,addr_1607_6);

wire[3:0] wires_1608_6;

wire[31:0] addr_1608_6;

Selector_2 s1608_6(wires_402_5[0], addr_402_5, wires_1608_6,addr_1608_6);

wire[3:0] wires_1609_6;

wire[31:0] addr_1609_6;

Selector_2 s1609_6(wires_402_5[1], addr_402_5, wires_1609_6,addr_1609_6);

wire[3:0] wires_1610_6;

wire[31:0] addr_1610_6;

Selector_2 s1610_6(wires_402_5[2], addr_402_5, wires_1610_6,addr_1610_6);

wire[3:0] wires_1611_6;

wire[31:0] addr_1611_6;

Selector_2 s1611_6(wires_402_5[3], addr_402_5, wires_1611_6,addr_1611_6);

wire[3:0] wires_1612_6;

wire[31:0] addr_1612_6;

Selector_2 s1612_6(wires_403_5[0], addr_403_5, wires_1612_6,addr_1612_6);

wire[3:0] wires_1613_6;

wire[31:0] addr_1613_6;

Selector_2 s1613_6(wires_403_5[1], addr_403_5, wires_1613_6,addr_1613_6);

wire[3:0] wires_1614_6;

wire[31:0] addr_1614_6;

Selector_2 s1614_6(wires_403_5[2], addr_403_5, wires_1614_6,addr_1614_6);

wire[3:0] wires_1615_6;

wire[31:0] addr_1615_6;

Selector_2 s1615_6(wires_403_5[3], addr_403_5, wires_1615_6,addr_1615_6);

wire[3:0] wires_1616_6;

wire[31:0] addr_1616_6;

Selector_2 s1616_6(wires_404_5[0], addr_404_5, wires_1616_6,addr_1616_6);

wire[3:0] wires_1617_6;

wire[31:0] addr_1617_6;

Selector_2 s1617_6(wires_404_5[1], addr_404_5, wires_1617_6,addr_1617_6);

wire[3:0] wires_1618_6;

wire[31:0] addr_1618_6;

Selector_2 s1618_6(wires_404_5[2], addr_404_5, wires_1618_6,addr_1618_6);

wire[3:0] wires_1619_6;

wire[31:0] addr_1619_6;

Selector_2 s1619_6(wires_404_5[3], addr_404_5, wires_1619_6,addr_1619_6);

wire[3:0] wires_1620_6;

wire[31:0] addr_1620_6;

Selector_2 s1620_6(wires_405_5[0], addr_405_5, wires_1620_6,addr_1620_6);

wire[3:0] wires_1621_6;

wire[31:0] addr_1621_6;

Selector_2 s1621_6(wires_405_5[1], addr_405_5, wires_1621_6,addr_1621_6);

wire[3:0] wires_1622_6;

wire[31:0] addr_1622_6;

Selector_2 s1622_6(wires_405_5[2], addr_405_5, wires_1622_6,addr_1622_6);

wire[3:0] wires_1623_6;

wire[31:0] addr_1623_6;

Selector_2 s1623_6(wires_405_5[3], addr_405_5, wires_1623_6,addr_1623_6);

wire[3:0] wires_1624_6;

wire[31:0] addr_1624_6;

Selector_2 s1624_6(wires_406_5[0], addr_406_5, wires_1624_6,addr_1624_6);

wire[3:0] wires_1625_6;

wire[31:0] addr_1625_6;

Selector_2 s1625_6(wires_406_5[1], addr_406_5, wires_1625_6,addr_1625_6);

wire[3:0] wires_1626_6;

wire[31:0] addr_1626_6;

Selector_2 s1626_6(wires_406_5[2], addr_406_5, wires_1626_6,addr_1626_6);

wire[3:0] wires_1627_6;

wire[31:0] addr_1627_6;

Selector_2 s1627_6(wires_406_5[3], addr_406_5, wires_1627_6,addr_1627_6);

wire[3:0] wires_1628_6;

wire[31:0] addr_1628_6;

Selector_2 s1628_6(wires_407_5[0], addr_407_5, wires_1628_6,addr_1628_6);

wire[3:0] wires_1629_6;

wire[31:0] addr_1629_6;

Selector_2 s1629_6(wires_407_5[1], addr_407_5, wires_1629_6,addr_1629_6);

wire[3:0] wires_1630_6;

wire[31:0] addr_1630_6;

Selector_2 s1630_6(wires_407_5[2], addr_407_5, wires_1630_6,addr_1630_6);

wire[3:0] wires_1631_6;

wire[31:0] addr_1631_6;

Selector_2 s1631_6(wires_407_5[3], addr_407_5, wires_1631_6,addr_1631_6);

wire[3:0] wires_1632_6;

wire[31:0] addr_1632_6;

Selector_2 s1632_6(wires_408_5[0], addr_408_5, wires_1632_6,addr_1632_6);

wire[3:0] wires_1633_6;

wire[31:0] addr_1633_6;

Selector_2 s1633_6(wires_408_5[1], addr_408_5, wires_1633_6,addr_1633_6);

wire[3:0] wires_1634_6;

wire[31:0] addr_1634_6;

Selector_2 s1634_6(wires_408_5[2], addr_408_5, wires_1634_6,addr_1634_6);

wire[3:0] wires_1635_6;

wire[31:0] addr_1635_6;

Selector_2 s1635_6(wires_408_5[3], addr_408_5, wires_1635_6,addr_1635_6);

wire[3:0] wires_1636_6;

wire[31:0] addr_1636_6;

Selector_2 s1636_6(wires_409_5[0], addr_409_5, wires_1636_6,addr_1636_6);

wire[3:0] wires_1637_6;

wire[31:0] addr_1637_6;

Selector_2 s1637_6(wires_409_5[1], addr_409_5, wires_1637_6,addr_1637_6);

wire[3:0] wires_1638_6;

wire[31:0] addr_1638_6;

Selector_2 s1638_6(wires_409_5[2], addr_409_5, wires_1638_6,addr_1638_6);

wire[3:0] wires_1639_6;

wire[31:0] addr_1639_6;

Selector_2 s1639_6(wires_409_5[3], addr_409_5, wires_1639_6,addr_1639_6);

wire[3:0] wires_1640_6;

wire[31:0] addr_1640_6;

Selector_2 s1640_6(wires_410_5[0], addr_410_5, wires_1640_6,addr_1640_6);

wire[3:0] wires_1641_6;

wire[31:0] addr_1641_6;

Selector_2 s1641_6(wires_410_5[1], addr_410_5, wires_1641_6,addr_1641_6);

wire[3:0] wires_1642_6;

wire[31:0] addr_1642_6;

Selector_2 s1642_6(wires_410_5[2], addr_410_5, wires_1642_6,addr_1642_6);

wire[3:0] wires_1643_6;

wire[31:0] addr_1643_6;

Selector_2 s1643_6(wires_410_5[3], addr_410_5, wires_1643_6,addr_1643_6);

wire[3:0] wires_1644_6;

wire[31:0] addr_1644_6;

Selector_2 s1644_6(wires_411_5[0], addr_411_5, wires_1644_6,addr_1644_6);

wire[3:0] wires_1645_6;

wire[31:0] addr_1645_6;

Selector_2 s1645_6(wires_411_5[1], addr_411_5, wires_1645_6,addr_1645_6);

wire[3:0] wires_1646_6;

wire[31:0] addr_1646_6;

Selector_2 s1646_6(wires_411_5[2], addr_411_5, wires_1646_6,addr_1646_6);

wire[3:0] wires_1647_6;

wire[31:0] addr_1647_6;

Selector_2 s1647_6(wires_411_5[3], addr_411_5, wires_1647_6,addr_1647_6);

wire[3:0] wires_1648_6;

wire[31:0] addr_1648_6;

Selector_2 s1648_6(wires_412_5[0], addr_412_5, wires_1648_6,addr_1648_6);

wire[3:0] wires_1649_6;

wire[31:0] addr_1649_6;

Selector_2 s1649_6(wires_412_5[1], addr_412_5, wires_1649_6,addr_1649_6);

wire[3:0] wires_1650_6;

wire[31:0] addr_1650_6;

Selector_2 s1650_6(wires_412_5[2], addr_412_5, wires_1650_6,addr_1650_6);

wire[3:0] wires_1651_6;

wire[31:0] addr_1651_6;

Selector_2 s1651_6(wires_412_5[3], addr_412_5, wires_1651_6,addr_1651_6);

wire[3:0] wires_1652_6;

wire[31:0] addr_1652_6;

Selector_2 s1652_6(wires_413_5[0], addr_413_5, wires_1652_6,addr_1652_6);

wire[3:0] wires_1653_6;

wire[31:0] addr_1653_6;

Selector_2 s1653_6(wires_413_5[1], addr_413_5, wires_1653_6,addr_1653_6);

wire[3:0] wires_1654_6;

wire[31:0] addr_1654_6;

Selector_2 s1654_6(wires_413_5[2], addr_413_5, wires_1654_6,addr_1654_6);

wire[3:0] wires_1655_6;

wire[31:0] addr_1655_6;

Selector_2 s1655_6(wires_413_5[3], addr_413_5, wires_1655_6,addr_1655_6);

wire[3:0] wires_1656_6;

wire[31:0] addr_1656_6;

Selector_2 s1656_6(wires_414_5[0], addr_414_5, wires_1656_6,addr_1656_6);

wire[3:0] wires_1657_6;

wire[31:0] addr_1657_6;

Selector_2 s1657_6(wires_414_5[1], addr_414_5, wires_1657_6,addr_1657_6);

wire[3:0] wires_1658_6;

wire[31:0] addr_1658_6;

Selector_2 s1658_6(wires_414_5[2], addr_414_5, wires_1658_6,addr_1658_6);

wire[3:0] wires_1659_6;

wire[31:0] addr_1659_6;

Selector_2 s1659_6(wires_414_5[3], addr_414_5, wires_1659_6,addr_1659_6);

wire[3:0] wires_1660_6;

wire[31:0] addr_1660_6;

Selector_2 s1660_6(wires_415_5[0], addr_415_5, wires_1660_6,addr_1660_6);

wire[3:0] wires_1661_6;

wire[31:0] addr_1661_6;

Selector_2 s1661_6(wires_415_5[1], addr_415_5, wires_1661_6,addr_1661_6);

wire[3:0] wires_1662_6;

wire[31:0] addr_1662_6;

Selector_2 s1662_6(wires_415_5[2], addr_415_5, wires_1662_6,addr_1662_6);

wire[3:0] wires_1663_6;

wire[31:0] addr_1663_6;

Selector_2 s1663_6(wires_415_5[3], addr_415_5, wires_1663_6,addr_1663_6);

wire[3:0] wires_1664_6;

wire[31:0] addr_1664_6;

Selector_2 s1664_6(wires_416_5[0], addr_416_5, wires_1664_6,addr_1664_6);

wire[3:0] wires_1665_6;

wire[31:0] addr_1665_6;

Selector_2 s1665_6(wires_416_5[1], addr_416_5, wires_1665_6,addr_1665_6);

wire[3:0] wires_1666_6;

wire[31:0] addr_1666_6;

Selector_2 s1666_6(wires_416_5[2], addr_416_5, wires_1666_6,addr_1666_6);

wire[3:0] wires_1667_6;

wire[31:0] addr_1667_6;

Selector_2 s1667_6(wires_416_5[3], addr_416_5, wires_1667_6,addr_1667_6);

wire[3:0] wires_1668_6;

wire[31:0] addr_1668_6;

Selector_2 s1668_6(wires_417_5[0], addr_417_5, wires_1668_6,addr_1668_6);

wire[3:0] wires_1669_6;

wire[31:0] addr_1669_6;

Selector_2 s1669_6(wires_417_5[1], addr_417_5, wires_1669_6,addr_1669_6);

wire[3:0] wires_1670_6;

wire[31:0] addr_1670_6;

Selector_2 s1670_6(wires_417_5[2], addr_417_5, wires_1670_6,addr_1670_6);

wire[3:0] wires_1671_6;

wire[31:0] addr_1671_6;

Selector_2 s1671_6(wires_417_5[3], addr_417_5, wires_1671_6,addr_1671_6);

wire[3:0] wires_1672_6;

wire[31:0] addr_1672_6;

Selector_2 s1672_6(wires_418_5[0], addr_418_5, wires_1672_6,addr_1672_6);

wire[3:0] wires_1673_6;

wire[31:0] addr_1673_6;

Selector_2 s1673_6(wires_418_5[1], addr_418_5, wires_1673_6,addr_1673_6);

wire[3:0] wires_1674_6;

wire[31:0] addr_1674_6;

Selector_2 s1674_6(wires_418_5[2], addr_418_5, wires_1674_6,addr_1674_6);

wire[3:0] wires_1675_6;

wire[31:0] addr_1675_6;

Selector_2 s1675_6(wires_418_5[3], addr_418_5, wires_1675_6,addr_1675_6);

wire[3:0] wires_1676_6;

wire[31:0] addr_1676_6;

Selector_2 s1676_6(wires_419_5[0], addr_419_5, wires_1676_6,addr_1676_6);

wire[3:0] wires_1677_6;

wire[31:0] addr_1677_6;

Selector_2 s1677_6(wires_419_5[1], addr_419_5, wires_1677_6,addr_1677_6);

wire[3:0] wires_1678_6;

wire[31:0] addr_1678_6;

Selector_2 s1678_6(wires_419_5[2], addr_419_5, wires_1678_6,addr_1678_6);

wire[3:0] wires_1679_6;

wire[31:0] addr_1679_6;

Selector_2 s1679_6(wires_419_5[3], addr_419_5, wires_1679_6,addr_1679_6);

wire[3:0] wires_1680_6;

wire[31:0] addr_1680_6;

Selector_2 s1680_6(wires_420_5[0], addr_420_5, wires_1680_6,addr_1680_6);

wire[3:0] wires_1681_6;

wire[31:0] addr_1681_6;

Selector_2 s1681_6(wires_420_5[1], addr_420_5, wires_1681_6,addr_1681_6);

wire[3:0] wires_1682_6;

wire[31:0] addr_1682_6;

Selector_2 s1682_6(wires_420_5[2], addr_420_5, wires_1682_6,addr_1682_6);

wire[3:0] wires_1683_6;

wire[31:0] addr_1683_6;

Selector_2 s1683_6(wires_420_5[3], addr_420_5, wires_1683_6,addr_1683_6);

wire[3:0] wires_1684_6;

wire[31:0] addr_1684_6;

Selector_2 s1684_6(wires_421_5[0], addr_421_5, wires_1684_6,addr_1684_6);

wire[3:0] wires_1685_6;

wire[31:0] addr_1685_6;

Selector_2 s1685_6(wires_421_5[1], addr_421_5, wires_1685_6,addr_1685_6);

wire[3:0] wires_1686_6;

wire[31:0] addr_1686_6;

Selector_2 s1686_6(wires_421_5[2], addr_421_5, wires_1686_6,addr_1686_6);

wire[3:0] wires_1687_6;

wire[31:0] addr_1687_6;

Selector_2 s1687_6(wires_421_5[3], addr_421_5, wires_1687_6,addr_1687_6);

wire[3:0] wires_1688_6;

wire[31:0] addr_1688_6;

Selector_2 s1688_6(wires_422_5[0], addr_422_5, wires_1688_6,addr_1688_6);

wire[3:0] wires_1689_6;

wire[31:0] addr_1689_6;

Selector_2 s1689_6(wires_422_5[1], addr_422_5, wires_1689_6,addr_1689_6);

wire[3:0] wires_1690_6;

wire[31:0] addr_1690_6;

Selector_2 s1690_6(wires_422_5[2], addr_422_5, wires_1690_6,addr_1690_6);

wire[3:0] wires_1691_6;

wire[31:0] addr_1691_6;

Selector_2 s1691_6(wires_422_5[3], addr_422_5, wires_1691_6,addr_1691_6);

wire[3:0] wires_1692_6;

wire[31:0] addr_1692_6;

Selector_2 s1692_6(wires_423_5[0], addr_423_5, wires_1692_6,addr_1692_6);

wire[3:0] wires_1693_6;

wire[31:0] addr_1693_6;

Selector_2 s1693_6(wires_423_5[1], addr_423_5, wires_1693_6,addr_1693_6);

wire[3:0] wires_1694_6;

wire[31:0] addr_1694_6;

Selector_2 s1694_6(wires_423_5[2], addr_423_5, wires_1694_6,addr_1694_6);

wire[3:0] wires_1695_6;

wire[31:0] addr_1695_6;

Selector_2 s1695_6(wires_423_5[3], addr_423_5, wires_1695_6,addr_1695_6);

wire[3:0] wires_1696_6;

wire[31:0] addr_1696_6;

Selector_2 s1696_6(wires_424_5[0], addr_424_5, wires_1696_6,addr_1696_6);

wire[3:0] wires_1697_6;

wire[31:0] addr_1697_6;

Selector_2 s1697_6(wires_424_5[1], addr_424_5, wires_1697_6,addr_1697_6);

wire[3:0] wires_1698_6;

wire[31:0] addr_1698_6;

Selector_2 s1698_6(wires_424_5[2], addr_424_5, wires_1698_6,addr_1698_6);

wire[3:0] wires_1699_6;

wire[31:0] addr_1699_6;

Selector_2 s1699_6(wires_424_5[3], addr_424_5, wires_1699_6,addr_1699_6);

wire[3:0] wires_1700_6;

wire[31:0] addr_1700_6;

Selector_2 s1700_6(wires_425_5[0], addr_425_5, wires_1700_6,addr_1700_6);

wire[3:0] wires_1701_6;

wire[31:0] addr_1701_6;

Selector_2 s1701_6(wires_425_5[1], addr_425_5, wires_1701_6,addr_1701_6);

wire[3:0] wires_1702_6;

wire[31:0] addr_1702_6;

Selector_2 s1702_6(wires_425_5[2], addr_425_5, wires_1702_6,addr_1702_6);

wire[3:0] wires_1703_6;

wire[31:0] addr_1703_6;

Selector_2 s1703_6(wires_425_5[3], addr_425_5, wires_1703_6,addr_1703_6);

wire[3:0] wires_1704_6;

wire[31:0] addr_1704_6;

Selector_2 s1704_6(wires_426_5[0], addr_426_5, wires_1704_6,addr_1704_6);

wire[3:0] wires_1705_6;

wire[31:0] addr_1705_6;

Selector_2 s1705_6(wires_426_5[1], addr_426_5, wires_1705_6,addr_1705_6);

wire[3:0] wires_1706_6;

wire[31:0] addr_1706_6;

Selector_2 s1706_6(wires_426_5[2], addr_426_5, wires_1706_6,addr_1706_6);

wire[3:0] wires_1707_6;

wire[31:0] addr_1707_6;

Selector_2 s1707_6(wires_426_5[3], addr_426_5, wires_1707_6,addr_1707_6);

wire[3:0] wires_1708_6;

wire[31:0] addr_1708_6;

Selector_2 s1708_6(wires_427_5[0], addr_427_5, wires_1708_6,addr_1708_6);

wire[3:0] wires_1709_6;

wire[31:0] addr_1709_6;

Selector_2 s1709_6(wires_427_5[1], addr_427_5, wires_1709_6,addr_1709_6);

wire[3:0] wires_1710_6;

wire[31:0] addr_1710_6;

Selector_2 s1710_6(wires_427_5[2], addr_427_5, wires_1710_6,addr_1710_6);

wire[3:0] wires_1711_6;

wire[31:0] addr_1711_6;

Selector_2 s1711_6(wires_427_5[3], addr_427_5, wires_1711_6,addr_1711_6);

wire[3:0] wires_1712_6;

wire[31:0] addr_1712_6;

Selector_2 s1712_6(wires_428_5[0], addr_428_5, wires_1712_6,addr_1712_6);

wire[3:0] wires_1713_6;

wire[31:0] addr_1713_6;

Selector_2 s1713_6(wires_428_5[1], addr_428_5, wires_1713_6,addr_1713_6);

wire[3:0] wires_1714_6;

wire[31:0] addr_1714_6;

Selector_2 s1714_6(wires_428_5[2], addr_428_5, wires_1714_6,addr_1714_6);

wire[3:0] wires_1715_6;

wire[31:0] addr_1715_6;

Selector_2 s1715_6(wires_428_5[3], addr_428_5, wires_1715_6,addr_1715_6);

wire[3:0] wires_1716_6;

wire[31:0] addr_1716_6;

Selector_2 s1716_6(wires_429_5[0], addr_429_5, wires_1716_6,addr_1716_6);

wire[3:0] wires_1717_6;

wire[31:0] addr_1717_6;

Selector_2 s1717_6(wires_429_5[1], addr_429_5, wires_1717_6,addr_1717_6);

wire[3:0] wires_1718_6;

wire[31:0] addr_1718_6;

Selector_2 s1718_6(wires_429_5[2], addr_429_5, wires_1718_6,addr_1718_6);

wire[3:0] wires_1719_6;

wire[31:0] addr_1719_6;

Selector_2 s1719_6(wires_429_5[3], addr_429_5, wires_1719_6,addr_1719_6);

wire[3:0] wires_1720_6;

wire[31:0] addr_1720_6;

Selector_2 s1720_6(wires_430_5[0], addr_430_5, wires_1720_6,addr_1720_6);

wire[3:0] wires_1721_6;

wire[31:0] addr_1721_6;

Selector_2 s1721_6(wires_430_5[1], addr_430_5, wires_1721_6,addr_1721_6);

wire[3:0] wires_1722_6;

wire[31:0] addr_1722_6;

Selector_2 s1722_6(wires_430_5[2], addr_430_5, wires_1722_6,addr_1722_6);

wire[3:0] wires_1723_6;

wire[31:0] addr_1723_6;

Selector_2 s1723_6(wires_430_5[3], addr_430_5, wires_1723_6,addr_1723_6);

wire[3:0] wires_1724_6;

wire[31:0] addr_1724_6;

Selector_2 s1724_6(wires_431_5[0], addr_431_5, wires_1724_6,addr_1724_6);

wire[3:0] wires_1725_6;

wire[31:0] addr_1725_6;

Selector_2 s1725_6(wires_431_5[1], addr_431_5, wires_1725_6,addr_1725_6);

wire[3:0] wires_1726_6;

wire[31:0] addr_1726_6;

Selector_2 s1726_6(wires_431_5[2], addr_431_5, wires_1726_6,addr_1726_6);

wire[3:0] wires_1727_6;

wire[31:0] addr_1727_6;

Selector_2 s1727_6(wires_431_5[3], addr_431_5, wires_1727_6,addr_1727_6);

wire[3:0] wires_1728_6;

wire[31:0] addr_1728_6;

Selector_2 s1728_6(wires_432_5[0], addr_432_5, wires_1728_6,addr_1728_6);

wire[3:0] wires_1729_6;

wire[31:0] addr_1729_6;

Selector_2 s1729_6(wires_432_5[1], addr_432_5, wires_1729_6,addr_1729_6);

wire[3:0] wires_1730_6;

wire[31:0] addr_1730_6;

Selector_2 s1730_6(wires_432_5[2], addr_432_5, wires_1730_6,addr_1730_6);

wire[3:0] wires_1731_6;

wire[31:0] addr_1731_6;

Selector_2 s1731_6(wires_432_5[3], addr_432_5, wires_1731_6,addr_1731_6);

wire[3:0] wires_1732_6;

wire[31:0] addr_1732_6;

Selector_2 s1732_6(wires_433_5[0], addr_433_5, wires_1732_6,addr_1732_6);

wire[3:0] wires_1733_6;

wire[31:0] addr_1733_6;

Selector_2 s1733_6(wires_433_5[1], addr_433_5, wires_1733_6,addr_1733_6);

wire[3:0] wires_1734_6;

wire[31:0] addr_1734_6;

Selector_2 s1734_6(wires_433_5[2], addr_433_5, wires_1734_6,addr_1734_6);

wire[3:0] wires_1735_6;

wire[31:0] addr_1735_6;

Selector_2 s1735_6(wires_433_5[3], addr_433_5, wires_1735_6,addr_1735_6);

wire[3:0] wires_1736_6;

wire[31:0] addr_1736_6;

Selector_2 s1736_6(wires_434_5[0], addr_434_5, wires_1736_6,addr_1736_6);

wire[3:0] wires_1737_6;

wire[31:0] addr_1737_6;

Selector_2 s1737_6(wires_434_5[1], addr_434_5, wires_1737_6,addr_1737_6);

wire[3:0] wires_1738_6;

wire[31:0] addr_1738_6;

Selector_2 s1738_6(wires_434_5[2], addr_434_5, wires_1738_6,addr_1738_6);

wire[3:0] wires_1739_6;

wire[31:0] addr_1739_6;

Selector_2 s1739_6(wires_434_5[3], addr_434_5, wires_1739_6,addr_1739_6);

wire[3:0] wires_1740_6;

wire[31:0] addr_1740_6;

Selector_2 s1740_6(wires_435_5[0], addr_435_5, wires_1740_6,addr_1740_6);

wire[3:0] wires_1741_6;

wire[31:0] addr_1741_6;

Selector_2 s1741_6(wires_435_5[1], addr_435_5, wires_1741_6,addr_1741_6);

wire[3:0] wires_1742_6;

wire[31:0] addr_1742_6;

Selector_2 s1742_6(wires_435_5[2], addr_435_5, wires_1742_6,addr_1742_6);

wire[3:0] wires_1743_6;

wire[31:0] addr_1743_6;

Selector_2 s1743_6(wires_435_5[3], addr_435_5, wires_1743_6,addr_1743_6);

wire[3:0] wires_1744_6;

wire[31:0] addr_1744_6;

Selector_2 s1744_6(wires_436_5[0], addr_436_5, wires_1744_6,addr_1744_6);

wire[3:0] wires_1745_6;

wire[31:0] addr_1745_6;

Selector_2 s1745_6(wires_436_5[1], addr_436_5, wires_1745_6,addr_1745_6);

wire[3:0] wires_1746_6;

wire[31:0] addr_1746_6;

Selector_2 s1746_6(wires_436_5[2], addr_436_5, wires_1746_6,addr_1746_6);

wire[3:0] wires_1747_6;

wire[31:0] addr_1747_6;

Selector_2 s1747_6(wires_436_5[3], addr_436_5, wires_1747_6,addr_1747_6);

wire[3:0] wires_1748_6;

wire[31:0] addr_1748_6;

Selector_2 s1748_6(wires_437_5[0], addr_437_5, wires_1748_6,addr_1748_6);

wire[3:0] wires_1749_6;

wire[31:0] addr_1749_6;

Selector_2 s1749_6(wires_437_5[1], addr_437_5, wires_1749_6,addr_1749_6);

wire[3:0] wires_1750_6;

wire[31:0] addr_1750_6;

Selector_2 s1750_6(wires_437_5[2], addr_437_5, wires_1750_6,addr_1750_6);

wire[3:0] wires_1751_6;

wire[31:0] addr_1751_6;

Selector_2 s1751_6(wires_437_5[3], addr_437_5, wires_1751_6,addr_1751_6);

wire[3:0] wires_1752_6;

wire[31:0] addr_1752_6;

Selector_2 s1752_6(wires_438_5[0], addr_438_5, wires_1752_6,addr_1752_6);

wire[3:0] wires_1753_6;

wire[31:0] addr_1753_6;

Selector_2 s1753_6(wires_438_5[1], addr_438_5, wires_1753_6,addr_1753_6);

wire[3:0] wires_1754_6;

wire[31:0] addr_1754_6;

Selector_2 s1754_6(wires_438_5[2], addr_438_5, wires_1754_6,addr_1754_6);

wire[3:0] wires_1755_6;

wire[31:0] addr_1755_6;

Selector_2 s1755_6(wires_438_5[3], addr_438_5, wires_1755_6,addr_1755_6);

wire[3:0] wires_1756_6;

wire[31:0] addr_1756_6;

Selector_2 s1756_6(wires_439_5[0], addr_439_5, wires_1756_6,addr_1756_6);

wire[3:0] wires_1757_6;

wire[31:0] addr_1757_6;

Selector_2 s1757_6(wires_439_5[1], addr_439_5, wires_1757_6,addr_1757_6);

wire[3:0] wires_1758_6;

wire[31:0] addr_1758_6;

Selector_2 s1758_6(wires_439_5[2], addr_439_5, wires_1758_6,addr_1758_6);

wire[3:0] wires_1759_6;

wire[31:0] addr_1759_6;

Selector_2 s1759_6(wires_439_5[3], addr_439_5, wires_1759_6,addr_1759_6);

wire[3:0] wires_1760_6;

wire[31:0] addr_1760_6;

Selector_2 s1760_6(wires_440_5[0], addr_440_5, wires_1760_6,addr_1760_6);

wire[3:0] wires_1761_6;

wire[31:0] addr_1761_6;

Selector_2 s1761_6(wires_440_5[1], addr_440_5, wires_1761_6,addr_1761_6);

wire[3:0] wires_1762_6;

wire[31:0] addr_1762_6;

Selector_2 s1762_6(wires_440_5[2], addr_440_5, wires_1762_6,addr_1762_6);

wire[3:0] wires_1763_6;

wire[31:0] addr_1763_6;

Selector_2 s1763_6(wires_440_5[3], addr_440_5, wires_1763_6,addr_1763_6);

wire[3:0] wires_1764_6;

wire[31:0] addr_1764_6;

Selector_2 s1764_6(wires_441_5[0], addr_441_5, wires_1764_6,addr_1764_6);

wire[3:0] wires_1765_6;

wire[31:0] addr_1765_6;

Selector_2 s1765_6(wires_441_5[1], addr_441_5, wires_1765_6,addr_1765_6);

wire[3:0] wires_1766_6;

wire[31:0] addr_1766_6;

Selector_2 s1766_6(wires_441_5[2], addr_441_5, wires_1766_6,addr_1766_6);

wire[3:0] wires_1767_6;

wire[31:0] addr_1767_6;

Selector_2 s1767_6(wires_441_5[3], addr_441_5, wires_1767_6,addr_1767_6);

wire[3:0] wires_1768_6;

wire[31:0] addr_1768_6;

Selector_2 s1768_6(wires_442_5[0], addr_442_5, wires_1768_6,addr_1768_6);

wire[3:0] wires_1769_6;

wire[31:0] addr_1769_6;

Selector_2 s1769_6(wires_442_5[1], addr_442_5, wires_1769_6,addr_1769_6);

wire[3:0] wires_1770_6;

wire[31:0] addr_1770_6;

Selector_2 s1770_6(wires_442_5[2], addr_442_5, wires_1770_6,addr_1770_6);

wire[3:0] wires_1771_6;

wire[31:0] addr_1771_6;

Selector_2 s1771_6(wires_442_5[3], addr_442_5, wires_1771_6,addr_1771_6);

wire[3:0] wires_1772_6;

wire[31:0] addr_1772_6;

Selector_2 s1772_6(wires_443_5[0], addr_443_5, wires_1772_6,addr_1772_6);

wire[3:0] wires_1773_6;

wire[31:0] addr_1773_6;

Selector_2 s1773_6(wires_443_5[1], addr_443_5, wires_1773_6,addr_1773_6);

wire[3:0] wires_1774_6;

wire[31:0] addr_1774_6;

Selector_2 s1774_6(wires_443_5[2], addr_443_5, wires_1774_6,addr_1774_6);

wire[3:0] wires_1775_6;

wire[31:0] addr_1775_6;

Selector_2 s1775_6(wires_443_5[3], addr_443_5, wires_1775_6,addr_1775_6);

wire[3:0] wires_1776_6;

wire[31:0] addr_1776_6;

Selector_2 s1776_6(wires_444_5[0], addr_444_5, wires_1776_6,addr_1776_6);

wire[3:0] wires_1777_6;

wire[31:0] addr_1777_6;

Selector_2 s1777_6(wires_444_5[1], addr_444_5, wires_1777_6,addr_1777_6);

wire[3:0] wires_1778_6;

wire[31:0] addr_1778_6;

Selector_2 s1778_6(wires_444_5[2], addr_444_5, wires_1778_6,addr_1778_6);

wire[3:0] wires_1779_6;

wire[31:0] addr_1779_6;

Selector_2 s1779_6(wires_444_5[3], addr_444_5, wires_1779_6,addr_1779_6);

wire[3:0] wires_1780_6;

wire[31:0] addr_1780_6;

Selector_2 s1780_6(wires_445_5[0], addr_445_5, wires_1780_6,addr_1780_6);

wire[3:0] wires_1781_6;

wire[31:0] addr_1781_6;

Selector_2 s1781_6(wires_445_5[1], addr_445_5, wires_1781_6,addr_1781_6);

wire[3:0] wires_1782_6;

wire[31:0] addr_1782_6;

Selector_2 s1782_6(wires_445_5[2], addr_445_5, wires_1782_6,addr_1782_6);

wire[3:0] wires_1783_6;

wire[31:0] addr_1783_6;

Selector_2 s1783_6(wires_445_5[3], addr_445_5, wires_1783_6,addr_1783_6);

wire[3:0] wires_1784_6;

wire[31:0] addr_1784_6;

Selector_2 s1784_6(wires_446_5[0], addr_446_5, wires_1784_6,addr_1784_6);

wire[3:0] wires_1785_6;

wire[31:0] addr_1785_6;

Selector_2 s1785_6(wires_446_5[1], addr_446_5, wires_1785_6,addr_1785_6);

wire[3:0] wires_1786_6;

wire[31:0] addr_1786_6;

Selector_2 s1786_6(wires_446_5[2], addr_446_5, wires_1786_6,addr_1786_6);

wire[3:0] wires_1787_6;

wire[31:0] addr_1787_6;

Selector_2 s1787_6(wires_446_5[3], addr_446_5, wires_1787_6,addr_1787_6);

wire[3:0] wires_1788_6;

wire[31:0] addr_1788_6;

Selector_2 s1788_6(wires_447_5[0], addr_447_5, wires_1788_6,addr_1788_6);

wire[3:0] wires_1789_6;

wire[31:0] addr_1789_6;

Selector_2 s1789_6(wires_447_5[1], addr_447_5, wires_1789_6,addr_1789_6);

wire[3:0] wires_1790_6;

wire[31:0] addr_1790_6;

Selector_2 s1790_6(wires_447_5[2], addr_447_5, wires_1790_6,addr_1790_6);

wire[3:0] wires_1791_6;

wire[31:0] addr_1791_6;

Selector_2 s1791_6(wires_447_5[3], addr_447_5, wires_1791_6,addr_1791_6);

wire[3:0] wires_1792_6;

wire[31:0] addr_1792_6;

Selector_2 s1792_6(wires_448_5[0], addr_448_5, wires_1792_6,addr_1792_6);

wire[3:0] wires_1793_6;

wire[31:0] addr_1793_6;

Selector_2 s1793_6(wires_448_5[1], addr_448_5, wires_1793_6,addr_1793_6);

wire[3:0] wires_1794_6;

wire[31:0] addr_1794_6;

Selector_2 s1794_6(wires_448_5[2], addr_448_5, wires_1794_6,addr_1794_6);

wire[3:0] wires_1795_6;

wire[31:0] addr_1795_6;

Selector_2 s1795_6(wires_448_5[3], addr_448_5, wires_1795_6,addr_1795_6);

wire[3:0] wires_1796_6;

wire[31:0] addr_1796_6;

Selector_2 s1796_6(wires_449_5[0], addr_449_5, wires_1796_6,addr_1796_6);

wire[3:0] wires_1797_6;

wire[31:0] addr_1797_6;

Selector_2 s1797_6(wires_449_5[1], addr_449_5, wires_1797_6,addr_1797_6);

wire[3:0] wires_1798_6;

wire[31:0] addr_1798_6;

Selector_2 s1798_6(wires_449_5[2], addr_449_5, wires_1798_6,addr_1798_6);

wire[3:0] wires_1799_6;

wire[31:0] addr_1799_6;

Selector_2 s1799_6(wires_449_5[3], addr_449_5, wires_1799_6,addr_1799_6);

wire[3:0] wires_1800_6;

wire[31:0] addr_1800_6;

Selector_2 s1800_6(wires_450_5[0], addr_450_5, wires_1800_6,addr_1800_6);

wire[3:0] wires_1801_6;

wire[31:0] addr_1801_6;

Selector_2 s1801_6(wires_450_5[1], addr_450_5, wires_1801_6,addr_1801_6);

wire[3:0] wires_1802_6;

wire[31:0] addr_1802_6;

Selector_2 s1802_6(wires_450_5[2], addr_450_5, wires_1802_6,addr_1802_6);

wire[3:0] wires_1803_6;

wire[31:0] addr_1803_6;

Selector_2 s1803_6(wires_450_5[3], addr_450_5, wires_1803_6,addr_1803_6);

wire[3:0] wires_1804_6;

wire[31:0] addr_1804_6;

Selector_2 s1804_6(wires_451_5[0], addr_451_5, wires_1804_6,addr_1804_6);

wire[3:0] wires_1805_6;

wire[31:0] addr_1805_6;

Selector_2 s1805_6(wires_451_5[1], addr_451_5, wires_1805_6,addr_1805_6);

wire[3:0] wires_1806_6;

wire[31:0] addr_1806_6;

Selector_2 s1806_6(wires_451_5[2], addr_451_5, wires_1806_6,addr_1806_6);

wire[3:0] wires_1807_6;

wire[31:0] addr_1807_6;

Selector_2 s1807_6(wires_451_5[3], addr_451_5, wires_1807_6,addr_1807_6);

wire[3:0] wires_1808_6;

wire[31:0] addr_1808_6;

Selector_2 s1808_6(wires_452_5[0], addr_452_5, wires_1808_6,addr_1808_6);

wire[3:0] wires_1809_6;

wire[31:0] addr_1809_6;

Selector_2 s1809_6(wires_452_5[1], addr_452_5, wires_1809_6,addr_1809_6);

wire[3:0] wires_1810_6;

wire[31:0] addr_1810_6;

Selector_2 s1810_6(wires_452_5[2], addr_452_5, wires_1810_6,addr_1810_6);

wire[3:0] wires_1811_6;

wire[31:0] addr_1811_6;

Selector_2 s1811_6(wires_452_5[3], addr_452_5, wires_1811_6,addr_1811_6);

wire[3:0] wires_1812_6;

wire[31:0] addr_1812_6;

Selector_2 s1812_6(wires_453_5[0], addr_453_5, wires_1812_6,addr_1812_6);

wire[3:0] wires_1813_6;

wire[31:0] addr_1813_6;

Selector_2 s1813_6(wires_453_5[1], addr_453_5, wires_1813_6,addr_1813_6);

wire[3:0] wires_1814_6;

wire[31:0] addr_1814_6;

Selector_2 s1814_6(wires_453_5[2], addr_453_5, wires_1814_6,addr_1814_6);

wire[3:0] wires_1815_6;

wire[31:0] addr_1815_6;

Selector_2 s1815_6(wires_453_5[3], addr_453_5, wires_1815_6,addr_1815_6);

wire[3:0] wires_1816_6;

wire[31:0] addr_1816_6;

Selector_2 s1816_6(wires_454_5[0], addr_454_5, wires_1816_6,addr_1816_6);

wire[3:0] wires_1817_6;

wire[31:0] addr_1817_6;

Selector_2 s1817_6(wires_454_5[1], addr_454_5, wires_1817_6,addr_1817_6);

wire[3:0] wires_1818_6;

wire[31:0] addr_1818_6;

Selector_2 s1818_6(wires_454_5[2], addr_454_5, wires_1818_6,addr_1818_6);

wire[3:0] wires_1819_6;

wire[31:0] addr_1819_6;

Selector_2 s1819_6(wires_454_5[3], addr_454_5, wires_1819_6,addr_1819_6);

wire[3:0] wires_1820_6;

wire[31:0] addr_1820_6;

Selector_2 s1820_6(wires_455_5[0], addr_455_5, wires_1820_6,addr_1820_6);

wire[3:0] wires_1821_6;

wire[31:0] addr_1821_6;

Selector_2 s1821_6(wires_455_5[1], addr_455_5, wires_1821_6,addr_1821_6);

wire[3:0] wires_1822_6;

wire[31:0] addr_1822_6;

Selector_2 s1822_6(wires_455_5[2], addr_455_5, wires_1822_6,addr_1822_6);

wire[3:0] wires_1823_6;

wire[31:0] addr_1823_6;

Selector_2 s1823_6(wires_455_5[3], addr_455_5, wires_1823_6,addr_1823_6);

wire[3:0] wires_1824_6;

wire[31:0] addr_1824_6;

Selector_2 s1824_6(wires_456_5[0], addr_456_5, wires_1824_6,addr_1824_6);

wire[3:0] wires_1825_6;

wire[31:0] addr_1825_6;

Selector_2 s1825_6(wires_456_5[1], addr_456_5, wires_1825_6,addr_1825_6);

wire[3:0] wires_1826_6;

wire[31:0] addr_1826_6;

Selector_2 s1826_6(wires_456_5[2], addr_456_5, wires_1826_6,addr_1826_6);

wire[3:0] wires_1827_6;

wire[31:0] addr_1827_6;

Selector_2 s1827_6(wires_456_5[3], addr_456_5, wires_1827_6,addr_1827_6);

wire[3:0] wires_1828_6;

wire[31:0] addr_1828_6;

Selector_2 s1828_6(wires_457_5[0], addr_457_5, wires_1828_6,addr_1828_6);

wire[3:0] wires_1829_6;

wire[31:0] addr_1829_6;

Selector_2 s1829_6(wires_457_5[1], addr_457_5, wires_1829_6,addr_1829_6);

wire[3:0] wires_1830_6;

wire[31:0] addr_1830_6;

Selector_2 s1830_6(wires_457_5[2], addr_457_5, wires_1830_6,addr_1830_6);

wire[3:0] wires_1831_6;

wire[31:0] addr_1831_6;

Selector_2 s1831_6(wires_457_5[3], addr_457_5, wires_1831_6,addr_1831_6);

wire[3:0] wires_1832_6;

wire[31:0] addr_1832_6;

Selector_2 s1832_6(wires_458_5[0], addr_458_5, wires_1832_6,addr_1832_6);

wire[3:0] wires_1833_6;

wire[31:0] addr_1833_6;

Selector_2 s1833_6(wires_458_5[1], addr_458_5, wires_1833_6,addr_1833_6);

wire[3:0] wires_1834_6;

wire[31:0] addr_1834_6;

Selector_2 s1834_6(wires_458_5[2], addr_458_5, wires_1834_6,addr_1834_6);

wire[3:0] wires_1835_6;

wire[31:0] addr_1835_6;

Selector_2 s1835_6(wires_458_5[3], addr_458_5, wires_1835_6,addr_1835_6);

wire[3:0] wires_1836_6;

wire[31:0] addr_1836_6;

Selector_2 s1836_6(wires_459_5[0], addr_459_5, wires_1836_6,addr_1836_6);

wire[3:0] wires_1837_6;

wire[31:0] addr_1837_6;

Selector_2 s1837_6(wires_459_5[1], addr_459_5, wires_1837_6,addr_1837_6);

wire[3:0] wires_1838_6;

wire[31:0] addr_1838_6;

Selector_2 s1838_6(wires_459_5[2], addr_459_5, wires_1838_6,addr_1838_6);

wire[3:0] wires_1839_6;

wire[31:0] addr_1839_6;

Selector_2 s1839_6(wires_459_5[3], addr_459_5, wires_1839_6,addr_1839_6);

wire[3:0] wires_1840_6;

wire[31:0] addr_1840_6;

Selector_2 s1840_6(wires_460_5[0], addr_460_5, wires_1840_6,addr_1840_6);

wire[3:0] wires_1841_6;

wire[31:0] addr_1841_6;

Selector_2 s1841_6(wires_460_5[1], addr_460_5, wires_1841_6,addr_1841_6);

wire[3:0] wires_1842_6;

wire[31:0] addr_1842_6;

Selector_2 s1842_6(wires_460_5[2], addr_460_5, wires_1842_6,addr_1842_6);

wire[3:0] wires_1843_6;

wire[31:0] addr_1843_6;

Selector_2 s1843_6(wires_460_5[3], addr_460_5, wires_1843_6,addr_1843_6);

wire[3:0] wires_1844_6;

wire[31:0] addr_1844_6;

Selector_2 s1844_6(wires_461_5[0], addr_461_5, wires_1844_6,addr_1844_6);

wire[3:0] wires_1845_6;

wire[31:0] addr_1845_6;

Selector_2 s1845_6(wires_461_5[1], addr_461_5, wires_1845_6,addr_1845_6);

wire[3:0] wires_1846_6;

wire[31:0] addr_1846_6;

Selector_2 s1846_6(wires_461_5[2], addr_461_5, wires_1846_6,addr_1846_6);

wire[3:0] wires_1847_6;

wire[31:0] addr_1847_6;

Selector_2 s1847_6(wires_461_5[3], addr_461_5, wires_1847_6,addr_1847_6);

wire[3:0] wires_1848_6;

wire[31:0] addr_1848_6;

Selector_2 s1848_6(wires_462_5[0], addr_462_5, wires_1848_6,addr_1848_6);

wire[3:0] wires_1849_6;

wire[31:0] addr_1849_6;

Selector_2 s1849_6(wires_462_5[1], addr_462_5, wires_1849_6,addr_1849_6);

wire[3:0] wires_1850_6;

wire[31:0] addr_1850_6;

Selector_2 s1850_6(wires_462_5[2], addr_462_5, wires_1850_6,addr_1850_6);

wire[3:0] wires_1851_6;

wire[31:0] addr_1851_6;

Selector_2 s1851_6(wires_462_5[3], addr_462_5, wires_1851_6,addr_1851_6);

wire[3:0] wires_1852_6;

wire[31:0] addr_1852_6;

Selector_2 s1852_6(wires_463_5[0], addr_463_5, wires_1852_6,addr_1852_6);

wire[3:0] wires_1853_6;

wire[31:0] addr_1853_6;

Selector_2 s1853_6(wires_463_5[1], addr_463_5, wires_1853_6,addr_1853_6);

wire[3:0] wires_1854_6;

wire[31:0] addr_1854_6;

Selector_2 s1854_6(wires_463_5[2], addr_463_5, wires_1854_6,addr_1854_6);

wire[3:0] wires_1855_6;

wire[31:0] addr_1855_6;

Selector_2 s1855_6(wires_463_5[3], addr_463_5, wires_1855_6,addr_1855_6);

wire[3:0] wires_1856_6;

wire[31:0] addr_1856_6;

Selector_2 s1856_6(wires_464_5[0], addr_464_5, wires_1856_6,addr_1856_6);

wire[3:0] wires_1857_6;

wire[31:0] addr_1857_6;

Selector_2 s1857_6(wires_464_5[1], addr_464_5, wires_1857_6,addr_1857_6);

wire[3:0] wires_1858_6;

wire[31:0] addr_1858_6;

Selector_2 s1858_6(wires_464_5[2], addr_464_5, wires_1858_6,addr_1858_6);

wire[3:0] wires_1859_6;

wire[31:0] addr_1859_6;

Selector_2 s1859_6(wires_464_5[3], addr_464_5, wires_1859_6,addr_1859_6);

wire[3:0] wires_1860_6;

wire[31:0] addr_1860_6;

Selector_2 s1860_6(wires_465_5[0], addr_465_5, wires_1860_6,addr_1860_6);

wire[3:0] wires_1861_6;

wire[31:0] addr_1861_6;

Selector_2 s1861_6(wires_465_5[1], addr_465_5, wires_1861_6,addr_1861_6);

wire[3:0] wires_1862_6;

wire[31:0] addr_1862_6;

Selector_2 s1862_6(wires_465_5[2], addr_465_5, wires_1862_6,addr_1862_6);

wire[3:0] wires_1863_6;

wire[31:0] addr_1863_6;

Selector_2 s1863_6(wires_465_5[3], addr_465_5, wires_1863_6,addr_1863_6);

wire[3:0] wires_1864_6;

wire[31:0] addr_1864_6;

Selector_2 s1864_6(wires_466_5[0], addr_466_5, wires_1864_6,addr_1864_6);

wire[3:0] wires_1865_6;

wire[31:0] addr_1865_6;

Selector_2 s1865_6(wires_466_5[1], addr_466_5, wires_1865_6,addr_1865_6);

wire[3:0] wires_1866_6;

wire[31:0] addr_1866_6;

Selector_2 s1866_6(wires_466_5[2], addr_466_5, wires_1866_6,addr_1866_6);

wire[3:0] wires_1867_6;

wire[31:0] addr_1867_6;

Selector_2 s1867_6(wires_466_5[3], addr_466_5, wires_1867_6,addr_1867_6);

wire[3:0] wires_1868_6;

wire[31:0] addr_1868_6;

Selector_2 s1868_6(wires_467_5[0], addr_467_5, wires_1868_6,addr_1868_6);

wire[3:0] wires_1869_6;

wire[31:0] addr_1869_6;

Selector_2 s1869_6(wires_467_5[1], addr_467_5, wires_1869_6,addr_1869_6);

wire[3:0] wires_1870_6;

wire[31:0] addr_1870_6;

Selector_2 s1870_6(wires_467_5[2], addr_467_5, wires_1870_6,addr_1870_6);

wire[3:0] wires_1871_6;

wire[31:0] addr_1871_6;

Selector_2 s1871_6(wires_467_5[3], addr_467_5, wires_1871_6,addr_1871_6);

wire[3:0] wires_1872_6;

wire[31:0] addr_1872_6;

Selector_2 s1872_6(wires_468_5[0], addr_468_5, wires_1872_6,addr_1872_6);

wire[3:0] wires_1873_6;

wire[31:0] addr_1873_6;

Selector_2 s1873_6(wires_468_5[1], addr_468_5, wires_1873_6,addr_1873_6);

wire[3:0] wires_1874_6;

wire[31:0] addr_1874_6;

Selector_2 s1874_6(wires_468_5[2], addr_468_5, wires_1874_6,addr_1874_6);

wire[3:0] wires_1875_6;

wire[31:0] addr_1875_6;

Selector_2 s1875_6(wires_468_5[3], addr_468_5, wires_1875_6,addr_1875_6);

wire[3:0] wires_1876_6;

wire[31:0] addr_1876_6;

Selector_2 s1876_6(wires_469_5[0], addr_469_5, wires_1876_6,addr_1876_6);

wire[3:0] wires_1877_6;

wire[31:0] addr_1877_6;

Selector_2 s1877_6(wires_469_5[1], addr_469_5, wires_1877_6,addr_1877_6);

wire[3:0] wires_1878_6;

wire[31:0] addr_1878_6;

Selector_2 s1878_6(wires_469_5[2], addr_469_5, wires_1878_6,addr_1878_6);

wire[3:0] wires_1879_6;

wire[31:0] addr_1879_6;

Selector_2 s1879_6(wires_469_5[3], addr_469_5, wires_1879_6,addr_1879_6);

wire[3:0] wires_1880_6;

wire[31:0] addr_1880_6;

Selector_2 s1880_6(wires_470_5[0], addr_470_5, wires_1880_6,addr_1880_6);

wire[3:0] wires_1881_6;

wire[31:0] addr_1881_6;

Selector_2 s1881_6(wires_470_5[1], addr_470_5, wires_1881_6,addr_1881_6);

wire[3:0] wires_1882_6;

wire[31:0] addr_1882_6;

Selector_2 s1882_6(wires_470_5[2], addr_470_5, wires_1882_6,addr_1882_6);

wire[3:0] wires_1883_6;

wire[31:0] addr_1883_6;

Selector_2 s1883_6(wires_470_5[3], addr_470_5, wires_1883_6,addr_1883_6);

wire[3:0] wires_1884_6;

wire[31:0] addr_1884_6;

Selector_2 s1884_6(wires_471_5[0], addr_471_5, wires_1884_6,addr_1884_6);

wire[3:0] wires_1885_6;

wire[31:0] addr_1885_6;

Selector_2 s1885_6(wires_471_5[1], addr_471_5, wires_1885_6,addr_1885_6);

wire[3:0] wires_1886_6;

wire[31:0] addr_1886_6;

Selector_2 s1886_6(wires_471_5[2], addr_471_5, wires_1886_6,addr_1886_6);

wire[3:0] wires_1887_6;

wire[31:0] addr_1887_6;

Selector_2 s1887_6(wires_471_5[3], addr_471_5, wires_1887_6,addr_1887_6);

wire[3:0] wires_1888_6;

wire[31:0] addr_1888_6;

Selector_2 s1888_6(wires_472_5[0], addr_472_5, wires_1888_6,addr_1888_6);

wire[3:0] wires_1889_6;

wire[31:0] addr_1889_6;

Selector_2 s1889_6(wires_472_5[1], addr_472_5, wires_1889_6,addr_1889_6);

wire[3:0] wires_1890_6;

wire[31:0] addr_1890_6;

Selector_2 s1890_6(wires_472_5[2], addr_472_5, wires_1890_6,addr_1890_6);

wire[3:0] wires_1891_6;

wire[31:0] addr_1891_6;

Selector_2 s1891_6(wires_472_5[3], addr_472_5, wires_1891_6,addr_1891_6);

wire[3:0] wires_1892_6;

wire[31:0] addr_1892_6;

Selector_2 s1892_6(wires_473_5[0], addr_473_5, wires_1892_6,addr_1892_6);

wire[3:0] wires_1893_6;

wire[31:0] addr_1893_6;

Selector_2 s1893_6(wires_473_5[1], addr_473_5, wires_1893_6,addr_1893_6);

wire[3:0] wires_1894_6;

wire[31:0] addr_1894_6;

Selector_2 s1894_6(wires_473_5[2], addr_473_5, wires_1894_6,addr_1894_6);

wire[3:0] wires_1895_6;

wire[31:0] addr_1895_6;

Selector_2 s1895_6(wires_473_5[3], addr_473_5, wires_1895_6,addr_1895_6);

wire[3:0] wires_1896_6;

wire[31:0] addr_1896_6;

Selector_2 s1896_6(wires_474_5[0], addr_474_5, wires_1896_6,addr_1896_6);

wire[3:0] wires_1897_6;

wire[31:0] addr_1897_6;

Selector_2 s1897_6(wires_474_5[1], addr_474_5, wires_1897_6,addr_1897_6);

wire[3:0] wires_1898_6;

wire[31:0] addr_1898_6;

Selector_2 s1898_6(wires_474_5[2], addr_474_5, wires_1898_6,addr_1898_6);

wire[3:0] wires_1899_6;

wire[31:0] addr_1899_6;

Selector_2 s1899_6(wires_474_5[3], addr_474_5, wires_1899_6,addr_1899_6);

wire[3:0] wires_1900_6;

wire[31:0] addr_1900_6;

Selector_2 s1900_6(wires_475_5[0], addr_475_5, wires_1900_6,addr_1900_6);

wire[3:0] wires_1901_6;

wire[31:0] addr_1901_6;

Selector_2 s1901_6(wires_475_5[1], addr_475_5, wires_1901_6,addr_1901_6);

wire[3:0] wires_1902_6;

wire[31:0] addr_1902_6;

Selector_2 s1902_6(wires_475_5[2], addr_475_5, wires_1902_6,addr_1902_6);

wire[3:0] wires_1903_6;

wire[31:0] addr_1903_6;

Selector_2 s1903_6(wires_475_5[3], addr_475_5, wires_1903_6,addr_1903_6);

wire[3:0] wires_1904_6;

wire[31:0] addr_1904_6;

Selector_2 s1904_6(wires_476_5[0], addr_476_5, wires_1904_6,addr_1904_6);

wire[3:0] wires_1905_6;

wire[31:0] addr_1905_6;

Selector_2 s1905_6(wires_476_5[1], addr_476_5, wires_1905_6,addr_1905_6);

wire[3:0] wires_1906_6;

wire[31:0] addr_1906_6;

Selector_2 s1906_6(wires_476_5[2], addr_476_5, wires_1906_6,addr_1906_6);

wire[3:0] wires_1907_6;

wire[31:0] addr_1907_6;

Selector_2 s1907_6(wires_476_5[3], addr_476_5, wires_1907_6,addr_1907_6);

wire[3:0] wires_1908_6;

wire[31:0] addr_1908_6;

Selector_2 s1908_6(wires_477_5[0], addr_477_5, wires_1908_6,addr_1908_6);

wire[3:0] wires_1909_6;

wire[31:0] addr_1909_6;

Selector_2 s1909_6(wires_477_5[1], addr_477_5, wires_1909_6,addr_1909_6);

wire[3:0] wires_1910_6;

wire[31:0] addr_1910_6;

Selector_2 s1910_6(wires_477_5[2], addr_477_5, wires_1910_6,addr_1910_6);

wire[3:0] wires_1911_6;

wire[31:0] addr_1911_6;

Selector_2 s1911_6(wires_477_5[3], addr_477_5, wires_1911_6,addr_1911_6);

wire[3:0] wires_1912_6;

wire[31:0] addr_1912_6;

Selector_2 s1912_6(wires_478_5[0], addr_478_5, wires_1912_6,addr_1912_6);

wire[3:0] wires_1913_6;

wire[31:0] addr_1913_6;

Selector_2 s1913_6(wires_478_5[1], addr_478_5, wires_1913_6,addr_1913_6);

wire[3:0] wires_1914_6;

wire[31:0] addr_1914_6;

Selector_2 s1914_6(wires_478_5[2], addr_478_5, wires_1914_6,addr_1914_6);

wire[3:0] wires_1915_6;

wire[31:0] addr_1915_6;

Selector_2 s1915_6(wires_478_5[3], addr_478_5, wires_1915_6,addr_1915_6);

wire[3:0] wires_1916_6;

wire[31:0] addr_1916_6;

Selector_2 s1916_6(wires_479_5[0], addr_479_5, wires_1916_6,addr_1916_6);

wire[3:0] wires_1917_6;

wire[31:0] addr_1917_6;

Selector_2 s1917_6(wires_479_5[1], addr_479_5, wires_1917_6,addr_1917_6);

wire[3:0] wires_1918_6;

wire[31:0] addr_1918_6;

Selector_2 s1918_6(wires_479_5[2], addr_479_5, wires_1918_6,addr_1918_6);

wire[3:0] wires_1919_6;

wire[31:0] addr_1919_6;

Selector_2 s1919_6(wires_479_5[3], addr_479_5, wires_1919_6,addr_1919_6);

wire[3:0] wires_1920_6;

wire[31:0] addr_1920_6;

Selector_2 s1920_6(wires_480_5[0], addr_480_5, wires_1920_6,addr_1920_6);

wire[3:0] wires_1921_6;

wire[31:0] addr_1921_6;

Selector_2 s1921_6(wires_480_5[1], addr_480_5, wires_1921_6,addr_1921_6);

wire[3:0] wires_1922_6;

wire[31:0] addr_1922_6;

Selector_2 s1922_6(wires_480_5[2], addr_480_5, wires_1922_6,addr_1922_6);

wire[3:0] wires_1923_6;

wire[31:0] addr_1923_6;

Selector_2 s1923_6(wires_480_5[3], addr_480_5, wires_1923_6,addr_1923_6);

wire[3:0] wires_1924_6;

wire[31:0] addr_1924_6;

Selector_2 s1924_6(wires_481_5[0], addr_481_5, wires_1924_6,addr_1924_6);

wire[3:0] wires_1925_6;

wire[31:0] addr_1925_6;

Selector_2 s1925_6(wires_481_5[1], addr_481_5, wires_1925_6,addr_1925_6);

wire[3:0] wires_1926_6;

wire[31:0] addr_1926_6;

Selector_2 s1926_6(wires_481_5[2], addr_481_5, wires_1926_6,addr_1926_6);

wire[3:0] wires_1927_6;

wire[31:0] addr_1927_6;

Selector_2 s1927_6(wires_481_5[3], addr_481_5, wires_1927_6,addr_1927_6);

wire[3:0] wires_1928_6;

wire[31:0] addr_1928_6;

Selector_2 s1928_6(wires_482_5[0], addr_482_5, wires_1928_6,addr_1928_6);

wire[3:0] wires_1929_6;

wire[31:0] addr_1929_6;

Selector_2 s1929_6(wires_482_5[1], addr_482_5, wires_1929_6,addr_1929_6);

wire[3:0] wires_1930_6;

wire[31:0] addr_1930_6;

Selector_2 s1930_6(wires_482_5[2], addr_482_5, wires_1930_6,addr_1930_6);

wire[3:0] wires_1931_6;

wire[31:0] addr_1931_6;

Selector_2 s1931_6(wires_482_5[3], addr_482_5, wires_1931_6,addr_1931_6);

wire[3:0] wires_1932_6;

wire[31:0] addr_1932_6;

Selector_2 s1932_6(wires_483_5[0], addr_483_5, wires_1932_6,addr_1932_6);

wire[3:0] wires_1933_6;

wire[31:0] addr_1933_6;

Selector_2 s1933_6(wires_483_5[1], addr_483_5, wires_1933_6,addr_1933_6);

wire[3:0] wires_1934_6;

wire[31:0] addr_1934_6;

Selector_2 s1934_6(wires_483_5[2], addr_483_5, wires_1934_6,addr_1934_6);

wire[3:0] wires_1935_6;

wire[31:0] addr_1935_6;

Selector_2 s1935_6(wires_483_5[3], addr_483_5, wires_1935_6,addr_1935_6);

wire[3:0] wires_1936_6;

wire[31:0] addr_1936_6;

Selector_2 s1936_6(wires_484_5[0], addr_484_5, wires_1936_6,addr_1936_6);

wire[3:0] wires_1937_6;

wire[31:0] addr_1937_6;

Selector_2 s1937_6(wires_484_5[1], addr_484_5, wires_1937_6,addr_1937_6);

wire[3:0] wires_1938_6;

wire[31:0] addr_1938_6;

Selector_2 s1938_6(wires_484_5[2], addr_484_5, wires_1938_6,addr_1938_6);

wire[3:0] wires_1939_6;

wire[31:0] addr_1939_6;

Selector_2 s1939_6(wires_484_5[3], addr_484_5, wires_1939_6,addr_1939_6);

wire[3:0] wires_1940_6;

wire[31:0] addr_1940_6;

Selector_2 s1940_6(wires_485_5[0], addr_485_5, wires_1940_6,addr_1940_6);

wire[3:0] wires_1941_6;

wire[31:0] addr_1941_6;

Selector_2 s1941_6(wires_485_5[1], addr_485_5, wires_1941_6,addr_1941_6);

wire[3:0] wires_1942_6;

wire[31:0] addr_1942_6;

Selector_2 s1942_6(wires_485_5[2], addr_485_5, wires_1942_6,addr_1942_6);

wire[3:0] wires_1943_6;

wire[31:0] addr_1943_6;

Selector_2 s1943_6(wires_485_5[3], addr_485_5, wires_1943_6,addr_1943_6);

wire[3:0] wires_1944_6;

wire[31:0] addr_1944_6;

Selector_2 s1944_6(wires_486_5[0], addr_486_5, wires_1944_6,addr_1944_6);

wire[3:0] wires_1945_6;

wire[31:0] addr_1945_6;

Selector_2 s1945_6(wires_486_5[1], addr_486_5, wires_1945_6,addr_1945_6);

wire[3:0] wires_1946_6;

wire[31:0] addr_1946_6;

Selector_2 s1946_6(wires_486_5[2], addr_486_5, wires_1946_6,addr_1946_6);

wire[3:0] wires_1947_6;

wire[31:0] addr_1947_6;

Selector_2 s1947_6(wires_486_5[3], addr_486_5, wires_1947_6,addr_1947_6);

wire[3:0] wires_1948_6;

wire[31:0] addr_1948_6;

Selector_2 s1948_6(wires_487_5[0], addr_487_5, wires_1948_6,addr_1948_6);

wire[3:0] wires_1949_6;

wire[31:0] addr_1949_6;

Selector_2 s1949_6(wires_487_5[1], addr_487_5, wires_1949_6,addr_1949_6);

wire[3:0] wires_1950_6;

wire[31:0] addr_1950_6;

Selector_2 s1950_6(wires_487_5[2], addr_487_5, wires_1950_6,addr_1950_6);

wire[3:0] wires_1951_6;

wire[31:0] addr_1951_6;

Selector_2 s1951_6(wires_487_5[3], addr_487_5, wires_1951_6,addr_1951_6);

wire[3:0] wires_1952_6;

wire[31:0] addr_1952_6;

Selector_2 s1952_6(wires_488_5[0], addr_488_5, wires_1952_6,addr_1952_6);

wire[3:0] wires_1953_6;

wire[31:0] addr_1953_6;

Selector_2 s1953_6(wires_488_5[1], addr_488_5, wires_1953_6,addr_1953_6);

wire[3:0] wires_1954_6;

wire[31:0] addr_1954_6;

Selector_2 s1954_6(wires_488_5[2], addr_488_5, wires_1954_6,addr_1954_6);

wire[3:0] wires_1955_6;

wire[31:0] addr_1955_6;

Selector_2 s1955_6(wires_488_5[3], addr_488_5, wires_1955_6,addr_1955_6);

wire[3:0] wires_1956_6;

wire[31:0] addr_1956_6;

Selector_2 s1956_6(wires_489_5[0], addr_489_5, wires_1956_6,addr_1956_6);

wire[3:0] wires_1957_6;

wire[31:0] addr_1957_6;

Selector_2 s1957_6(wires_489_5[1], addr_489_5, wires_1957_6,addr_1957_6);

wire[3:0] wires_1958_6;

wire[31:0] addr_1958_6;

Selector_2 s1958_6(wires_489_5[2], addr_489_5, wires_1958_6,addr_1958_6);

wire[3:0] wires_1959_6;

wire[31:0] addr_1959_6;

Selector_2 s1959_6(wires_489_5[3], addr_489_5, wires_1959_6,addr_1959_6);

wire[3:0] wires_1960_6;

wire[31:0] addr_1960_6;

Selector_2 s1960_6(wires_490_5[0], addr_490_5, wires_1960_6,addr_1960_6);

wire[3:0] wires_1961_6;

wire[31:0] addr_1961_6;

Selector_2 s1961_6(wires_490_5[1], addr_490_5, wires_1961_6,addr_1961_6);

wire[3:0] wires_1962_6;

wire[31:0] addr_1962_6;

Selector_2 s1962_6(wires_490_5[2], addr_490_5, wires_1962_6,addr_1962_6);

wire[3:0] wires_1963_6;

wire[31:0] addr_1963_6;

Selector_2 s1963_6(wires_490_5[3], addr_490_5, wires_1963_6,addr_1963_6);

wire[3:0] wires_1964_6;

wire[31:0] addr_1964_6;

Selector_2 s1964_6(wires_491_5[0], addr_491_5, wires_1964_6,addr_1964_6);

wire[3:0] wires_1965_6;

wire[31:0] addr_1965_6;

Selector_2 s1965_6(wires_491_5[1], addr_491_5, wires_1965_6,addr_1965_6);

wire[3:0] wires_1966_6;

wire[31:0] addr_1966_6;

Selector_2 s1966_6(wires_491_5[2], addr_491_5, wires_1966_6,addr_1966_6);

wire[3:0] wires_1967_6;

wire[31:0] addr_1967_6;

Selector_2 s1967_6(wires_491_5[3], addr_491_5, wires_1967_6,addr_1967_6);

wire[3:0] wires_1968_6;

wire[31:0] addr_1968_6;

Selector_2 s1968_6(wires_492_5[0], addr_492_5, wires_1968_6,addr_1968_6);

wire[3:0] wires_1969_6;

wire[31:0] addr_1969_6;

Selector_2 s1969_6(wires_492_5[1], addr_492_5, wires_1969_6,addr_1969_6);

wire[3:0] wires_1970_6;

wire[31:0] addr_1970_6;

Selector_2 s1970_6(wires_492_5[2], addr_492_5, wires_1970_6,addr_1970_6);

wire[3:0] wires_1971_6;

wire[31:0] addr_1971_6;

Selector_2 s1971_6(wires_492_5[3], addr_492_5, wires_1971_6,addr_1971_6);

wire[3:0] wires_1972_6;

wire[31:0] addr_1972_6;

Selector_2 s1972_6(wires_493_5[0], addr_493_5, wires_1972_6,addr_1972_6);

wire[3:0] wires_1973_6;

wire[31:0] addr_1973_6;

Selector_2 s1973_6(wires_493_5[1], addr_493_5, wires_1973_6,addr_1973_6);

wire[3:0] wires_1974_6;

wire[31:0] addr_1974_6;

Selector_2 s1974_6(wires_493_5[2], addr_493_5, wires_1974_6,addr_1974_6);

wire[3:0] wires_1975_6;

wire[31:0] addr_1975_6;

Selector_2 s1975_6(wires_493_5[3], addr_493_5, wires_1975_6,addr_1975_6);

wire[3:0] wires_1976_6;

wire[31:0] addr_1976_6;

Selector_2 s1976_6(wires_494_5[0], addr_494_5, wires_1976_6,addr_1976_6);

wire[3:0] wires_1977_6;

wire[31:0] addr_1977_6;

Selector_2 s1977_6(wires_494_5[1], addr_494_5, wires_1977_6,addr_1977_6);

wire[3:0] wires_1978_6;

wire[31:0] addr_1978_6;

Selector_2 s1978_6(wires_494_5[2], addr_494_5, wires_1978_6,addr_1978_6);

wire[3:0] wires_1979_6;

wire[31:0] addr_1979_6;

Selector_2 s1979_6(wires_494_5[3], addr_494_5, wires_1979_6,addr_1979_6);

wire[3:0] wires_1980_6;

wire[31:0] addr_1980_6;

Selector_2 s1980_6(wires_495_5[0], addr_495_5, wires_1980_6,addr_1980_6);

wire[3:0] wires_1981_6;

wire[31:0] addr_1981_6;

Selector_2 s1981_6(wires_495_5[1], addr_495_5, wires_1981_6,addr_1981_6);

wire[3:0] wires_1982_6;

wire[31:0] addr_1982_6;

Selector_2 s1982_6(wires_495_5[2], addr_495_5, wires_1982_6,addr_1982_6);

wire[3:0] wires_1983_6;

wire[31:0] addr_1983_6;

Selector_2 s1983_6(wires_495_5[3], addr_495_5, wires_1983_6,addr_1983_6);

wire[3:0] wires_1984_6;

wire[31:0] addr_1984_6;

Selector_2 s1984_6(wires_496_5[0], addr_496_5, wires_1984_6,addr_1984_6);

wire[3:0] wires_1985_6;

wire[31:0] addr_1985_6;

Selector_2 s1985_6(wires_496_5[1], addr_496_5, wires_1985_6,addr_1985_6);

wire[3:0] wires_1986_6;

wire[31:0] addr_1986_6;

Selector_2 s1986_6(wires_496_5[2], addr_496_5, wires_1986_6,addr_1986_6);

wire[3:0] wires_1987_6;

wire[31:0] addr_1987_6;

Selector_2 s1987_6(wires_496_5[3], addr_496_5, wires_1987_6,addr_1987_6);

wire[3:0] wires_1988_6;

wire[31:0] addr_1988_6;

Selector_2 s1988_6(wires_497_5[0], addr_497_5, wires_1988_6,addr_1988_6);

wire[3:0] wires_1989_6;

wire[31:0] addr_1989_6;

Selector_2 s1989_6(wires_497_5[1], addr_497_5, wires_1989_6,addr_1989_6);

wire[3:0] wires_1990_6;

wire[31:0] addr_1990_6;

Selector_2 s1990_6(wires_497_5[2], addr_497_5, wires_1990_6,addr_1990_6);

wire[3:0] wires_1991_6;

wire[31:0] addr_1991_6;

Selector_2 s1991_6(wires_497_5[3], addr_497_5, wires_1991_6,addr_1991_6);

wire[3:0] wires_1992_6;

wire[31:0] addr_1992_6;

Selector_2 s1992_6(wires_498_5[0], addr_498_5, wires_1992_6,addr_1992_6);

wire[3:0] wires_1993_6;

wire[31:0] addr_1993_6;

Selector_2 s1993_6(wires_498_5[1], addr_498_5, wires_1993_6,addr_1993_6);

wire[3:0] wires_1994_6;

wire[31:0] addr_1994_6;

Selector_2 s1994_6(wires_498_5[2], addr_498_5, wires_1994_6,addr_1994_6);

wire[3:0] wires_1995_6;

wire[31:0] addr_1995_6;

Selector_2 s1995_6(wires_498_5[3], addr_498_5, wires_1995_6,addr_1995_6);

wire[3:0] wires_1996_6;

wire[31:0] addr_1996_6;

Selector_2 s1996_6(wires_499_5[0], addr_499_5, wires_1996_6,addr_1996_6);

wire[3:0] wires_1997_6;

wire[31:0] addr_1997_6;

Selector_2 s1997_6(wires_499_5[1], addr_499_5, wires_1997_6,addr_1997_6);

wire[3:0] wires_1998_6;

wire[31:0] addr_1998_6;

Selector_2 s1998_6(wires_499_5[2], addr_499_5, wires_1998_6,addr_1998_6);

wire[3:0] wires_1999_6;

wire[31:0] addr_1999_6;

Selector_2 s1999_6(wires_499_5[3], addr_499_5, wires_1999_6,addr_1999_6);

wire[3:0] wires_2000_6;

wire[31:0] addr_2000_6;

Selector_2 s2000_6(wires_500_5[0], addr_500_5, wires_2000_6,addr_2000_6);

wire[3:0] wires_2001_6;

wire[31:0] addr_2001_6;

Selector_2 s2001_6(wires_500_5[1], addr_500_5, wires_2001_6,addr_2001_6);

wire[3:0] wires_2002_6;

wire[31:0] addr_2002_6;

Selector_2 s2002_6(wires_500_5[2], addr_500_5, wires_2002_6,addr_2002_6);

wire[3:0] wires_2003_6;

wire[31:0] addr_2003_6;

Selector_2 s2003_6(wires_500_5[3], addr_500_5, wires_2003_6,addr_2003_6);

wire[3:0] wires_2004_6;

wire[31:0] addr_2004_6;

Selector_2 s2004_6(wires_501_5[0], addr_501_5, wires_2004_6,addr_2004_6);

wire[3:0] wires_2005_6;

wire[31:0] addr_2005_6;

Selector_2 s2005_6(wires_501_5[1], addr_501_5, wires_2005_6,addr_2005_6);

wire[3:0] wires_2006_6;

wire[31:0] addr_2006_6;

Selector_2 s2006_6(wires_501_5[2], addr_501_5, wires_2006_6,addr_2006_6);

wire[3:0] wires_2007_6;

wire[31:0] addr_2007_6;

Selector_2 s2007_6(wires_501_5[3], addr_501_5, wires_2007_6,addr_2007_6);

wire[3:0] wires_2008_6;

wire[31:0] addr_2008_6;

Selector_2 s2008_6(wires_502_5[0], addr_502_5, wires_2008_6,addr_2008_6);

wire[3:0] wires_2009_6;

wire[31:0] addr_2009_6;

Selector_2 s2009_6(wires_502_5[1], addr_502_5, wires_2009_6,addr_2009_6);

wire[3:0] wires_2010_6;

wire[31:0] addr_2010_6;

Selector_2 s2010_6(wires_502_5[2], addr_502_5, wires_2010_6,addr_2010_6);

wire[3:0] wires_2011_6;

wire[31:0] addr_2011_6;

Selector_2 s2011_6(wires_502_5[3], addr_502_5, wires_2011_6,addr_2011_6);

wire[3:0] wires_2012_6;

wire[31:0] addr_2012_6;

Selector_2 s2012_6(wires_503_5[0], addr_503_5, wires_2012_6,addr_2012_6);

wire[3:0] wires_2013_6;

wire[31:0] addr_2013_6;

Selector_2 s2013_6(wires_503_5[1], addr_503_5, wires_2013_6,addr_2013_6);

wire[3:0] wires_2014_6;

wire[31:0] addr_2014_6;

Selector_2 s2014_6(wires_503_5[2], addr_503_5, wires_2014_6,addr_2014_6);

wire[3:0] wires_2015_6;

wire[31:0] addr_2015_6;

Selector_2 s2015_6(wires_503_5[3], addr_503_5, wires_2015_6,addr_2015_6);

wire[3:0] wires_2016_6;

wire[31:0] addr_2016_6;

Selector_2 s2016_6(wires_504_5[0], addr_504_5, wires_2016_6,addr_2016_6);

wire[3:0] wires_2017_6;

wire[31:0] addr_2017_6;

Selector_2 s2017_6(wires_504_5[1], addr_504_5, wires_2017_6,addr_2017_6);

wire[3:0] wires_2018_6;

wire[31:0] addr_2018_6;

Selector_2 s2018_6(wires_504_5[2], addr_504_5, wires_2018_6,addr_2018_6);

wire[3:0] wires_2019_6;

wire[31:0] addr_2019_6;

Selector_2 s2019_6(wires_504_5[3], addr_504_5, wires_2019_6,addr_2019_6);

wire[3:0] wires_2020_6;

wire[31:0] addr_2020_6;

Selector_2 s2020_6(wires_505_5[0], addr_505_5, wires_2020_6,addr_2020_6);

wire[3:0] wires_2021_6;

wire[31:0] addr_2021_6;

Selector_2 s2021_6(wires_505_5[1], addr_505_5, wires_2021_6,addr_2021_6);

wire[3:0] wires_2022_6;

wire[31:0] addr_2022_6;

Selector_2 s2022_6(wires_505_5[2], addr_505_5, wires_2022_6,addr_2022_6);

wire[3:0] wires_2023_6;

wire[31:0] addr_2023_6;

Selector_2 s2023_6(wires_505_5[3], addr_505_5, wires_2023_6,addr_2023_6);

wire[3:0] wires_2024_6;

wire[31:0] addr_2024_6;

Selector_2 s2024_6(wires_506_5[0], addr_506_5, wires_2024_6,addr_2024_6);

wire[3:0] wires_2025_6;

wire[31:0] addr_2025_6;

Selector_2 s2025_6(wires_506_5[1], addr_506_5, wires_2025_6,addr_2025_6);

wire[3:0] wires_2026_6;

wire[31:0] addr_2026_6;

Selector_2 s2026_6(wires_506_5[2], addr_506_5, wires_2026_6,addr_2026_6);

wire[3:0] wires_2027_6;

wire[31:0] addr_2027_6;

Selector_2 s2027_6(wires_506_5[3], addr_506_5, wires_2027_6,addr_2027_6);

wire[3:0] wires_2028_6;

wire[31:0] addr_2028_6;

Selector_2 s2028_6(wires_507_5[0], addr_507_5, wires_2028_6,addr_2028_6);

wire[3:0] wires_2029_6;

wire[31:0] addr_2029_6;

Selector_2 s2029_6(wires_507_5[1], addr_507_5, wires_2029_6,addr_2029_6);

wire[3:0] wires_2030_6;

wire[31:0] addr_2030_6;

Selector_2 s2030_6(wires_507_5[2], addr_507_5, wires_2030_6,addr_2030_6);

wire[3:0] wires_2031_6;

wire[31:0] addr_2031_6;

Selector_2 s2031_6(wires_507_5[3], addr_507_5, wires_2031_6,addr_2031_6);

wire[3:0] wires_2032_6;

wire[31:0] addr_2032_6;

Selector_2 s2032_6(wires_508_5[0], addr_508_5, wires_2032_6,addr_2032_6);

wire[3:0] wires_2033_6;

wire[31:0] addr_2033_6;

Selector_2 s2033_6(wires_508_5[1], addr_508_5, wires_2033_6,addr_2033_6);

wire[3:0] wires_2034_6;

wire[31:0] addr_2034_6;

Selector_2 s2034_6(wires_508_5[2], addr_508_5, wires_2034_6,addr_2034_6);

wire[3:0] wires_2035_6;

wire[31:0] addr_2035_6;

Selector_2 s2035_6(wires_508_5[3], addr_508_5, wires_2035_6,addr_2035_6);

wire[3:0] wires_2036_6;

wire[31:0] addr_2036_6;

Selector_2 s2036_6(wires_509_5[0], addr_509_5, wires_2036_6,addr_2036_6);

wire[3:0] wires_2037_6;

wire[31:0] addr_2037_6;

Selector_2 s2037_6(wires_509_5[1], addr_509_5, wires_2037_6,addr_2037_6);

wire[3:0] wires_2038_6;

wire[31:0] addr_2038_6;

Selector_2 s2038_6(wires_509_5[2], addr_509_5, wires_2038_6,addr_2038_6);

wire[3:0] wires_2039_6;

wire[31:0] addr_2039_6;

Selector_2 s2039_6(wires_509_5[3], addr_509_5, wires_2039_6,addr_2039_6);

wire[3:0] wires_2040_6;

wire[31:0] addr_2040_6;

Selector_2 s2040_6(wires_510_5[0], addr_510_5, wires_2040_6,addr_2040_6);

wire[3:0] wires_2041_6;

wire[31:0] addr_2041_6;

Selector_2 s2041_6(wires_510_5[1], addr_510_5, wires_2041_6,addr_2041_6);

wire[3:0] wires_2042_6;

wire[31:0] addr_2042_6;

Selector_2 s2042_6(wires_510_5[2], addr_510_5, wires_2042_6,addr_2042_6);

wire[3:0] wires_2043_6;

wire[31:0] addr_2043_6;

Selector_2 s2043_6(wires_510_5[3], addr_510_5, wires_2043_6,addr_2043_6);

wire[3:0] wires_2044_6;

wire[31:0] addr_2044_6;

Selector_2 s2044_6(wires_511_5[0], addr_511_5, wires_2044_6,addr_2044_6);

wire[3:0] wires_2045_6;

wire[31:0] addr_2045_6;

Selector_2 s2045_6(wires_511_5[1], addr_511_5, wires_2045_6,addr_2045_6);

wire[3:0] wires_2046_6;

wire[31:0] addr_2046_6;

Selector_2 s2046_6(wires_511_5[2], addr_511_5, wires_2046_6,addr_2046_6);

wire[3:0] wires_2047_6;

wire[31:0] addr_2047_6;

Selector_2 s2047_6(wires_511_5[3], addr_511_5, wires_2047_6,addr_2047_6);

wire[3:0] wires_2048_6;

wire[31:0] addr_2048_6;

Selector_2 s2048_6(wires_512_5[0], addr_512_5, wires_2048_6,addr_2048_6);

wire[3:0] wires_2049_6;

wire[31:0] addr_2049_6;

Selector_2 s2049_6(wires_512_5[1], addr_512_5, wires_2049_6,addr_2049_6);

wire[3:0] wires_2050_6;

wire[31:0] addr_2050_6;

Selector_2 s2050_6(wires_512_5[2], addr_512_5, wires_2050_6,addr_2050_6);

wire[3:0] wires_2051_6;

wire[31:0] addr_2051_6;

Selector_2 s2051_6(wires_512_5[3], addr_512_5, wires_2051_6,addr_2051_6);

wire[3:0] wires_2052_6;

wire[31:0] addr_2052_6;

Selector_2 s2052_6(wires_513_5[0], addr_513_5, wires_2052_6,addr_2052_6);

wire[3:0] wires_2053_6;

wire[31:0] addr_2053_6;

Selector_2 s2053_6(wires_513_5[1], addr_513_5, wires_2053_6,addr_2053_6);

wire[3:0] wires_2054_6;

wire[31:0] addr_2054_6;

Selector_2 s2054_6(wires_513_5[2], addr_513_5, wires_2054_6,addr_2054_6);

wire[3:0] wires_2055_6;

wire[31:0] addr_2055_6;

Selector_2 s2055_6(wires_513_5[3], addr_513_5, wires_2055_6,addr_2055_6);

wire[3:0] wires_2056_6;

wire[31:0] addr_2056_6;

Selector_2 s2056_6(wires_514_5[0], addr_514_5, wires_2056_6,addr_2056_6);

wire[3:0] wires_2057_6;

wire[31:0] addr_2057_6;

Selector_2 s2057_6(wires_514_5[1], addr_514_5, wires_2057_6,addr_2057_6);

wire[3:0] wires_2058_6;

wire[31:0] addr_2058_6;

Selector_2 s2058_6(wires_514_5[2], addr_514_5, wires_2058_6,addr_2058_6);

wire[3:0] wires_2059_6;

wire[31:0] addr_2059_6;

Selector_2 s2059_6(wires_514_5[3], addr_514_5, wires_2059_6,addr_2059_6);

wire[3:0] wires_2060_6;

wire[31:0] addr_2060_6;

Selector_2 s2060_6(wires_515_5[0], addr_515_5, wires_2060_6,addr_2060_6);

wire[3:0] wires_2061_6;

wire[31:0] addr_2061_6;

Selector_2 s2061_6(wires_515_5[1], addr_515_5, wires_2061_6,addr_2061_6);

wire[3:0] wires_2062_6;

wire[31:0] addr_2062_6;

Selector_2 s2062_6(wires_515_5[2], addr_515_5, wires_2062_6,addr_2062_6);

wire[3:0] wires_2063_6;

wire[31:0] addr_2063_6;

Selector_2 s2063_6(wires_515_5[3], addr_515_5, wires_2063_6,addr_2063_6);

wire[3:0] wires_2064_6;

wire[31:0] addr_2064_6;

Selector_2 s2064_6(wires_516_5[0], addr_516_5, wires_2064_6,addr_2064_6);

wire[3:0] wires_2065_6;

wire[31:0] addr_2065_6;

Selector_2 s2065_6(wires_516_5[1], addr_516_5, wires_2065_6,addr_2065_6);

wire[3:0] wires_2066_6;

wire[31:0] addr_2066_6;

Selector_2 s2066_6(wires_516_5[2], addr_516_5, wires_2066_6,addr_2066_6);

wire[3:0] wires_2067_6;

wire[31:0] addr_2067_6;

Selector_2 s2067_6(wires_516_5[3], addr_516_5, wires_2067_6,addr_2067_6);

wire[3:0] wires_2068_6;

wire[31:0] addr_2068_6;

Selector_2 s2068_6(wires_517_5[0], addr_517_5, wires_2068_6,addr_2068_6);

wire[3:0] wires_2069_6;

wire[31:0] addr_2069_6;

Selector_2 s2069_6(wires_517_5[1], addr_517_5, wires_2069_6,addr_2069_6);

wire[3:0] wires_2070_6;

wire[31:0] addr_2070_6;

Selector_2 s2070_6(wires_517_5[2], addr_517_5, wires_2070_6,addr_2070_6);

wire[3:0] wires_2071_6;

wire[31:0] addr_2071_6;

Selector_2 s2071_6(wires_517_5[3], addr_517_5, wires_2071_6,addr_2071_6);

wire[3:0] wires_2072_6;

wire[31:0] addr_2072_6;

Selector_2 s2072_6(wires_518_5[0], addr_518_5, wires_2072_6,addr_2072_6);

wire[3:0] wires_2073_6;

wire[31:0] addr_2073_6;

Selector_2 s2073_6(wires_518_5[1], addr_518_5, wires_2073_6,addr_2073_6);

wire[3:0] wires_2074_6;

wire[31:0] addr_2074_6;

Selector_2 s2074_6(wires_518_5[2], addr_518_5, wires_2074_6,addr_2074_6);

wire[3:0] wires_2075_6;

wire[31:0] addr_2075_6;

Selector_2 s2075_6(wires_518_5[3], addr_518_5, wires_2075_6,addr_2075_6);

wire[3:0] wires_2076_6;

wire[31:0] addr_2076_6;

Selector_2 s2076_6(wires_519_5[0], addr_519_5, wires_2076_6,addr_2076_6);

wire[3:0] wires_2077_6;

wire[31:0] addr_2077_6;

Selector_2 s2077_6(wires_519_5[1], addr_519_5, wires_2077_6,addr_2077_6);

wire[3:0] wires_2078_6;

wire[31:0] addr_2078_6;

Selector_2 s2078_6(wires_519_5[2], addr_519_5, wires_2078_6,addr_2078_6);

wire[3:0] wires_2079_6;

wire[31:0] addr_2079_6;

Selector_2 s2079_6(wires_519_5[3], addr_519_5, wires_2079_6,addr_2079_6);

wire[3:0] wires_2080_6;

wire[31:0] addr_2080_6;

Selector_2 s2080_6(wires_520_5[0], addr_520_5, wires_2080_6,addr_2080_6);

wire[3:0] wires_2081_6;

wire[31:0] addr_2081_6;

Selector_2 s2081_6(wires_520_5[1], addr_520_5, wires_2081_6,addr_2081_6);

wire[3:0] wires_2082_6;

wire[31:0] addr_2082_6;

Selector_2 s2082_6(wires_520_5[2], addr_520_5, wires_2082_6,addr_2082_6);

wire[3:0] wires_2083_6;

wire[31:0] addr_2083_6;

Selector_2 s2083_6(wires_520_5[3], addr_520_5, wires_2083_6,addr_2083_6);

wire[3:0] wires_2084_6;

wire[31:0] addr_2084_6;

Selector_2 s2084_6(wires_521_5[0], addr_521_5, wires_2084_6,addr_2084_6);

wire[3:0] wires_2085_6;

wire[31:0] addr_2085_6;

Selector_2 s2085_6(wires_521_5[1], addr_521_5, wires_2085_6,addr_2085_6);

wire[3:0] wires_2086_6;

wire[31:0] addr_2086_6;

Selector_2 s2086_6(wires_521_5[2], addr_521_5, wires_2086_6,addr_2086_6);

wire[3:0] wires_2087_6;

wire[31:0] addr_2087_6;

Selector_2 s2087_6(wires_521_5[3], addr_521_5, wires_2087_6,addr_2087_6);

wire[3:0] wires_2088_6;

wire[31:0] addr_2088_6;

Selector_2 s2088_6(wires_522_5[0], addr_522_5, wires_2088_6,addr_2088_6);

wire[3:0] wires_2089_6;

wire[31:0] addr_2089_6;

Selector_2 s2089_6(wires_522_5[1], addr_522_5, wires_2089_6,addr_2089_6);

wire[3:0] wires_2090_6;

wire[31:0] addr_2090_6;

Selector_2 s2090_6(wires_522_5[2], addr_522_5, wires_2090_6,addr_2090_6);

wire[3:0] wires_2091_6;

wire[31:0] addr_2091_6;

Selector_2 s2091_6(wires_522_5[3], addr_522_5, wires_2091_6,addr_2091_6);

wire[3:0] wires_2092_6;

wire[31:0] addr_2092_6;

Selector_2 s2092_6(wires_523_5[0], addr_523_5, wires_2092_6,addr_2092_6);

wire[3:0] wires_2093_6;

wire[31:0] addr_2093_6;

Selector_2 s2093_6(wires_523_5[1], addr_523_5, wires_2093_6,addr_2093_6);

wire[3:0] wires_2094_6;

wire[31:0] addr_2094_6;

Selector_2 s2094_6(wires_523_5[2], addr_523_5, wires_2094_6,addr_2094_6);

wire[3:0] wires_2095_6;

wire[31:0] addr_2095_6;

Selector_2 s2095_6(wires_523_5[3], addr_523_5, wires_2095_6,addr_2095_6);

wire[3:0] wires_2096_6;

wire[31:0] addr_2096_6;

Selector_2 s2096_6(wires_524_5[0], addr_524_5, wires_2096_6,addr_2096_6);

wire[3:0] wires_2097_6;

wire[31:0] addr_2097_6;

Selector_2 s2097_6(wires_524_5[1], addr_524_5, wires_2097_6,addr_2097_6);

wire[3:0] wires_2098_6;

wire[31:0] addr_2098_6;

Selector_2 s2098_6(wires_524_5[2], addr_524_5, wires_2098_6,addr_2098_6);

wire[3:0] wires_2099_6;

wire[31:0] addr_2099_6;

Selector_2 s2099_6(wires_524_5[3], addr_524_5, wires_2099_6,addr_2099_6);

wire[3:0] wires_2100_6;

wire[31:0] addr_2100_6;

Selector_2 s2100_6(wires_525_5[0], addr_525_5, wires_2100_6,addr_2100_6);

wire[3:0] wires_2101_6;

wire[31:0] addr_2101_6;

Selector_2 s2101_6(wires_525_5[1], addr_525_5, wires_2101_6,addr_2101_6);

wire[3:0] wires_2102_6;

wire[31:0] addr_2102_6;

Selector_2 s2102_6(wires_525_5[2], addr_525_5, wires_2102_6,addr_2102_6);

wire[3:0] wires_2103_6;

wire[31:0] addr_2103_6;

Selector_2 s2103_6(wires_525_5[3], addr_525_5, wires_2103_6,addr_2103_6);

wire[3:0] wires_2104_6;

wire[31:0] addr_2104_6;

Selector_2 s2104_6(wires_526_5[0], addr_526_5, wires_2104_6,addr_2104_6);

wire[3:0] wires_2105_6;

wire[31:0] addr_2105_6;

Selector_2 s2105_6(wires_526_5[1], addr_526_5, wires_2105_6,addr_2105_6);

wire[3:0] wires_2106_6;

wire[31:0] addr_2106_6;

Selector_2 s2106_6(wires_526_5[2], addr_526_5, wires_2106_6,addr_2106_6);

wire[3:0] wires_2107_6;

wire[31:0] addr_2107_6;

Selector_2 s2107_6(wires_526_5[3], addr_526_5, wires_2107_6,addr_2107_6);

wire[3:0] wires_2108_6;

wire[31:0] addr_2108_6;

Selector_2 s2108_6(wires_527_5[0], addr_527_5, wires_2108_6,addr_2108_6);

wire[3:0] wires_2109_6;

wire[31:0] addr_2109_6;

Selector_2 s2109_6(wires_527_5[1], addr_527_5, wires_2109_6,addr_2109_6);

wire[3:0] wires_2110_6;

wire[31:0] addr_2110_6;

Selector_2 s2110_6(wires_527_5[2], addr_527_5, wires_2110_6,addr_2110_6);

wire[3:0] wires_2111_6;

wire[31:0] addr_2111_6;

Selector_2 s2111_6(wires_527_5[3], addr_527_5, wires_2111_6,addr_2111_6);

wire[3:0] wires_2112_6;

wire[31:0] addr_2112_6;

Selector_2 s2112_6(wires_528_5[0], addr_528_5, wires_2112_6,addr_2112_6);

wire[3:0] wires_2113_6;

wire[31:0] addr_2113_6;

Selector_2 s2113_6(wires_528_5[1], addr_528_5, wires_2113_6,addr_2113_6);

wire[3:0] wires_2114_6;

wire[31:0] addr_2114_6;

Selector_2 s2114_6(wires_528_5[2], addr_528_5, wires_2114_6,addr_2114_6);

wire[3:0] wires_2115_6;

wire[31:0] addr_2115_6;

Selector_2 s2115_6(wires_528_5[3], addr_528_5, wires_2115_6,addr_2115_6);

wire[3:0] wires_2116_6;

wire[31:0] addr_2116_6;

Selector_2 s2116_6(wires_529_5[0], addr_529_5, wires_2116_6,addr_2116_6);

wire[3:0] wires_2117_6;

wire[31:0] addr_2117_6;

Selector_2 s2117_6(wires_529_5[1], addr_529_5, wires_2117_6,addr_2117_6);

wire[3:0] wires_2118_6;

wire[31:0] addr_2118_6;

Selector_2 s2118_6(wires_529_5[2], addr_529_5, wires_2118_6,addr_2118_6);

wire[3:0] wires_2119_6;

wire[31:0] addr_2119_6;

Selector_2 s2119_6(wires_529_5[3], addr_529_5, wires_2119_6,addr_2119_6);

wire[3:0] wires_2120_6;

wire[31:0] addr_2120_6;

Selector_2 s2120_6(wires_530_5[0], addr_530_5, wires_2120_6,addr_2120_6);

wire[3:0] wires_2121_6;

wire[31:0] addr_2121_6;

Selector_2 s2121_6(wires_530_5[1], addr_530_5, wires_2121_6,addr_2121_6);

wire[3:0] wires_2122_6;

wire[31:0] addr_2122_6;

Selector_2 s2122_6(wires_530_5[2], addr_530_5, wires_2122_6,addr_2122_6);

wire[3:0] wires_2123_6;

wire[31:0] addr_2123_6;

Selector_2 s2123_6(wires_530_5[3], addr_530_5, wires_2123_6,addr_2123_6);

wire[3:0] wires_2124_6;

wire[31:0] addr_2124_6;

Selector_2 s2124_6(wires_531_5[0], addr_531_5, wires_2124_6,addr_2124_6);

wire[3:0] wires_2125_6;

wire[31:0] addr_2125_6;

Selector_2 s2125_6(wires_531_5[1], addr_531_5, wires_2125_6,addr_2125_6);

wire[3:0] wires_2126_6;

wire[31:0] addr_2126_6;

Selector_2 s2126_6(wires_531_5[2], addr_531_5, wires_2126_6,addr_2126_6);

wire[3:0] wires_2127_6;

wire[31:0] addr_2127_6;

Selector_2 s2127_6(wires_531_5[3], addr_531_5, wires_2127_6,addr_2127_6);

wire[3:0] wires_2128_6;

wire[31:0] addr_2128_6;

Selector_2 s2128_6(wires_532_5[0], addr_532_5, wires_2128_6,addr_2128_6);

wire[3:0] wires_2129_6;

wire[31:0] addr_2129_6;

Selector_2 s2129_6(wires_532_5[1], addr_532_5, wires_2129_6,addr_2129_6);

wire[3:0] wires_2130_6;

wire[31:0] addr_2130_6;

Selector_2 s2130_6(wires_532_5[2], addr_532_5, wires_2130_6,addr_2130_6);

wire[3:0] wires_2131_6;

wire[31:0] addr_2131_6;

Selector_2 s2131_6(wires_532_5[3], addr_532_5, wires_2131_6,addr_2131_6);

wire[3:0] wires_2132_6;

wire[31:0] addr_2132_6;

Selector_2 s2132_6(wires_533_5[0], addr_533_5, wires_2132_6,addr_2132_6);

wire[3:0] wires_2133_6;

wire[31:0] addr_2133_6;

Selector_2 s2133_6(wires_533_5[1], addr_533_5, wires_2133_6,addr_2133_6);

wire[3:0] wires_2134_6;

wire[31:0] addr_2134_6;

Selector_2 s2134_6(wires_533_5[2], addr_533_5, wires_2134_6,addr_2134_6);

wire[3:0] wires_2135_6;

wire[31:0] addr_2135_6;

Selector_2 s2135_6(wires_533_5[3], addr_533_5, wires_2135_6,addr_2135_6);

wire[3:0] wires_2136_6;

wire[31:0] addr_2136_6;

Selector_2 s2136_6(wires_534_5[0], addr_534_5, wires_2136_6,addr_2136_6);

wire[3:0] wires_2137_6;

wire[31:0] addr_2137_6;

Selector_2 s2137_6(wires_534_5[1], addr_534_5, wires_2137_6,addr_2137_6);

wire[3:0] wires_2138_6;

wire[31:0] addr_2138_6;

Selector_2 s2138_6(wires_534_5[2], addr_534_5, wires_2138_6,addr_2138_6);

wire[3:0] wires_2139_6;

wire[31:0] addr_2139_6;

Selector_2 s2139_6(wires_534_5[3], addr_534_5, wires_2139_6,addr_2139_6);

wire[3:0] wires_2140_6;

wire[31:0] addr_2140_6;

Selector_2 s2140_6(wires_535_5[0], addr_535_5, wires_2140_6,addr_2140_6);

wire[3:0] wires_2141_6;

wire[31:0] addr_2141_6;

Selector_2 s2141_6(wires_535_5[1], addr_535_5, wires_2141_6,addr_2141_6);

wire[3:0] wires_2142_6;

wire[31:0] addr_2142_6;

Selector_2 s2142_6(wires_535_5[2], addr_535_5, wires_2142_6,addr_2142_6);

wire[3:0] wires_2143_6;

wire[31:0] addr_2143_6;

Selector_2 s2143_6(wires_535_5[3], addr_535_5, wires_2143_6,addr_2143_6);

wire[3:0] wires_2144_6;

wire[31:0] addr_2144_6;

Selector_2 s2144_6(wires_536_5[0], addr_536_5, wires_2144_6,addr_2144_6);

wire[3:0] wires_2145_6;

wire[31:0] addr_2145_6;

Selector_2 s2145_6(wires_536_5[1], addr_536_5, wires_2145_6,addr_2145_6);

wire[3:0] wires_2146_6;

wire[31:0] addr_2146_6;

Selector_2 s2146_6(wires_536_5[2], addr_536_5, wires_2146_6,addr_2146_6);

wire[3:0] wires_2147_6;

wire[31:0] addr_2147_6;

Selector_2 s2147_6(wires_536_5[3], addr_536_5, wires_2147_6,addr_2147_6);

wire[3:0] wires_2148_6;

wire[31:0] addr_2148_6;

Selector_2 s2148_6(wires_537_5[0], addr_537_5, wires_2148_6,addr_2148_6);

wire[3:0] wires_2149_6;

wire[31:0] addr_2149_6;

Selector_2 s2149_6(wires_537_5[1], addr_537_5, wires_2149_6,addr_2149_6);

wire[3:0] wires_2150_6;

wire[31:0] addr_2150_6;

Selector_2 s2150_6(wires_537_5[2], addr_537_5, wires_2150_6,addr_2150_6);

wire[3:0] wires_2151_6;

wire[31:0] addr_2151_6;

Selector_2 s2151_6(wires_537_5[3], addr_537_5, wires_2151_6,addr_2151_6);

wire[3:0] wires_2152_6;

wire[31:0] addr_2152_6;

Selector_2 s2152_6(wires_538_5[0], addr_538_5, wires_2152_6,addr_2152_6);

wire[3:0] wires_2153_6;

wire[31:0] addr_2153_6;

Selector_2 s2153_6(wires_538_5[1], addr_538_5, wires_2153_6,addr_2153_6);

wire[3:0] wires_2154_6;

wire[31:0] addr_2154_6;

Selector_2 s2154_6(wires_538_5[2], addr_538_5, wires_2154_6,addr_2154_6);

wire[3:0] wires_2155_6;

wire[31:0] addr_2155_6;

Selector_2 s2155_6(wires_538_5[3], addr_538_5, wires_2155_6,addr_2155_6);

wire[3:0] wires_2156_6;

wire[31:0] addr_2156_6;

Selector_2 s2156_6(wires_539_5[0], addr_539_5, wires_2156_6,addr_2156_6);

wire[3:0] wires_2157_6;

wire[31:0] addr_2157_6;

Selector_2 s2157_6(wires_539_5[1], addr_539_5, wires_2157_6,addr_2157_6);

wire[3:0] wires_2158_6;

wire[31:0] addr_2158_6;

Selector_2 s2158_6(wires_539_5[2], addr_539_5, wires_2158_6,addr_2158_6);

wire[3:0] wires_2159_6;

wire[31:0] addr_2159_6;

Selector_2 s2159_6(wires_539_5[3], addr_539_5, wires_2159_6,addr_2159_6);

wire[3:0] wires_2160_6;

wire[31:0] addr_2160_6;

Selector_2 s2160_6(wires_540_5[0], addr_540_5, wires_2160_6,addr_2160_6);

wire[3:0] wires_2161_6;

wire[31:0] addr_2161_6;

Selector_2 s2161_6(wires_540_5[1], addr_540_5, wires_2161_6,addr_2161_6);

wire[3:0] wires_2162_6;

wire[31:0] addr_2162_6;

Selector_2 s2162_6(wires_540_5[2], addr_540_5, wires_2162_6,addr_2162_6);

wire[3:0] wires_2163_6;

wire[31:0] addr_2163_6;

Selector_2 s2163_6(wires_540_5[3], addr_540_5, wires_2163_6,addr_2163_6);

wire[3:0] wires_2164_6;

wire[31:0] addr_2164_6;

Selector_2 s2164_6(wires_541_5[0], addr_541_5, wires_2164_6,addr_2164_6);

wire[3:0] wires_2165_6;

wire[31:0] addr_2165_6;

Selector_2 s2165_6(wires_541_5[1], addr_541_5, wires_2165_6,addr_2165_6);

wire[3:0] wires_2166_6;

wire[31:0] addr_2166_6;

Selector_2 s2166_6(wires_541_5[2], addr_541_5, wires_2166_6,addr_2166_6);

wire[3:0] wires_2167_6;

wire[31:0] addr_2167_6;

Selector_2 s2167_6(wires_541_5[3], addr_541_5, wires_2167_6,addr_2167_6);

wire[3:0] wires_2168_6;

wire[31:0] addr_2168_6;

Selector_2 s2168_6(wires_542_5[0], addr_542_5, wires_2168_6,addr_2168_6);

wire[3:0] wires_2169_6;

wire[31:0] addr_2169_6;

Selector_2 s2169_6(wires_542_5[1], addr_542_5, wires_2169_6,addr_2169_6);

wire[3:0] wires_2170_6;

wire[31:0] addr_2170_6;

Selector_2 s2170_6(wires_542_5[2], addr_542_5, wires_2170_6,addr_2170_6);

wire[3:0] wires_2171_6;

wire[31:0] addr_2171_6;

Selector_2 s2171_6(wires_542_5[3], addr_542_5, wires_2171_6,addr_2171_6);

wire[3:0] wires_2172_6;

wire[31:0] addr_2172_6;

Selector_2 s2172_6(wires_543_5[0], addr_543_5, wires_2172_6,addr_2172_6);

wire[3:0] wires_2173_6;

wire[31:0] addr_2173_6;

Selector_2 s2173_6(wires_543_5[1], addr_543_5, wires_2173_6,addr_2173_6);

wire[3:0] wires_2174_6;

wire[31:0] addr_2174_6;

Selector_2 s2174_6(wires_543_5[2], addr_543_5, wires_2174_6,addr_2174_6);

wire[3:0] wires_2175_6;

wire[31:0] addr_2175_6;

Selector_2 s2175_6(wires_543_5[3], addr_543_5, wires_2175_6,addr_2175_6);

wire[3:0] wires_2176_6;

wire[31:0] addr_2176_6;

Selector_2 s2176_6(wires_544_5[0], addr_544_5, wires_2176_6,addr_2176_6);

wire[3:0] wires_2177_6;

wire[31:0] addr_2177_6;

Selector_2 s2177_6(wires_544_5[1], addr_544_5, wires_2177_6,addr_2177_6);

wire[3:0] wires_2178_6;

wire[31:0] addr_2178_6;

Selector_2 s2178_6(wires_544_5[2], addr_544_5, wires_2178_6,addr_2178_6);

wire[3:0] wires_2179_6;

wire[31:0] addr_2179_6;

Selector_2 s2179_6(wires_544_5[3], addr_544_5, wires_2179_6,addr_2179_6);

wire[3:0] wires_2180_6;

wire[31:0] addr_2180_6;

Selector_2 s2180_6(wires_545_5[0], addr_545_5, wires_2180_6,addr_2180_6);

wire[3:0] wires_2181_6;

wire[31:0] addr_2181_6;

Selector_2 s2181_6(wires_545_5[1], addr_545_5, wires_2181_6,addr_2181_6);

wire[3:0] wires_2182_6;

wire[31:0] addr_2182_6;

Selector_2 s2182_6(wires_545_5[2], addr_545_5, wires_2182_6,addr_2182_6);

wire[3:0] wires_2183_6;

wire[31:0] addr_2183_6;

Selector_2 s2183_6(wires_545_5[3], addr_545_5, wires_2183_6,addr_2183_6);

wire[3:0] wires_2184_6;

wire[31:0] addr_2184_6;

Selector_2 s2184_6(wires_546_5[0], addr_546_5, wires_2184_6,addr_2184_6);

wire[3:0] wires_2185_6;

wire[31:0] addr_2185_6;

Selector_2 s2185_6(wires_546_5[1], addr_546_5, wires_2185_6,addr_2185_6);

wire[3:0] wires_2186_6;

wire[31:0] addr_2186_6;

Selector_2 s2186_6(wires_546_5[2], addr_546_5, wires_2186_6,addr_2186_6);

wire[3:0] wires_2187_6;

wire[31:0] addr_2187_6;

Selector_2 s2187_6(wires_546_5[3], addr_546_5, wires_2187_6,addr_2187_6);

wire[3:0] wires_2188_6;

wire[31:0] addr_2188_6;

Selector_2 s2188_6(wires_547_5[0], addr_547_5, wires_2188_6,addr_2188_6);

wire[3:0] wires_2189_6;

wire[31:0] addr_2189_6;

Selector_2 s2189_6(wires_547_5[1], addr_547_5, wires_2189_6,addr_2189_6);

wire[3:0] wires_2190_6;

wire[31:0] addr_2190_6;

Selector_2 s2190_6(wires_547_5[2], addr_547_5, wires_2190_6,addr_2190_6);

wire[3:0] wires_2191_6;

wire[31:0] addr_2191_6;

Selector_2 s2191_6(wires_547_5[3], addr_547_5, wires_2191_6,addr_2191_6);

wire[3:0] wires_2192_6;

wire[31:0] addr_2192_6;

Selector_2 s2192_6(wires_548_5[0], addr_548_5, wires_2192_6,addr_2192_6);

wire[3:0] wires_2193_6;

wire[31:0] addr_2193_6;

Selector_2 s2193_6(wires_548_5[1], addr_548_5, wires_2193_6,addr_2193_6);

wire[3:0] wires_2194_6;

wire[31:0] addr_2194_6;

Selector_2 s2194_6(wires_548_5[2], addr_548_5, wires_2194_6,addr_2194_6);

wire[3:0] wires_2195_6;

wire[31:0] addr_2195_6;

Selector_2 s2195_6(wires_548_5[3], addr_548_5, wires_2195_6,addr_2195_6);

wire[3:0] wires_2196_6;

wire[31:0] addr_2196_6;

Selector_2 s2196_6(wires_549_5[0], addr_549_5, wires_2196_6,addr_2196_6);

wire[3:0] wires_2197_6;

wire[31:0] addr_2197_6;

Selector_2 s2197_6(wires_549_5[1], addr_549_5, wires_2197_6,addr_2197_6);

wire[3:0] wires_2198_6;

wire[31:0] addr_2198_6;

Selector_2 s2198_6(wires_549_5[2], addr_549_5, wires_2198_6,addr_2198_6);

wire[3:0] wires_2199_6;

wire[31:0] addr_2199_6;

Selector_2 s2199_6(wires_549_5[3], addr_549_5, wires_2199_6,addr_2199_6);

wire[3:0] wires_2200_6;

wire[31:0] addr_2200_6;

Selector_2 s2200_6(wires_550_5[0], addr_550_5, wires_2200_6,addr_2200_6);

wire[3:0] wires_2201_6;

wire[31:0] addr_2201_6;

Selector_2 s2201_6(wires_550_5[1], addr_550_5, wires_2201_6,addr_2201_6);

wire[3:0] wires_2202_6;

wire[31:0] addr_2202_6;

Selector_2 s2202_6(wires_550_5[2], addr_550_5, wires_2202_6,addr_2202_6);

wire[3:0] wires_2203_6;

wire[31:0] addr_2203_6;

Selector_2 s2203_6(wires_550_5[3], addr_550_5, wires_2203_6,addr_2203_6);

wire[3:0] wires_2204_6;

wire[31:0] addr_2204_6;

Selector_2 s2204_6(wires_551_5[0], addr_551_5, wires_2204_6,addr_2204_6);

wire[3:0] wires_2205_6;

wire[31:0] addr_2205_6;

Selector_2 s2205_6(wires_551_5[1], addr_551_5, wires_2205_6,addr_2205_6);

wire[3:0] wires_2206_6;

wire[31:0] addr_2206_6;

Selector_2 s2206_6(wires_551_5[2], addr_551_5, wires_2206_6,addr_2206_6);

wire[3:0] wires_2207_6;

wire[31:0] addr_2207_6;

Selector_2 s2207_6(wires_551_5[3], addr_551_5, wires_2207_6,addr_2207_6);

wire[3:0] wires_2208_6;

wire[31:0] addr_2208_6;

Selector_2 s2208_6(wires_552_5[0], addr_552_5, wires_2208_6,addr_2208_6);

wire[3:0] wires_2209_6;

wire[31:0] addr_2209_6;

Selector_2 s2209_6(wires_552_5[1], addr_552_5, wires_2209_6,addr_2209_6);

wire[3:0] wires_2210_6;

wire[31:0] addr_2210_6;

Selector_2 s2210_6(wires_552_5[2], addr_552_5, wires_2210_6,addr_2210_6);

wire[3:0] wires_2211_6;

wire[31:0] addr_2211_6;

Selector_2 s2211_6(wires_552_5[3], addr_552_5, wires_2211_6,addr_2211_6);

wire[3:0] wires_2212_6;

wire[31:0] addr_2212_6;

Selector_2 s2212_6(wires_553_5[0], addr_553_5, wires_2212_6,addr_2212_6);

wire[3:0] wires_2213_6;

wire[31:0] addr_2213_6;

Selector_2 s2213_6(wires_553_5[1], addr_553_5, wires_2213_6,addr_2213_6);

wire[3:0] wires_2214_6;

wire[31:0] addr_2214_6;

Selector_2 s2214_6(wires_553_5[2], addr_553_5, wires_2214_6,addr_2214_6);

wire[3:0] wires_2215_6;

wire[31:0] addr_2215_6;

Selector_2 s2215_6(wires_553_5[3], addr_553_5, wires_2215_6,addr_2215_6);

wire[3:0] wires_2216_6;

wire[31:0] addr_2216_6;

Selector_2 s2216_6(wires_554_5[0], addr_554_5, wires_2216_6,addr_2216_6);

wire[3:0] wires_2217_6;

wire[31:0] addr_2217_6;

Selector_2 s2217_6(wires_554_5[1], addr_554_5, wires_2217_6,addr_2217_6);

wire[3:0] wires_2218_6;

wire[31:0] addr_2218_6;

Selector_2 s2218_6(wires_554_5[2], addr_554_5, wires_2218_6,addr_2218_6);

wire[3:0] wires_2219_6;

wire[31:0] addr_2219_6;

Selector_2 s2219_6(wires_554_5[3], addr_554_5, wires_2219_6,addr_2219_6);

wire[3:0] wires_2220_6;

wire[31:0] addr_2220_6;

Selector_2 s2220_6(wires_555_5[0], addr_555_5, wires_2220_6,addr_2220_6);

wire[3:0] wires_2221_6;

wire[31:0] addr_2221_6;

Selector_2 s2221_6(wires_555_5[1], addr_555_5, wires_2221_6,addr_2221_6);

wire[3:0] wires_2222_6;

wire[31:0] addr_2222_6;

Selector_2 s2222_6(wires_555_5[2], addr_555_5, wires_2222_6,addr_2222_6);

wire[3:0] wires_2223_6;

wire[31:0] addr_2223_6;

Selector_2 s2223_6(wires_555_5[3], addr_555_5, wires_2223_6,addr_2223_6);

wire[3:0] wires_2224_6;

wire[31:0] addr_2224_6;

Selector_2 s2224_6(wires_556_5[0], addr_556_5, wires_2224_6,addr_2224_6);

wire[3:0] wires_2225_6;

wire[31:0] addr_2225_6;

Selector_2 s2225_6(wires_556_5[1], addr_556_5, wires_2225_6,addr_2225_6);

wire[3:0] wires_2226_6;

wire[31:0] addr_2226_6;

Selector_2 s2226_6(wires_556_5[2], addr_556_5, wires_2226_6,addr_2226_6);

wire[3:0] wires_2227_6;

wire[31:0] addr_2227_6;

Selector_2 s2227_6(wires_556_5[3], addr_556_5, wires_2227_6,addr_2227_6);

wire[3:0] wires_2228_6;

wire[31:0] addr_2228_6;

Selector_2 s2228_6(wires_557_5[0], addr_557_5, wires_2228_6,addr_2228_6);

wire[3:0] wires_2229_6;

wire[31:0] addr_2229_6;

Selector_2 s2229_6(wires_557_5[1], addr_557_5, wires_2229_6,addr_2229_6);

wire[3:0] wires_2230_6;

wire[31:0] addr_2230_6;

Selector_2 s2230_6(wires_557_5[2], addr_557_5, wires_2230_6,addr_2230_6);

wire[3:0] wires_2231_6;

wire[31:0] addr_2231_6;

Selector_2 s2231_6(wires_557_5[3], addr_557_5, wires_2231_6,addr_2231_6);

wire[3:0] wires_2232_6;

wire[31:0] addr_2232_6;

Selector_2 s2232_6(wires_558_5[0], addr_558_5, wires_2232_6,addr_2232_6);

wire[3:0] wires_2233_6;

wire[31:0] addr_2233_6;

Selector_2 s2233_6(wires_558_5[1], addr_558_5, wires_2233_6,addr_2233_6);

wire[3:0] wires_2234_6;

wire[31:0] addr_2234_6;

Selector_2 s2234_6(wires_558_5[2], addr_558_5, wires_2234_6,addr_2234_6);

wire[3:0] wires_2235_6;

wire[31:0] addr_2235_6;

Selector_2 s2235_6(wires_558_5[3], addr_558_5, wires_2235_6,addr_2235_6);

wire[3:0] wires_2236_6;

wire[31:0] addr_2236_6;

Selector_2 s2236_6(wires_559_5[0], addr_559_5, wires_2236_6,addr_2236_6);

wire[3:0] wires_2237_6;

wire[31:0] addr_2237_6;

Selector_2 s2237_6(wires_559_5[1], addr_559_5, wires_2237_6,addr_2237_6);

wire[3:0] wires_2238_6;

wire[31:0] addr_2238_6;

Selector_2 s2238_6(wires_559_5[2], addr_559_5, wires_2238_6,addr_2238_6);

wire[3:0] wires_2239_6;

wire[31:0] addr_2239_6;

Selector_2 s2239_6(wires_559_5[3], addr_559_5, wires_2239_6,addr_2239_6);

wire[3:0] wires_2240_6;

wire[31:0] addr_2240_6;

Selector_2 s2240_6(wires_560_5[0], addr_560_5, wires_2240_6,addr_2240_6);

wire[3:0] wires_2241_6;

wire[31:0] addr_2241_6;

Selector_2 s2241_6(wires_560_5[1], addr_560_5, wires_2241_6,addr_2241_6);

wire[3:0] wires_2242_6;

wire[31:0] addr_2242_6;

Selector_2 s2242_6(wires_560_5[2], addr_560_5, wires_2242_6,addr_2242_6);

wire[3:0] wires_2243_6;

wire[31:0] addr_2243_6;

Selector_2 s2243_6(wires_560_5[3], addr_560_5, wires_2243_6,addr_2243_6);

wire[3:0] wires_2244_6;

wire[31:0] addr_2244_6;

Selector_2 s2244_6(wires_561_5[0], addr_561_5, wires_2244_6,addr_2244_6);

wire[3:0] wires_2245_6;

wire[31:0] addr_2245_6;

Selector_2 s2245_6(wires_561_5[1], addr_561_5, wires_2245_6,addr_2245_6);

wire[3:0] wires_2246_6;

wire[31:0] addr_2246_6;

Selector_2 s2246_6(wires_561_5[2], addr_561_5, wires_2246_6,addr_2246_6);

wire[3:0] wires_2247_6;

wire[31:0] addr_2247_6;

Selector_2 s2247_6(wires_561_5[3], addr_561_5, wires_2247_6,addr_2247_6);

wire[3:0] wires_2248_6;

wire[31:0] addr_2248_6;

Selector_2 s2248_6(wires_562_5[0], addr_562_5, wires_2248_6,addr_2248_6);

wire[3:0] wires_2249_6;

wire[31:0] addr_2249_6;

Selector_2 s2249_6(wires_562_5[1], addr_562_5, wires_2249_6,addr_2249_6);

wire[3:0] wires_2250_6;

wire[31:0] addr_2250_6;

Selector_2 s2250_6(wires_562_5[2], addr_562_5, wires_2250_6,addr_2250_6);

wire[3:0] wires_2251_6;

wire[31:0] addr_2251_6;

Selector_2 s2251_6(wires_562_5[3], addr_562_5, wires_2251_6,addr_2251_6);

wire[3:0] wires_2252_6;

wire[31:0] addr_2252_6;

Selector_2 s2252_6(wires_563_5[0], addr_563_5, wires_2252_6,addr_2252_6);

wire[3:0] wires_2253_6;

wire[31:0] addr_2253_6;

Selector_2 s2253_6(wires_563_5[1], addr_563_5, wires_2253_6,addr_2253_6);

wire[3:0] wires_2254_6;

wire[31:0] addr_2254_6;

Selector_2 s2254_6(wires_563_5[2], addr_563_5, wires_2254_6,addr_2254_6);

wire[3:0] wires_2255_6;

wire[31:0] addr_2255_6;

Selector_2 s2255_6(wires_563_5[3], addr_563_5, wires_2255_6,addr_2255_6);

wire[3:0] wires_2256_6;

wire[31:0] addr_2256_6;

Selector_2 s2256_6(wires_564_5[0], addr_564_5, wires_2256_6,addr_2256_6);

wire[3:0] wires_2257_6;

wire[31:0] addr_2257_6;

Selector_2 s2257_6(wires_564_5[1], addr_564_5, wires_2257_6,addr_2257_6);

wire[3:0] wires_2258_6;

wire[31:0] addr_2258_6;

Selector_2 s2258_6(wires_564_5[2], addr_564_5, wires_2258_6,addr_2258_6);

wire[3:0] wires_2259_6;

wire[31:0] addr_2259_6;

Selector_2 s2259_6(wires_564_5[3], addr_564_5, wires_2259_6,addr_2259_6);

wire[3:0] wires_2260_6;

wire[31:0] addr_2260_6;

Selector_2 s2260_6(wires_565_5[0], addr_565_5, wires_2260_6,addr_2260_6);

wire[3:0] wires_2261_6;

wire[31:0] addr_2261_6;

Selector_2 s2261_6(wires_565_5[1], addr_565_5, wires_2261_6,addr_2261_6);

wire[3:0] wires_2262_6;

wire[31:0] addr_2262_6;

Selector_2 s2262_6(wires_565_5[2], addr_565_5, wires_2262_6,addr_2262_6);

wire[3:0] wires_2263_6;

wire[31:0] addr_2263_6;

Selector_2 s2263_6(wires_565_5[3], addr_565_5, wires_2263_6,addr_2263_6);

wire[3:0] wires_2264_6;

wire[31:0] addr_2264_6;

Selector_2 s2264_6(wires_566_5[0], addr_566_5, wires_2264_6,addr_2264_6);

wire[3:0] wires_2265_6;

wire[31:0] addr_2265_6;

Selector_2 s2265_6(wires_566_5[1], addr_566_5, wires_2265_6,addr_2265_6);

wire[3:0] wires_2266_6;

wire[31:0] addr_2266_6;

Selector_2 s2266_6(wires_566_5[2], addr_566_5, wires_2266_6,addr_2266_6);

wire[3:0] wires_2267_6;

wire[31:0] addr_2267_6;

Selector_2 s2267_6(wires_566_5[3], addr_566_5, wires_2267_6,addr_2267_6);

wire[3:0] wires_2268_6;

wire[31:0] addr_2268_6;

Selector_2 s2268_6(wires_567_5[0], addr_567_5, wires_2268_6,addr_2268_6);

wire[3:0] wires_2269_6;

wire[31:0] addr_2269_6;

Selector_2 s2269_6(wires_567_5[1], addr_567_5, wires_2269_6,addr_2269_6);

wire[3:0] wires_2270_6;

wire[31:0] addr_2270_6;

Selector_2 s2270_6(wires_567_5[2], addr_567_5, wires_2270_6,addr_2270_6);

wire[3:0] wires_2271_6;

wire[31:0] addr_2271_6;

Selector_2 s2271_6(wires_567_5[3], addr_567_5, wires_2271_6,addr_2271_6);

wire[3:0] wires_2272_6;

wire[31:0] addr_2272_6;

Selector_2 s2272_6(wires_568_5[0], addr_568_5, wires_2272_6,addr_2272_6);

wire[3:0] wires_2273_6;

wire[31:0] addr_2273_6;

Selector_2 s2273_6(wires_568_5[1], addr_568_5, wires_2273_6,addr_2273_6);

wire[3:0] wires_2274_6;

wire[31:0] addr_2274_6;

Selector_2 s2274_6(wires_568_5[2], addr_568_5, wires_2274_6,addr_2274_6);

wire[3:0] wires_2275_6;

wire[31:0] addr_2275_6;

Selector_2 s2275_6(wires_568_5[3], addr_568_5, wires_2275_6,addr_2275_6);

wire[3:0] wires_2276_6;

wire[31:0] addr_2276_6;

Selector_2 s2276_6(wires_569_5[0], addr_569_5, wires_2276_6,addr_2276_6);

wire[3:0] wires_2277_6;

wire[31:0] addr_2277_6;

Selector_2 s2277_6(wires_569_5[1], addr_569_5, wires_2277_6,addr_2277_6);

wire[3:0] wires_2278_6;

wire[31:0] addr_2278_6;

Selector_2 s2278_6(wires_569_5[2], addr_569_5, wires_2278_6,addr_2278_6);

wire[3:0] wires_2279_6;

wire[31:0] addr_2279_6;

Selector_2 s2279_6(wires_569_5[3], addr_569_5, wires_2279_6,addr_2279_6);

wire[3:0] wires_2280_6;

wire[31:0] addr_2280_6;

Selector_2 s2280_6(wires_570_5[0], addr_570_5, wires_2280_6,addr_2280_6);

wire[3:0] wires_2281_6;

wire[31:0] addr_2281_6;

Selector_2 s2281_6(wires_570_5[1], addr_570_5, wires_2281_6,addr_2281_6);

wire[3:0] wires_2282_6;

wire[31:0] addr_2282_6;

Selector_2 s2282_6(wires_570_5[2], addr_570_5, wires_2282_6,addr_2282_6);

wire[3:0] wires_2283_6;

wire[31:0] addr_2283_6;

Selector_2 s2283_6(wires_570_5[3], addr_570_5, wires_2283_6,addr_2283_6);

wire[3:0] wires_2284_6;

wire[31:0] addr_2284_6;

Selector_2 s2284_6(wires_571_5[0], addr_571_5, wires_2284_6,addr_2284_6);

wire[3:0] wires_2285_6;

wire[31:0] addr_2285_6;

Selector_2 s2285_6(wires_571_5[1], addr_571_5, wires_2285_6,addr_2285_6);

wire[3:0] wires_2286_6;

wire[31:0] addr_2286_6;

Selector_2 s2286_6(wires_571_5[2], addr_571_5, wires_2286_6,addr_2286_6);

wire[3:0] wires_2287_6;

wire[31:0] addr_2287_6;

Selector_2 s2287_6(wires_571_5[3], addr_571_5, wires_2287_6,addr_2287_6);

wire[3:0] wires_2288_6;

wire[31:0] addr_2288_6;

Selector_2 s2288_6(wires_572_5[0], addr_572_5, wires_2288_6,addr_2288_6);

wire[3:0] wires_2289_6;

wire[31:0] addr_2289_6;

Selector_2 s2289_6(wires_572_5[1], addr_572_5, wires_2289_6,addr_2289_6);

wire[3:0] wires_2290_6;

wire[31:0] addr_2290_6;

Selector_2 s2290_6(wires_572_5[2], addr_572_5, wires_2290_6,addr_2290_6);

wire[3:0] wires_2291_6;

wire[31:0] addr_2291_6;

Selector_2 s2291_6(wires_572_5[3], addr_572_5, wires_2291_6,addr_2291_6);

wire[3:0] wires_2292_6;

wire[31:0] addr_2292_6;

Selector_2 s2292_6(wires_573_5[0], addr_573_5, wires_2292_6,addr_2292_6);

wire[3:0] wires_2293_6;

wire[31:0] addr_2293_6;

Selector_2 s2293_6(wires_573_5[1], addr_573_5, wires_2293_6,addr_2293_6);

wire[3:0] wires_2294_6;

wire[31:0] addr_2294_6;

Selector_2 s2294_6(wires_573_5[2], addr_573_5, wires_2294_6,addr_2294_6);

wire[3:0] wires_2295_6;

wire[31:0] addr_2295_6;

Selector_2 s2295_6(wires_573_5[3], addr_573_5, wires_2295_6,addr_2295_6);

wire[3:0] wires_2296_6;

wire[31:0] addr_2296_6;

Selector_2 s2296_6(wires_574_5[0], addr_574_5, wires_2296_6,addr_2296_6);

wire[3:0] wires_2297_6;

wire[31:0] addr_2297_6;

Selector_2 s2297_6(wires_574_5[1], addr_574_5, wires_2297_6,addr_2297_6);

wire[3:0] wires_2298_6;

wire[31:0] addr_2298_6;

Selector_2 s2298_6(wires_574_5[2], addr_574_5, wires_2298_6,addr_2298_6);

wire[3:0] wires_2299_6;

wire[31:0] addr_2299_6;

Selector_2 s2299_6(wires_574_5[3], addr_574_5, wires_2299_6,addr_2299_6);

wire[3:0] wires_2300_6;

wire[31:0] addr_2300_6;

Selector_2 s2300_6(wires_575_5[0], addr_575_5, wires_2300_6,addr_2300_6);

wire[3:0] wires_2301_6;

wire[31:0] addr_2301_6;

Selector_2 s2301_6(wires_575_5[1], addr_575_5, wires_2301_6,addr_2301_6);

wire[3:0] wires_2302_6;

wire[31:0] addr_2302_6;

Selector_2 s2302_6(wires_575_5[2], addr_575_5, wires_2302_6,addr_2302_6);

wire[3:0] wires_2303_6;

wire[31:0] addr_2303_6;

Selector_2 s2303_6(wires_575_5[3], addr_575_5, wires_2303_6,addr_2303_6);

wire[3:0] wires_2304_6;

wire[31:0] addr_2304_6;

Selector_2 s2304_6(wires_576_5[0], addr_576_5, wires_2304_6,addr_2304_6);

wire[3:0] wires_2305_6;

wire[31:0] addr_2305_6;

Selector_2 s2305_6(wires_576_5[1], addr_576_5, wires_2305_6,addr_2305_6);

wire[3:0] wires_2306_6;

wire[31:0] addr_2306_6;

Selector_2 s2306_6(wires_576_5[2], addr_576_5, wires_2306_6,addr_2306_6);

wire[3:0] wires_2307_6;

wire[31:0] addr_2307_6;

Selector_2 s2307_6(wires_576_5[3], addr_576_5, wires_2307_6,addr_2307_6);

wire[3:0] wires_2308_6;

wire[31:0] addr_2308_6;

Selector_2 s2308_6(wires_577_5[0], addr_577_5, wires_2308_6,addr_2308_6);

wire[3:0] wires_2309_6;

wire[31:0] addr_2309_6;

Selector_2 s2309_6(wires_577_5[1], addr_577_5, wires_2309_6,addr_2309_6);

wire[3:0] wires_2310_6;

wire[31:0] addr_2310_6;

Selector_2 s2310_6(wires_577_5[2], addr_577_5, wires_2310_6,addr_2310_6);

wire[3:0] wires_2311_6;

wire[31:0] addr_2311_6;

Selector_2 s2311_6(wires_577_5[3], addr_577_5, wires_2311_6,addr_2311_6);

wire[3:0] wires_2312_6;

wire[31:0] addr_2312_6;

Selector_2 s2312_6(wires_578_5[0], addr_578_5, wires_2312_6,addr_2312_6);

wire[3:0] wires_2313_6;

wire[31:0] addr_2313_6;

Selector_2 s2313_6(wires_578_5[1], addr_578_5, wires_2313_6,addr_2313_6);

wire[3:0] wires_2314_6;

wire[31:0] addr_2314_6;

Selector_2 s2314_6(wires_578_5[2], addr_578_5, wires_2314_6,addr_2314_6);

wire[3:0] wires_2315_6;

wire[31:0] addr_2315_6;

Selector_2 s2315_6(wires_578_5[3], addr_578_5, wires_2315_6,addr_2315_6);

wire[3:0] wires_2316_6;

wire[31:0] addr_2316_6;

Selector_2 s2316_6(wires_579_5[0], addr_579_5, wires_2316_6,addr_2316_6);

wire[3:0] wires_2317_6;

wire[31:0] addr_2317_6;

Selector_2 s2317_6(wires_579_5[1], addr_579_5, wires_2317_6,addr_2317_6);

wire[3:0] wires_2318_6;

wire[31:0] addr_2318_6;

Selector_2 s2318_6(wires_579_5[2], addr_579_5, wires_2318_6,addr_2318_6);

wire[3:0] wires_2319_6;

wire[31:0] addr_2319_6;

Selector_2 s2319_6(wires_579_5[3], addr_579_5, wires_2319_6,addr_2319_6);

wire[3:0] wires_2320_6;

wire[31:0] addr_2320_6;

Selector_2 s2320_6(wires_580_5[0], addr_580_5, wires_2320_6,addr_2320_6);

wire[3:0] wires_2321_6;

wire[31:0] addr_2321_6;

Selector_2 s2321_6(wires_580_5[1], addr_580_5, wires_2321_6,addr_2321_6);

wire[3:0] wires_2322_6;

wire[31:0] addr_2322_6;

Selector_2 s2322_6(wires_580_5[2], addr_580_5, wires_2322_6,addr_2322_6);

wire[3:0] wires_2323_6;

wire[31:0] addr_2323_6;

Selector_2 s2323_6(wires_580_5[3], addr_580_5, wires_2323_6,addr_2323_6);

wire[3:0] wires_2324_6;

wire[31:0] addr_2324_6;

Selector_2 s2324_6(wires_581_5[0], addr_581_5, wires_2324_6,addr_2324_6);

wire[3:0] wires_2325_6;

wire[31:0] addr_2325_6;

Selector_2 s2325_6(wires_581_5[1], addr_581_5, wires_2325_6,addr_2325_6);

wire[3:0] wires_2326_6;

wire[31:0] addr_2326_6;

Selector_2 s2326_6(wires_581_5[2], addr_581_5, wires_2326_6,addr_2326_6);

wire[3:0] wires_2327_6;

wire[31:0] addr_2327_6;

Selector_2 s2327_6(wires_581_5[3], addr_581_5, wires_2327_6,addr_2327_6);

wire[3:0] wires_2328_6;

wire[31:0] addr_2328_6;

Selector_2 s2328_6(wires_582_5[0], addr_582_5, wires_2328_6,addr_2328_6);

wire[3:0] wires_2329_6;

wire[31:0] addr_2329_6;

Selector_2 s2329_6(wires_582_5[1], addr_582_5, wires_2329_6,addr_2329_6);

wire[3:0] wires_2330_6;

wire[31:0] addr_2330_6;

Selector_2 s2330_6(wires_582_5[2], addr_582_5, wires_2330_6,addr_2330_6);

wire[3:0] wires_2331_6;

wire[31:0] addr_2331_6;

Selector_2 s2331_6(wires_582_5[3], addr_582_5, wires_2331_6,addr_2331_6);

wire[3:0] wires_2332_6;

wire[31:0] addr_2332_6;

Selector_2 s2332_6(wires_583_5[0], addr_583_5, wires_2332_6,addr_2332_6);

wire[3:0] wires_2333_6;

wire[31:0] addr_2333_6;

Selector_2 s2333_6(wires_583_5[1], addr_583_5, wires_2333_6,addr_2333_6);

wire[3:0] wires_2334_6;

wire[31:0] addr_2334_6;

Selector_2 s2334_6(wires_583_5[2], addr_583_5, wires_2334_6,addr_2334_6);

wire[3:0] wires_2335_6;

wire[31:0] addr_2335_6;

Selector_2 s2335_6(wires_583_5[3], addr_583_5, wires_2335_6,addr_2335_6);

wire[3:0] wires_2336_6;

wire[31:0] addr_2336_6;

Selector_2 s2336_6(wires_584_5[0], addr_584_5, wires_2336_6,addr_2336_6);

wire[3:0] wires_2337_6;

wire[31:0] addr_2337_6;

Selector_2 s2337_6(wires_584_5[1], addr_584_5, wires_2337_6,addr_2337_6);

wire[3:0] wires_2338_6;

wire[31:0] addr_2338_6;

Selector_2 s2338_6(wires_584_5[2], addr_584_5, wires_2338_6,addr_2338_6);

wire[3:0] wires_2339_6;

wire[31:0] addr_2339_6;

Selector_2 s2339_6(wires_584_5[3], addr_584_5, wires_2339_6,addr_2339_6);

wire[3:0] wires_2340_6;

wire[31:0] addr_2340_6;

Selector_2 s2340_6(wires_585_5[0], addr_585_5, wires_2340_6,addr_2340_6);

wire[3:0] wires_2341_6;

wire[31:0] addr_2341_6;

Selector_2 s2341_6(wires_585_5[1], addr_585_5, wires_2341_6,addr_2341_6);

wire[3:0] wires_2342_6;

wire[31:0] addr_2342_6;

Selector_2 s2342_6(wires_585_5[2], addr_585_5, wires_2342_6,addr_2342_6);

wire[3:0] wires_2343_6;

wire[31:0] addr_2343_6;

Selector_2 s2343_6(wires_585_5[3], addr_585_5, wires_2343_6,addr_2343_6);

wire[3:0] wires_2344_6;

wire[31:0] addr_2344_6;

Selector_2 s2344_6(wires_586_5[0], addr_586_5, wires_2344_6,addr_2344_6);

wire[3:0] wires_2345_6;

wire[31:0] addr_2345_6;

Selector_2 s2345_6(wires_586_5[1], addr_586_5, wires_2345_6,addr_2345_6);

wire[3:0] wires_2346_6;

wire[31:0] addr_2346_6;

Selector_2 s2346_6(wires_586_5[2], addr_586_5, wires_2346_6,addr_2346_6);

wire[3:0] wires_2347_6;

wire[31:0] addr_2347_6;

Selector_2 s2347_6(wires_586_5[3], addr_586_5, wires_2347_6,addr_2347_6);

wire[3:0] wires_2348_6;

wire[31:0] addr_2348_6;

Selector_2 s2348_6(wires_587_5[0], addr_587_5, wires_2348_6,addr_2348_6);

wire[3:0] wires_2349_6;

wire[31:0] addr_2349_6;

Selector_2 s2349_6(wires_587_5[1], addr_587_5, wires_2349_6,addr_2349_6);

wire[3:0] wires_2350_6;

wire[31:0] addr_2350_6;

Selector_2 s2350_6(wires_587_5[2], addr_587_5, wires_2350_6,addr_2350_6);

wire[3:0] wires_2351_6;

wire[31:0] addr_2351_6;

Selector_2 s2351_6(wires_587_5[3], addr_587_5, wires_2351_6,addr_2351_6);

wire[3:0] wires_2352_6;

wire[31:0] addr_2352_6;

Selector_2 s2352_6(wires_588_5[0], addr_588_5, wires_2352_6,addr_2352_6);

wire[3:0] wires_2353_6;

wire[31:0] addr_2353_6;

Selector_2 s2353_6(wires_588_5[1], addr_588_5, wires_2353_6,addr_2353_6);

wire[3:0] wires_2354_6;

wire[31:0] addr_2354_6;

Selector_2 s2354_6(wires_588_5[2], addr_588_5, wires_2354_6,addr_2354_6);

wire[3:0] wires_2355_6;

wire[31:0] addr_2355_6;

Selector_2 s2355_6(wires_588_5[3], addr_588_5, wires_2355_6,addr_2355_6);

wire[3:0] wires_2356_6;

wire[31:0] addr_2356_6;

Selector_2 s2356_6(wires_589_5[0], addr_589_5, wires_2356_6,addr_2356_6);

wire[3:0] wires_2357_6;

wire[31:0] addr_2357_6;

Selector_2 s2357_6(wires_589_5[1], addr_589_5, wires_2357_6,addr_2357_6);

wire[3:0] wires_2358_6;

wire[31:0] addr_2358_6;

Selector_2 s2358_6(wires_589_5[2], addr_589_5, wires_2358_6,addr_2358_6);

wire[3:0] wires_2359_6;

wire[31:0] addr_2359_6;

Selector_2 s2359_6(wires_589_5[3], addr_589_5, wires_2359_6,addr_2359_6);

wire[3:0] wires_2360_6;

wire[31:0] addr_2360_6;

Selector_2 s2360_6(wires_590_5[0], addr_590_5, wires_2360_6,addr_2360_6);

wire[3:0] wires_2361_6;

wire[31:0] addr_2361_6;

Selector_2 s2361_6(wires_590_5[1], addr_590_5, wires_2361_6,addr_2361_6);

wire[3:0] wires_2362_6;

wire[31:0] addr_2362_6;

Selector_2 s2362_6(wires_590_5[2], addr_590_5, wires_2362_6,addr_2362_6);

wire[3:0] wires_2363_6;

wire[31:0] addr_2363_6;

Selector_2 s2363_6(wires_590_5[3], addr_590_5, wires_2363_6,addr_2363_6);

wire[3:0] wires_2364_6;

wire[31:0] addr_2364_6;

Selector_2 s2364_6(wires_591_5[0], addr_591_5, wires_2364_6,addr_2364_6);

wire[3:0] wires_2365_6;

wire[31:0] addr_2365_6;

Selector_2 s2365_6(wires_591_5[1], addr_591_5, wires_2365_6,addr_2365_6);

wire[3:0] wires_2366_6;

wire[31:0] addr_2366_6;

Selector_2 s2366_6(wires_591_5[2], addr_591_5, wires_2366_6,addr_2366_6);

wire[3:0] wires_2367_6;

wire[31:0] addr_2367_6;

Selector_2 s2367_6(wires_591_5[3], addr_591_5, wires_2367_6,addr_2367_6);

wire[3:0] wires_2368_6;

wire[31:0] addr_2368_6;

Selector_2 s2368_6(wires_592_5[0], addr_592_5, wires_2368_6,addr_2368_6);

wire[3:0] wires_2369_6;

wire[31:0] addr_2369_6;

Selector_2 s2369_6(wires_592_5[1], addr_592_5, wires_2369_6,addr_2369_6);

wire[3:0] wires_2370_6;

wire[31:0] addr_2370_6;

Selector_2 s2370_6(wires_592_5[2], addr_592_5, wires_2370_6,addr_2370_6);

wire[3:0] wires_2371_6;

wire[31:0] addr_2371_6;

Selector_2 s2371_6(wires_592_5[3], addr_592_5, wires_2371_6,addr_2371_6);

wire[3:0] wires_2372_6;

wire[31:0] addr_2372_6;

Selector_2 s2372_6(wires_593_5[0], addr_593_5, wires_2372_6,addr_2372_6);

wire[3:0] wires_2373_6;

wire[31:0] addr_2373_6;

Selector_2 s2373_6(wires_593_5[1], addr_593_5, wires_2373_6,addr_2373_6);

wire[3:0] wires_2374_6;

wire[31:0] addr_2374_6;

Selector_2 s2374_6(wires_593_5[2], addr_593_5, wires_2374_6,addr_2374_6);

wire[3:0] wires_2375_6;

wire[31:0] addr_2375_6;

Selector_2 s2375_6(wires_593_5[3], addr_593_5, wires_2375_6,addr_2375_6);

wire[3:0] wires_2376_6;

wire[31:0] addr_2376_6;

Selector_2 s2376_6(wires_594_5[0], addr_594_5, wires_2376_6,addr_2376_6);

wire[3:0] wires_2377_6;

wire[31:0] addr_2377_6;

Selector_2 s2377_6(wires_594_5[1], addr_594_5, wires_2377_6,addr_2377_6);

wire[3:0] wires_2378_6;

wire[31:0] addr_2378_6;

Selector_2 s2378_6(wires_594_5[2], addr_594_5, wires_2378_6,addr_2378_6);

wire[3:0] wires_2379_6;

wire[31:0] addr_2379_6;

Selector_2 s2379_6(wires_594_5[3], addr_594_5, wires_2379_6,addr_2379_6);

wire[3:0] wires_2380_6;

wire[31:0] addr_2380_6;

Selector_2 s2380_6(wires_595_5[0], addr_595_5, wires_2380_6,addr_2380_6);

wire[3:0] wires_2381_6;

wire[31:0] addr_2381_6;

Selector_2 s2381_6(wires_595_5[1], addr_595_5, wires_2381_6,addr_2381_6);

wire[3:0] wires_2382_6;

wire[31:0] addr_2382_6;

Selector_2 s2382_6(wires_595_5[2], addr_595_5, wires_2382_6,addr_2382_6);

wire[3:0] wires_2383_6;

wire[31:0] addr_2383_6;

Selector_2 s2383_6(wires_595_5[3], addr_595_5, wires_2383_6,addr_2383_6);

wire[3:0] wires_2384_6;

wire[31:0] addr_2384_6;

Selector_2 s2384_6(wires_596_5[0], addr_596_5, wires_2384_6,addr_2384_6);

wire[3:0] wires_2385_6;

wire[31:0] addr_2385_6;

Selector_2 s2385_6(wires_596_5[1], addr_596_5, wires_2385_6,addr_2385_6);

wire[3:0] wires_2386_6;

wire[31:0] addr_2386_6;

Selector_2 s2386_6(wires_596_5[2], addr_596_5, wires_2386_6,addr_2386_6);

wire[3:0] wires_2387_6;

wire[31:0] addr_2387_6;

Selector_2 s2387_6(wires_596_5[3], addr_596_5, wires_2387_6,addr_2387_6);

wire[3:0] wires_2388_6;

wire[31:0] addr_2388_6;

Selector_2 s2388_6(wires_597_5[0], addr_597_5, wires_2388_6,addr_2388_6);

wire[3:0] wires_2389_6;

wire[31:0] addr_2389_6;

Selector_2 s2389_6(wires_597_5[1], addr_597_5, wires_2389_6,addr_2389_6);

wire[3:0] wires_2390_6;

wire[31:0] addr_2390_6;

Selector_2 s2390_6(wires_597_5[2], addr_597_5, wires_2390_6,addr_2390_6);

wire[3:0] wires_2391_6;

wire[31:0] addr_2391_6;

Selector_2 s2391_6(wires_597_5[3], addr_597_5, wires_2391_6,addr_2391_6);

wire[3:0] wires_2392_6;

wire[31:0] addr_2392_6;

Selector_2 s2392_6(wires_598_5[0], addr_598_5, wires_2392_6,addr_2392_6);

wire[3:0] wires_2393_6;

wire[31:0] addr_2393_6;

Selector_2 s2393_6(wires_598_5[1], addr_598_5, wires_2393_6,addr_2393_6);

wire[3:0] wires_2394_6;

wire[31:0] addr_2394_6;

Selector_2 s2394_6(wires_598_5[2], addr_598_5, wires_2394_6,addr_2394_6);

wire[3:0] wires_2395_6;

wire[31:0] addr_2395_6;

Selector_2 s2395_6(wires_598_5[3], addr_598_5, wires_2395_6,addr_2395_6);

wire[3:0] wires_2396_6;

wire[31:0] addr_2396_6;

Selector_2 s2396_6(wires_599_5[0], addr_599_5, wires_2396_6,addr_2396_6);

wire[3:0] wires_2397_6;

wire[31:0] addr_2397_6;

Selector_2 s2397_6(wires_599_5[1], addr_599_5, wires_2397_6,addr_2397_6);

wire[3:0] wires_2398_6;

wire[31:0] addr_2398_6;

Selector_2 s2398_6(wires_599_5[2], addr_599_5, wires_2398_6,addr_2398_6);

wire[3:0] wires_2399_6;

wire[31:0] addr_2399_6;

Selector_2 s2399_6(wires_599_5[3], addr_599_5, wires_2399_6,addr_2399_6);

wire[3:0] wires_2400_6;

wire[31:0] addr_2400_6;

Selector_2 s2400_6(wires_600_5[0], addr_600_5, wires_2400_6,addr_2400_6);

wire[3:0] wires_2401_6;

wire[31:0] addr_2401_6;

Selector_2 s2401_6(wires_600_5[1], addr_600_5, wires_2401_6,addr_2401_6);

wire[3:0] wires_2402_6;

wire[31:0] addr_2402_6;

Selector_2 s2402_6(wires_600_5[2], addr_600_5, wires_2402_6,addr_2402_6);

wire[3:0] wires_2403_6;

wire[31:0] addr_2403_6;

Selector_2 s2403_6(wires_600_5[3], addr_600_5, wires_2403_6,addr_2403_6);

wire[3:0] wires_2404_6;

wire[31:0] addr_2404_6;

Selector_2 s2404_6(wires_601_5[0], addr_601_5, wires_2404_6,addr_2404_6);

wire[3:0] wires_2405_6;

wire[31:0] addr_2405_6;

Selector_2 s2405_6(wires_601_5[1], addr_601_5, wires_2405_6,addr_2405_6);

wire[3:0] wires_2406_6;

wire[31:0] addr_2406_6;

Selector_2 s2406_6(wires_601_5[2], addr_601_5, wires_2406_6,addr_2406_6);

wire[3:0] wires_2407_6;

wire[31:0] addr_2407_6;

Selector_2 s2407_6(wires_601_5[3], addr_601_5, wires_2407_6,addr_2407_6);

wire[3:0] wires_2408_6;

wire[31:0] addr_2408_6;

Selector_2 s2408_6(wires_602_5[0], addr_602_5, wires_2408_6,addr_2408_6);

wire[3:0] wires_2409_6;

wire[31:0] addr_2409_6;

Selector_2 s2409_6(wires_602_5[1], addr_602_5, wires_2409_6,addr_2409_6);

wire[3:0] wires_2410_6;

wire[31:0] addr_2410_6;

Selector_2 s2410_6(wires_602_5[2], addr_602_5, wires_2410_6,addr_2410_6);

wire[3:0] wires_2411_6;

wire[31:0] addr_2411_6;

Selector_2 s2411_6(wires_602_5[3], addr_602_5, wires_2411_6,addr_2411_6);

wire[3:0] wires_2412_6;

wire[31:0] addr_2412_6;

Selector_2 s2412_6(wires_603_5[0], addr_603_5, wires_2412_6,addr_2412_6);

wire[3:0] wires_2413_6;

wire[31:0] addr_2413_6;

Selector_2 s2413_6(wires_603_5[1], addr_603_5, wires_2413_6,addr_2413_6);

wire[3:0] wires_2414_6;

wire[31:0] addr_2414_6;

Selector_2 s2414_6(wires_603_5[2], addr_603_5, wires_2414_6,addr_2414_6);

wire[3:0] wires_2415_6;

wire[31:0] addr_2415_6;

Selector_2 s2415_6(wires_603_5[3], addr_603_5, wires_2415_6,addr_2415_6);

wire[3:0] wires_2416_6;

wire[31:0] addr_2416_6;

Selector_2 s2416_6(wires_604_5[0], addr_604_5, wires_2416_6,addr_2416_6);

wire[3:0] wires_2417_6;

wire[31:0] addr_2417_6;

Selector_2 s2417_6(wires_604_5[1], addr_604_5, wires_2417_6,addr_2417_6);

wire[3:0] wires_2418_6;

wire[31:0] addr_2418_6;

Selector_2 s2418_6(wires_604_5[2], addr_604_5, wires_2418_6,addr_2418_6);

wire[3:0] wires_2419_6;

wire[31:0] addr_2419_6;

Selector_2 s2419_6(wires_604_5[3], addr_604_5, wires_2419_6,addr_2419_6);

wire[3:0] wires_2420_6;

wire[31:0] addr_2420_6;

Selector_2 s2420_6(wires_605_5[0], addr_605_5, wires_2420_6,addr_2420_6);

wire[3:0] wires_2421_6;

wire[31:0] addr_2421_6;

Selector_2 s2421_6(wires_605_5[1], addr_605_5, wires_2421_6,addr_2421_6);

wire[3:0] wires_2422_6;

wire[31:0] addr_2422_6;

Selector_2 s2422_6(wires_605_5[2], addr_605_5, wires_2422_6,addr_2422_6);

wire[3:0] wires_2423_6;

wire[31:0] addr_2423_6;

Selector_2 s2423_6(wires_605_5[3], addr_605_5, wires_2423_6,addr_2423_6);

wire[3:0] wires_2424_6;

wire[31:0] addr_2424_6;

Selector_2 s2424_6(wires_606_5[0], addr_606_5, wires_2424_6,addr_2424_6);

wire[3:0] wires_2425_6;

wire[31:0] addr_2425_6;

Selector_2 s2425_6(wires_606_5[1], addr_606_5, wires_2425_6,addr_2425_6);

wire[3:0] wires_2426_6;

wire[31:0] addr_2426_6;

Selector_2 s2426_6(wires_606_5[2], addr_606_5, wires_2426_6,addr_2426_6);

wire[3:0] wires_2427_6;

wire[31:0] addr_2427_6;

Selector_2 s2427_6(wires_606_5[3], addr_606_5, wires_2427_6,addr_2427_6);

wire[3:0] wires_2428_6;

wire[31:0] addr_2428_6;

Selector_2 s2428_6(wires_607_5[0], addr_607_5, wires_2428_6,addr_2428_6);

wire[3:0] wires_2429_6;

wire[31:0] addr_2429_6;

Selector_2 s2429_6(wires_607_5[1], addr_607_5, wires_2429_6,addr_2429_6);

wire[3:0] wires_2430_6;

wire[31:0] addr_2430_6;

Selector_2 s2430_6(wires_607_5[2], addr_607_5, wires_2430_6,addr_2430_6);

wire[3:0] wires_2431_6;

wire[31:0] addr_2431_6;

Selector_2 s2431_6(wires_607_5[3], addr_607_5, wires_2431_6,addr_2431_6);

wire[3:0] wires_2432_6;

wire[31:0] addr_2432_6;

Selector_2 s2432_6(wires_608_5[0], addr_608_5, wires_2432_6,addr_2432_6);

wire[3:0] wires_2433_6;

wire[31:0] addr_2433_6;

Selector_2 s2433_6(wires_608_5[1], addr_608_5, wires_2433_6,addr_2433_6);

wire[3:0] wires_2434_6;

wire[31:0] addr_2434_6;

Selector_2 s2434_6(wires_608_5[2], addr_608_5, wires_2434_6,addr_2434_6);

wire[3:0] wires_2435_6;

wire[31:0] addr_2435_6;

Selector_2 s2435_6(wires_608_5[3], addr_608_5, wires_2435_6,addr_2435_6);

wire[3:0] wires_2436_6;

wire[31:0] addr_2436_6;

Selector_2 s2436_6(wires_609_5[0], addr_609_5, wires_2436_6,addr_2436_6);

wire[3:0] wires_2437_6;

wire[31:0] addr_2437_6;

Selector_2 s2437_6(wires_609_5[1], addr_609_5, wires_2437_6,addr_2437_6);

wire[3:0] wires_2438_6;

wire[31:0] addr_2438_6;

Selector_2 s2438_6(wires_609_5[2], addr_609_5, wires_2438_6,addr_2438_6);

wire[3:0] wires_2439_6;

wire[31:0] addr_2439_6;

Selector_2 s2439_6(wires_609_5[3], addr_609_5, wires_2439_6,addr_2439_6);

wire[3:0] wires_2440_6;

wire[31:0] addr_2440_6;

Selector_2 s2440_6(wires_610_5[0], addr_610_5, wires_2440_6,addr_2440_6);

wire[3:0] wires_2441_6;

wire[31:0] addr_2441_6;

Selector_2 s2441_6(wires_610_5[1], addr_610_5, wires_2441_6,addr_2441_6);

wire[3:0] wires_2442_6;

wire[31:0] addr_2442_6;

Selector_2 s2442_6(wires_610_5[2], addr_610_5, wires_2442_6,addr_2442_6);

wire[3:0] wires_2443_6;

wire[31:0] addr_2443_6;

Selector_2 s2443_6(wires_610_5[3], addr_610_5, wires_2443_6,addr_2443_6);

wire[3:0] wires_2444_6;

wire[31:0] addr_2444_6;

Selector_2 s2444_6(wires_611_5[0], addr_611_5, wires_2444_6,addr_2444_6);

wire[3:0] wires_2445_6;

wire[31:0] addr_2445_6;

Selector_2 s2445_6(wires_611_5[1], addr_611_5, wires_2445_6,addr_2445_6);

wire[3:0] wires_2446_6;

wire[31:0] addr_2446_6;

Selector_2 s2446_6(wires_611_5[2], addr_611_5, wires_2446_6,addr_2446_6);

wire[3:0] wires_2447_6;

wire[31:0] addr_2447_6;

Selector_2 s2447_6(wires_611_5[3], addr_611_5, wires_2447_6,addr_2447_6);

wire[3:0] wires_2448_6;

wire[31:0] addr_2448_6;

Selector_2 s2448_6(wires_612_5[0], addr_612_5, wires_2448_6,addr_2448_6);

wire[3:0] wires_2449_6;

wire[31:0] addr_2449_6;

Selector_2 s2449_6(wires_612_5[1], addr_612_5, wires_2449_6,addr_2449_6);

wire[3:0] wires_2450_6;

wire[31:0] addr_2450_6;

Selector_2 s2450_6(wires_612_5[2], addr_612_5, wires_2450_6,addr_2450_6);

wire[3:0] wires_2451_6;

wire[31:0] addr_2451_6;

Selector_2 s2451_6(wires_612_5[3], addr_612_5, wires_2451_6,addr_2451_6);

wire[3:0] wires_2452_6;

wire[31:0] addr_2452_6;

Selector_2 s2452_6(wires_613_5[0], addr_613_5, wires_2452_6,addr_2452_6);

wire[3:0] wires_2453_6;

wire[31:0] addr_2453_6;

Selector_2 s2453_6(wires_613_5[1], addr_613_5, wires_2453_6,addr_2453_6);

wire[3:0] wires_2454_6;

wire[31:0] addr_2454_6;

Selector_2 s2454_6(wires_613_5[2], addr_613_5, wires_2454_6,addr_2454_6);

wire[3:0] wires_2455_6;

wire[31:0] addr_2455_6;

Selector_2 s2455_6(wires_613_5[3], addr_613_5, wires_2455_6,addr_2455_6);

wire[3:0] wires_2456_6;

wire[31:0] addr_2456_6;

Selector_2 s2456_6(wires_614_5[0], addr_614_5, wires_2456_6,addr_2456_6);

wire[3:0] wires_2457_6;

wire[31:0] addr_2457_6;

Selector_2 s2457_6(wires_614_5[1], addr_614_5, wires_2457_6,addr_2457_6);

wire[3:0] wires_2458_6;

wire[31:0] addr_2458_6;

Selector_2 s2458_6(wires_614_5[2], addr_614_5, wires_2458_6,addr_2458_6);

wire[3:0] wires_2459_6;

wire[31:0] addr_2459_6;

Selector_2 s2459_6(wires_614_5[3], addr_614_5, wires_2459_6,addr_2459_6);

wire[3:0] wires_2460_6;

wire[31:0] addr_2460_6;

Selector_2 s2460_6(wires_615_5[0], addr_615_5, wires_2460_6,addr_2460_6);

wire[3:0] wires_2461_6;

wire[31:0] addr_2461_6;

Selector_2 s2461_6(wires_615_5[1], addr_615_5, wires_2461_6,addr_2461_6);

wire[3:0] wires_2462_6;

wire[31:0] addr_2462_6;

Selector_2 s2462_6(wires_615_5[2], addr_615_5, wires_2462_6,addr_2462_6);

wire[3:0] wires_2463_6;

wire[31:0] addr_2463_6;

Selector_2 s2463_6(wires_615_5[3], addr_615_5, wires_2463_6,addr_2463_6);

wire[3:0] wires_2464_6;

wire[31:0] addr_2464_6;

Selector_2 s2464_6(wires_616_5[0], addr_616_5, wires_2464_6,addr_2464_6);

wire[3:0] wires_2465_6;

wire[31:0] addr_2465_6;

Selector_2 s2465_6(wires_616_5[1], addr_616_5, wires_2465_6,addr_2465_6);

wire[3:0] wires_2466_6;

wire[31:0] addr_2466_6;

Selector_2 s2466_6(wires_616_5[2], addr_616_5, wires_2466_6,addr_2466_6);

wire[3:0] wires_2467_6;

wire[31:0] addr_2467_6;

Selector_2 s2467_6(wires_616_5[3], addr_616_5, wires_2467_6,addr_2467_6);

wire[3:0] wires_2468_6;

wire[31:0] addr_2468_6;

Selector_2 s2468_6(wires_617_5[0], addr_617_5, wires_2468_6,addr_2468_6);

wire[3:0] wires_2469_6;

wire[31:0] addr_2469_6;

Selector_2 s2469_6(wires_617_5[1], addr_617_5, wires_2469_6,addr_2469_6);

wire[3:0] wires_2470_6;

wire[31:0] addr_2470_6;

Selector_2 s2470_6(wires_617_5[2], addr_617_5, wires_2470_6,addr_2470_6);

wire[3:0] wires_2471_6;

wire[31:0] addr_2471_6;

Selector_2 s2471_6(wires_617_5[3], addr_617_5, wires_2471_6,addr_2471_6);

wire[3:0] wires_2472_6;

wire[31:0] addr_2472_6;

Selector_2 s2472_6(wires_618_5[0], addr_618_5, wires_2472_6,addr_2472_6);

wire[3:0] wires_2473_6;

wire[31:0] addr_2473_6;

Selector_2 s2473_6(wires_618_5[1], addr_618_5, wires_2473_6,addr_2473_6);

wire[3:0] wires_2474_6;

wire[31:0] addr_2474_6;

Selector_2 s2474_6(wires_618_5[2], addr_618_5, wires_2474_6,addr_2474_6);

wire[3:0] wires_2475_6;

wire[31:0] addr_2475_6;

Selector_2 s2475_6(wires_618_5[3], addr_618_5, wires_2475_6,addr_2475_6);

wire[3:0] wires_2476_6;

wire[31:0] addr_2476_6;

Selector_2 s2476_6(wires_619_5[0], addr_619_5, wires_2476_6,addr_2476_6);

wire[3:0] wires_2477_6;

wire[31:0] addr_2477_6;

Selector_2 s2477_6(wires_619_5[1], addr_619_5, wires_2477_6,addr_2477_6);

wire[3:0] wires_2478_6;

wire[31:0] addr_2478_6;

Selector_2 s2478_6(wires_619_5[2], addr_619_5, wires_2478_6,addr_2478_6);

wire[3:0] wires_2479_6;

wire[31:0] addr_2479_6;

Selector_2 s2479_6(wires_619_5[3], addr_619_5, wires_2479_6,addr_2479_6);

wire[3:0] wires_2480_6;

wire[31:0] addr_2480_6;

Selector_2 s2480_6(wires_620_5[0], addr_620_5, wires_2480_6,addr_2480_6);

wire[3:0] wires_2481_6;

wire[31:0] addr_2481_6;

Selector_2 s2481_6(wires_620_5[1], addr_620_5, wires_2481_6,addr_2481_6);

wire[3:0] wires_2482_6;

wire[31:0] addr_2482_6;

Selector_2 s2482_6(wires_620_5[2], addr_620_5, wires_2482_6,addr_2482_6);

wire[3:0] wires_2483_6;

wire[31:0] addr_2483_6;

Selector_2 s2483_6(wires_620_5[3], addr_620_5, wires_2483_6,addr_2483_6);

wire[3:0] wires_2484_6;

wire[31:0] addr_2484_6;

Selector_2 s2484_6(wires_621_5[0], addr_621_5, wires_2484_6,addr_2484_6);

wire[3:0] wires_2485_6;

wire[31:0] addr_2485_6;

Selector_2 s2485_6(wires_621_5[1], addr_621_5, wires_2485_6,addr_2485_6);

wire[3:0] wires_2486_6;

wire[31:0] addr_2486_6;

Selector_2 s2486_6(wires_621_5[2], addr_621_5, wires_2486_6,addr_2486_6);

wire[3:0] wires_2487_6;

wire[31:0] addr_2487_6;

Selector_2 s2487_6(wires_621_5[3], addr_621_5, wires_2487_6,addr_2487_6);

wire[3:0] wires_2488_6;

wire[31:0] addr_2488_6;

Selector_2 s2488_6(wires_622_5[0], addr_622_5, wires_2488_6,addr_2488_6);

wire[3:0] wires_2489_6;

wire[31:0] addr_2489_6;

Selector_2 s2489_6(wires_622_5[1], addr_622_5, wires_2489_6,addr_2489_6);

wire[3:0] wires_2490_6;

wire[31:0] addr_2490_6;

Selector_2 s2490_6(wires_622_5[2], addr_622_5, wires_2490_6,addr_2490_6);

wire[3:0] wires_2491_6;

wire[31:0] addr_2491_6;

Selector_2 s2491_6(wires_622_5[3], addr_622_5, wires_2491_6,addr_2491_6);

wire[3:0] wires_2492_6;

wire[31:0] addr_2492_6;

Selector_2 s2492_6(wires_623_5[0], addr_623_5, wires_2492_6,addr_2492_6);

wire[3:0] wires_2493_6;

wire[31:0] addr_2493_6;

Selector_2 s2493_6(wires_623_5[1], addr_623_5, wires_2493_6,addr_2493_6);

wire[3:0] wires_2494_6;

wire[31:0] addr_2494_6;

Selector_2 s2494_6(wires_623_5[2], addr_623_5, wires_2494_6,addr_2494_6);

wire[3:0] wires_2495_6;

wire[31:0] addr_2495_6;

Selector_2 s2495_6(wires_623_5[3], addr_623_5, wires_2495_6,addr_2495_6);

wire[3:0] wires_2496_6;

wire[31:0] addr_2496_6;

Selector_2 s2496_6(wires_624_5[0], addr_624_5, wires_2496_6,addr_2496_6);

wire[3:0] wires_2497_6;

wire[31:0] addr_2497_6;

Selector_2 s2497_6(wires_624_5[1], addr_624_5, wires_2497_6,addr_2497_6);

wire[3:0] wires_2498_6;

wire[31:0] addr_2498_6;

Selector_2 s2498_6(wires_624_5[2], addr_624_5, wires_2498_6,addr_2498_6);

wire[3:0] wires_2499_6;

wire[31:0] addr_2499_6;

Selector_2 s2499_6(wires_624_5[3], addr_624_5, wires_2499_6,addr_2499_6);

wire[3:0] wires_2500_6;

wire[31:0] addr_2500_6;

Selector_2 s2500_6(wires_625_5[0], addr_625_5, wires_2500_6,addr_2500_6);

wire[3:0] wires_2501_6;

wire[31:0] addr_2501_6;

Selector_2 s2501_6(wires_625_5[1], addr_625_5, wires_2501_6,addr_2501_6);

wire[3:0] wires_2502_6;

wire[31:0] addr_2502_6;

Selector_2 s2502_6(wires_625_5[2], addr_625_5, wires_2502_6,addr_2502_6);

wire[3:0] wires_2503_6;

wire[31:0] addr_2503_6;

Selector_2 s2503_6(wires_625_5[3], addr_625_5, wires_2503_6,addr_2503_6);

wire[3:0] wires_2504_6;

wire[31:0] addr_2504_6;

Selector_2 s2504_6(wires_626_5[0], addr_626_5, wires_2504_6,addr_2504_6);

wire[3:0] wires_2505_6;

wire[31:0] addr_2505_6;

Selector_2 s2505_6(wires_626_5[1], addr_626_5, wires_2505_6,addr_2505_6);

wire[3:0] wires_2506_6;

wire[31:0] addr_2506_6;

Selector_2 s2506_6(wires_626_5[2], addr_626_5, wires_2506_6,addr_2506_6);

wire[3:0] wires_2507_6;

wire[31:0] addr_2507_6;

Selector_2 s2507_6(wires_626_5[3], addr_626_5, wires_2507_6,addr_2507_6);

wire[3:0] wires_2508_6;

wire[31:0] addr_2508_6;

Selector_2 s2508_6(wires_627_5[0], addr_627_5, wires_2508_6,addr_2508_6);

wire[3:0] wires_2509_6;

wire[31:0] addr_2509_6;

Selector_2 s2509_6(wires_627_5[1], addr_627_5, wires_2509_6,addr_2509_6);

wire[3:0] wires_2510_6;

wire[31:0] addr_2510_6;

Selector_2 s2510_6(wires_627_5[2], addr_627_5, wires_2510_6,addr_2510_6);

wire[3:0] wires_2511_6;

wire[31:0] addr_2511_6;

Selector_2 s2511_6(wires_627_5[3], addr_627_5, wires_2511_6,addr_2511_6);

wire[3:0] wires_2512_6;

wire[31:0] addr_2512_6;

Selector_2 s2512_6(wires_628_5[0], addr_628_5, wires_2512_6,addr_2512_6);

wire[3:0] wires_2513_6;

wire[31:0] addr_2513_6;

Selector_2 s2513_6(wires_628_5[1], addr_628_5, wires_2513_6,addr_2513_6);

wire[3:0] wires_2514_6;

wire[31:0] addr_2514_6;

Selector_2 s2514_6(wires_628_5[2], addr_628_5, wires_2514_6,addr_2514_6);

wire[3:0] wires_2515_6;

wire[31:0] addr_2515_6;

Selector_2 s2515_6(wires_628_5[3], addr_628_5, wires_2515_6,addr_2515_6);

wire[3:0] wires_2516_6;

wire[31:0] addr_2516_6;

Selector_2 s2516_6(wires_629_5[0], addr_629_5, wires_2516_6,addr_2516_6);

wire[3:0] wires_2517_6;

wire[31:0] addr_2517_6;

Selector_2 s2517_6(wires_629_5[1], addr_629_5, wires_2517_6,addr_2517_6);

wire[3:0] wires_2518_6;

wire[31:0] addr_2518_6;

Selector_2 s2518_6(wires_629_5[2], addr_629_5, wires_2518_6,addr_2518_6);

wire[3:0] wires_2519_6;

wire[31:0] addr_2519_6;

Selector_2 s2519_6(wires_629_5[3], addr_629_5, wires_2519_6,addr_2519_6);

wire[3:0] wires_2520_6;

wire[31:0] addr_2520_6;

Selector_2 s2520_6(wires_630_5[0], addr_630_5, wires_2520_6,addr_2520_6);

wire[3:0] wires_2521_6;

wire[31:0] addr_2521_6;

Selector_2 s2521_6(wires_630_5[1], addr_630_5, wires_2521_6,addr_2521_6);

wire[3:0] wires_2522_6;

wire[31:0] addr_2522_6;

Selector_2 s2522_6(wires_630_5[2], addr_630_5, wires_2522_6,addr_2522_6);

wire[3:0] wires_2523_6;

wire[31:0] addr_2523_6;

Selector_2 s2523_6(wires_630_5[3], addr_630_5, wires_2523_6,addr_2523_6);

wire[3:0] wires_2524_6;

wire[31:0] addr_2524_6;

Selector_2 s2524_6(wires_631_5[0], addr_631_5, wires_2524_6,addr_2524_6);

wire[3:0] wires_2525_6;

wire[31:0] addr_2525_6;

Selector_2 s2525_6(wires_631_5[1], addr_631_5, wires_2525_6,addr_2525_6);

wire[3:0] wires_2526_6;

wire[31:0] addr_2526_6;

Selector_2 s2526_6(wires_631_5[2], addr_631_5, wires_2526_6,addr_2526_6);

wire[3:0] wires_2527_6;

wire[31:0] addr_2527_6;

Selector_2 s2527_6(wires_631_5[3], addr_631_5, wires_2527_6,addr_2527_6);

wire[3:0] wires_2528_6;

wire[31:0] addr_2528_6;

Selector_2 s2528_6(wires_632_5[0], addr_632_5, wires_2528_6,addr_2528_6);

wire[3:0] wires_2529_6;

wire[31:0] addr_2529_6;

Selector_2 s2529_6(wires_632_5[1], addr_632_5, wires_2529_6,addr_2529_6);

wire[3:0] wires_2530_6;

wire[31:0] addr_2530_6;

Selector_2 s2530_6(wires_632_5[2], addr_632_5, wires_2530_6,addr_2530_6);

wire[3:0] wires_2531_6;

wire[31:0] addr_2531_6;

Selector_2 s2531_6(wires_632_5[3], addr_632_5, wires_2531_6,addr_2531_6);

wire[3:0] wires_2532_6;

wire[31:0] addr_2532_6;

Selector_2 s2532_6(wires_633_5[0], addr_633_5, wires_2532_6,addr_2532_6);

wire[3:0] wires_2533_6;

wire[31:0] addr_2533_6;

Selector_2 s2533_6(wires_633_5[1], addr_633_5, wires_2533_6,addr_2533_6);

wire[3:0] wires_2534_6;

wire[31:0] addr_2534_6;

Selector_2 s2534_6(wires_633_5[2], addr_633_5, wires_2534_6,addr_2534_6);

wire[3:0] wires_2535_6;

wire[31:0] addr_2535_6;

Selector_2 s2535_6(wires_633_5[3], addr_633_5, wires_2535_6,addr_2535_6);

wire[3:0] wires_2536_6;

wire[31:0] addr_2536_6;

Selector_2 s2536_6(wires_634_5[0], addr_634_5, wires_2536_6,addr_2536_6);

wire[3:0] wires_2537_6;

wire[31:0] addr_2537_6;

Selector_2 s2537_6(wires_634_5[1], addr_634_5, wires_2537_6,addr_2537_6);

wire[3:0] wires_2538_6;

wire[31:0] addr_2538_6;

Selector_2 s2538_6(wires_634_5[2], addr_634_5, wires_2538_6,addr_2538_6);

wire[3:0] wires_2539_6;

wire[31:0] addr_2539_6;

Selector_2 s2539_6(wires_634_5[3], addr_634_5, wires_2539_6,addr_2539_6);

wire[3:0] wires_2540_6;

wire[31:0] addr_2540_6;

Selector_2 s2540_6(wires_635_5[0], addr_635_5, wires_2540_6,addr_2540_6);

wire[3:0] wires_2541_6;

wire[31:0] addr_2541_6;

Selector_2 s2541_6(wires_635_5[1], addr_635_5, wires_2541_6,addr_2541_6);

wire[3:0] wires_2542_6;

wire[31:0] addr_2542_6;

Selector_2 s2542_6(wires_635_5[2], addr_635_5, wires_2542_6,addr_2542_6);

wire[3:0] wires_2543_6;

wire[31:0] addr_2543_6;

Selector_2 s2543_6(wires_635_5[3], addr_635_5, wires_2543_6,addr_2543_6);

wire[3:0] wires_2544_6;

wire[31:0] addr_2544_6;

Selector_2 s2544_6(wires_636_5[0], addr_636_5, wires_2544_6,addr_2544_6);

wire[3:0] wires_2545_6;

wire[31:0] addr_2545_6;

Selector_2 s2545_6(wires_636_5[1], addr_636_5, wires_2545_6,addr_2545_6);

wire[3:0] wires_2546_6;

wire[31:0] addr_2546_6;

Selector_2 s2546_6(wires_636_5[2], addr_636_5, wires_2546_6,addr_2546_6);

wire[3:0] wires_2547_6;

wire[31:0] addr_2547_6;

Selector_2 s2547_6(wires_636_5[3], addr_636_5, wires_2547_6,addr_2547_6);

wire[3:0] wires_2548_6;

wire[31:0] addr_2548_6;

Selector_2 s2548_6(wires_637_5[0], addr_637_5, wires_2548_6,addr_2548_6);

wire[3:0] wires_2549_6;

wire[31:0] addr_2549_6;

Selector_2 s2549_6(wires_637_5[1], addr_637_5, wires_2549_6,addr_2549_6);

wire[3:0] wires_2550_6;

wire[31:0] addr_2550_6;

Selector_2 s2550_6(wires_637_5[2], addr_637_5, wires_2550_6,addr_2550_6);

wire[3:0] wires_2551_6;

wire[31:0] addr_2551_6;

Selector_2 s2551_6(wires_637_5[3], addr_637_5, wires_2551_6,addr_2551_6);

wire[3:0] wires_2552_6;

wire[31:0] addr_2552_6;

Selector_2 s2552_6(wires_638_5[0], addr_638_5, wires_2552_6,addr_2552_6);

wire[3:0] wires_2553_6;

wire[31:0] addr_2553_6;

Selector_2 s2553_6(wires_638_5[1], addr_638_5, wires_2553_6,addr_2553_6);

wire[3:0] wires_2554_6;

wire[31:0] addr_2554_6;

Selector_2 s2554_6(wires_638_5[2], addr_638_5, wires_2554_6,addr_2554_6);

wire[3:0] wires_2555_6;

wire[31:0] addr_2555_6;

Selector_2 s2555_6(wires_638_5[3], addr_638_5, wires_2555_6,addr_2555_6);

wire[3:0] wires_2556_6;

wire[31:0] addr_2556_6;

Selector_2 s2556_6(wires_639_5[0], addr_639_5, wires_2556_6,addr_2556_6);

wire[3:0] wires_2557_6;

wire[31:0] addr_2557_6;

Selector_2 s2557_6(wires_639_5[1], addr_639_5, wires_2557_6,addr_2557_6);

wire[3:0] wires_2558_6;

wire[31:0] addr_2558_6;

Selector_2 s2558_6(wires_639_5[2], addr_639_5, wires_2558_6,addr_2558_6);

wire[3:0] wires_2559_6;

wire[31:0] addr_2559_6;

Selector_2 s2559_6(wires_639_5[3], addr_639_5, wires_2559_6,addr_2559_6);

wire[3:0] wires_2560_6;

wire[31:0] addr_2560_6;

Selector_2 s2560_6(wires_640_5[0], addr_640_5, wires_2560_6,addr_2560_6);

wire[3:0] wires_2561_6;

wire[31:0] addr_2561_6;

Selector_2 s2561_6(wires_640_5[1], addr_640_5, wires_2561_6,addr_2561_6);

wire[3:0] wires_2562_6;

wire[31:0] addr_2562_6;

Selector_2 s2562_6(wires_640_5[2], addr_640_5, wires_2562_6,addr_2562_6);

wire[3:0] wires_2563_6;

wire[31:0] addr_2563_6;

Selector_2 s2563_6(wires_640_5[3], addr_640_5, wires_2563_6,addr_2563_6);

wire[3:0] wires_2564_6;

wire[31:0] addr_2564_6;

Selector_2 s2564_6(wires_641_5[0], addr_641_5, wires_2564_6,addr_2564_6);

wire[3:0] wires_2565_6;

wire[31:0] addr_2565_6;

Selector_2 s2565_6(wires_641_5[1], addr_641_5, wires_2565_6,addr_2565_6);

wire[3:0] wires_2566_6;

wire[31:0] addr_2566_6;

Selector_2 s2566_6(wires_641_5[2], addr_641_5, wires_2566_6,addr_2566_6);

wire[3:0] wires_2567_6;

wire[31:0] addr_2567_6;

Selector_2 s2567_6(wires_641_5[3], addr_641_5, wires_2567_6,addr_2567_6);

wire[3:0] wires_2568_6;

wire[31:0] addr_2568_6;

Selector_2 s2568_6(wires_642_5[0], addr_642_5, wires_2568_6,addr_2568_6);

wire[3:0] wires_2569_6;

wire[31:0] addr_2569_6;

Selector_2 s2569_6(wires_642_5[1], addr_642_5, wires_2569_6,addr_2569_6);

wire[3:0] wires_2570_6;

wire[31:0] addr_2570_6;

Selector_2 s2570_6(wires_642_5[2], addr_642_5, wires_2570_6,addr_2570_6);

wire[3:0] wires_2571_6;

wire[31:0] addr_2571_6;

Selector_2 s2571_6(wires_642_5[3], addr_642_5, wires_2571_6,addr_2571_6);

wire[3:0] wires_2572_6;

wire[31:0] addr_2572_6;

Selector_2 s2572_6(wires_643_5[0], addr_643_5, wires_2572_6,addr_2572_6);

wire[3:0] wires_2573_6;

wire[31:0] addr_2573_6;

Selector_2 s2573_6(wires_643_5[1], addr_643_5, wires_2573_6,addr_2573_6);

wire[3:0] wires_2574_6;

wire[31:0] addr_2574_6;

Selector_2 s2574_6(wires_643_5[2], addr_643_5, wires_2574_6,addr_2574_6);

wire[3:0] wires_2575_6;

wire[31:0] addr_2575_6;

Selector_2 s2575_6(wires_643_5[3], addr_643_5, wires_2575_6,addr_2575_6);

wire[3:0] wires_2576_6;

wire[31:0] addr_2576_6;

Selector_2 s2576_6(wires_644_5[0], addr_644_5, wires_2576_6,addr_2576_6);

wire[3:0] wires_2577_6;

wire[31:0] addr_2577_6;

Selector_2 s2577_6(wires_644_5[1], addr_644_5, wires_2577_6,addr_2577_6);

wire[3:0] wires_2578_6;

wire[31:0] addr_2578_6;

Selector_2 s2578_6(wires_644_5[2], addr_644_5, wires_2578_6,addr_2578_6);

wire[3:0] wires_2579_6;

wire[31:0] addr_2579_6;

Selector_2 s2579_6(wires_644_5[3], addr_644_5, wires_2579_6,addr_2579_6);

wire[3:0] wires_2580_6;

wire[31:0] addr_2580_6;

Selector_2 s2580_6(wires_645_5[0], addr_645_5, wires_2580_6,addr_2580_6);

wire[3:0] wires_2581_6;

wire[31:0] addr_2581_6;

Selector_2 s2581_6(wires_645_5[1], addr_645_5, wires_2581_6,addr_2581_6);

wire[3:0] wires_2582_6;

wire[31:0] addr_2582_6;

Selector_2 s2582_6(wires_645_5[2], addr_645_5, wires_2582_6,addr_2582_6);

wire[3:0] wires_2583_6;

wire[31:0] addr_2583_6;

Selector_2 s2583_6(wires_645_5[3], addr_645_5, wires_2583_6,addr_2583_6);

wire[3:0] wires_2584_6;

wire[31:0] addr_2584_6;

Selector_2 s2584_6(wires_646_5[0], addr_646_5, wires_2584_6,addr_2584_6);

wire[3:0] wires_2585_6;

wire[31:0] addr_2585_6;

Selector_2 s2585_6(wires_646_5[1], addr_646_5, wires_2585_6,addr_2585_6);

wire[3:0] wires_2586_6;

wire[31:0] addr_2586_6;

Selector_2 s2586_6(wires_646_5[2], addr_646_5, wires_2586_6,addr_2586_6);

wire[3:0] wires_2587_6;

wire[31:0] addr_2587_6;

Selector_2 s2587_6(wires_646_5[3], addr_646_5, wires_2587_6,addr_2587_6);

wire[3:0] wires_2588_6;

wire[31:0] addr_2588_6;

Selector_2 s2588_6(wires_647_5[0], addr_647_5, wires_2588_6,addr_2588_6);

wire[3:0] wires_2589_6;

wire[31:0] addr_2589_6;

Selector_2 s2589_6(wires_647_5[1], addr_647_5, wires_2589_6,addr_2589_6);

wire[3:0] wires_2590_6;

wire[31:0] addr_2590_6;

Selector_2 s2590_6(wires_647_5[2], addr_647_5, wires_2590_6,addr_2590_6);

wire[3:0] wires_2591_6;

wire[31:0] addr_2591_6;

Selector_2 s2591_6(wires_647_5[3], addr_647_5, wires_2591_6,addr_2591_6);

wire[3:0] wires_2592_6;

wire[31:0] addr_2592_6;

Selector_2 s2592_6(wires_648_5[0], addr_648_5, wires_2592_6,addr_2592_6);

wire[3:0] wires_2593_6;

wire[31:0] addr_2593_6;

Selector_2 s2593_6(wires_648_5[1], addr_648_5, wires_2593_6,addr_2593_6);

wire[3:0] wires_2594_6;

wire[31:0] addr_2594_6;

Selector_2 s2594_6(wires_648_5[2], addr_648_5, wires_2594_6,addr_2594_6);

wire[3:0] wires_2595_6;

wire[31:0] addr_2595_6;

Selector_2 s2595_6(wires_648_5[3], addr_648_5, wires_2595_6,addr_2595_6);

wire[3:0] wires_2596_6;

wire[31:0] addr_2596_6;

Selector_2 s2596_6(wires_649_5[0], addr_649_5, wires_2596_6,addr_2596_6);

wire[3:0] wires_2597_6;

wire[31:0] addr_2597_6;

Selector_2 s2597_6(wires_649_5[1], addr_649_5, wires_2597_6,addr_2597_6);

wire[3:0] wires_2598_6;

wire[31:0] addr_2598_6;

Selector_2 s2598_6(wires_649_5[2], addr_649_5, wires_2598_6,addr_2598_6);

wire[3:0] wires_2599_6;

wire[31:0] addr_2599_6;

Selector_2 s2599_6(wires_649_5[3], addr_649_5, wires_2599_6,addr_2599_6);

wire[3:0] wires_2600_6;

wire[31:0] addr_2600_6;

Selector_2 s2600_6(wires_650_5[0], addr_650_5, wires_2600_6,addr_2600_6);

wire[3:0] wires_2601_6;

wire[31:0] addr_2601_6;

Selector_2 s2601_6(wires_650_5[1], addr_650_5, wires_2601_6,addr_2601_6);

wire[3:0] wires_2602_6;

wire[31:0] addr_2602_6;

Selector_2 s2602_6(wires_650_5[2], addr_650_5, wires_2602_6,addr_2602_6);

wire[3:0] wires_2603_6;

wire[31:0] addr_2603_6;

Selector_2 s2603_6(wires_650_5[3], addr_650_5, wires_2603_6,addr_2603_6);

wire[3:0] wires_2604_6;

wire[31:0] addr_2604_6;

Selector_2 s2604_6(wires_651_5[0], addr_651_5, wires_2604_6,addr_2604_6);

wire[3:0] wires_2605_6;

wire[31:0] addr_2605_6;

Selector_2 s2605_6(wires_651_5[1], addr_651_5, wires_2605_6,addr_2605_6);

wire[3:0] wires_2606_6;

wire[31:0] addr_2606_6;

Selector_2 s2606_6(wires_651_5[2], addr_651_5, wires_2606_6,addr_2606_6);

wire[3:0] wires_2607_6;

wire[31:0] addr_2607_6;

Selector_2 s2607_6(wires_651_5[3], addr_651_5, wires_2607_6,addr_2607_6);

wire[3:0] wires_2608_6;

wire[31:0] addr_2608_6;

Selector_2 s2608_6(wires_652_5[0], addr_652_5, wires_2608_6,addr_2608_6);

wire[3:0] wires_2609_6;

wire[31:0] addr_2609_6;

Selector_2 s2609_6(wires_652_5[1], addr_652_5, wires_2609_6,addr_2609_6);

wire[3:0] wires_2610_6;

wire[31:0] addr_2610_6;

Selector_2 s2610_6(wires_652_5[2], addr_652_5, wires_2610_6,addr_2610_6);

wire[3:0] wires_2611_6;

wire[31:0] addr_2611_6;

Selector_2 s2611_6(wires_652_5[3], addr_652_5, wires_2611_6,addr_2611_6);

wire[3:0] wires_2612_6;

wire[31:0] addr_2612_6;

Selector_2 s2612_6(wires_653_5[0], addr_653_5, wires_2612_6,addr_2612_6);

wire[3:0] wires_2613_6;

wire[31:0] addr_2613_6;

Selector_2 s2613_6(wires_653_5[1], addr_653_5, wires_2613_6,addr_2613_6);

wire[3:0] wires_2614_6;

wire[31:0] addr_2614_6;

Selector_2 s2614_6(wires_653_5[2], addr_653_5, wires_2614_6,addr_2614_6);

wire[3:0] wires_2615_6;

wire[31:0] addr_2615_6;

Selector_2 s2615_6(wires_653_5[3], addr_653_5, wires_2615_6,addr_2615_6);

wire[3:0] wires_2616_6;

wire[31:0] addr_2616_6;

Selector_2 s2616_6(wires_654_5[0], addr_654_5, wires_2616_6,addr_2616_6);

wire[3:0] wires_2617_6;

wire[31:0] addr_2617_6;

Selector_2 s2617_6(wires_654_5[1], addr_654_5, wires_2617_6,addr_2617_6);

wire[3:0] wires_2618_6;

wire[31:0] addr_2618_6;

Selector_2 s2618_6(wires_654_5[2], addr_654_5, wires_2618_6,addr_2618_6);

wire[3:0] wires_2619_6;

wire[31:0] addr_2619_6;

Selector_2 s2619_6(wires_654_5[3], addr_654_5, wires_2619_6,addr_2619_6);

wire[3:0] wires_2620_6;

wire[31:0] addr_2620_6;

Selector_2 s2620_6(wires_655_5[0], addr_655_5, wires_2620_6,addr_2620_6);

wire[3:0] wires_2621_6;

wire[31:0] addr_2621_6;

Selector_2 s2621_6(wires_655_5[1], addr_655_5, wires_2621_6,addr_2621_6);

wire[3:0] wires_2622_6;

wire[31:0] addr_2622_6;

Selector_2 s2622_6(wires_655_5[2], addr_655_5, wires_2622_6,addr_2622_6);

wire[3:0] wires_2623_6;

wire[31:0] addr_2623_6;

Selector_2 s2623_6(wires_655_5[3], addr_655_5, wires_2623_6,addr_2623_6);

wire[3:0] wires_2624_6;

wire[31:0] addr_2624_6;

Selector_2 s2624_6(wires_656_5[0], addr_656_5, wires_2624_6,addr_2624_6);

wire[3:0] wires_2625_6;

wire[31:0] addr_2625_6;

Selector_2 s2625_6(wires_656_5[1], addr_656_5, wires_2625_6,addr_2625_6);

wire[3:0] wires_2626_6;

wire[31:0] addr_2626_6;

Selector_2 s2626_6(wires_656_5[2], addr_656_5, wires_2626_6,addr_2626_6);

wire[3:0] wires_2627_6;

wire[31:0] addr_2627_6;

Selector_2 s2627_6(wires_656_5[3], addr_656_5, wires_2627_6,addr_2627_6);

wire[3:0] wires_2628_6;

wire[31:0] addr_2628_6;

Selector_2 s2628_6(wires_657_5[0], addr_657_5, wires_2628_6,addr_2628_6);

wire[3:0] wires_2629_6;

wire[31:0] addr_2629_6;

Selector_2 s2629_6(wires_657_5[1], addr_657_5, wires_2629_6,addr_2629_6);

wire[3:0] wires_2630_6;

wire[31:0] addr_2630_6;

Selector_2 s2630_6(wires_657_5[2], addr_657_5, wires_2630_6,addr_2630_6);

wire[3:0] wires_2631_6;

wire[31:0] addr_2631_6;

Selector_2 s2631_6(wires_657_5[3], addr_657_5, wires_2631_6,addr_2631_6);

wire[3:0] wires_2632_6;

wire[31:0] addr_2632_6;

Selector_2 s2632_6(wires_658_5[0], addr_658_5, wires_2632_6,addr_2632_6);

wire[3:0] wires_2633_6;

wire[31:0] addr_2633_6;

Selector_2 s2633_6(wires_658_5[1], addr_658_5, wires_2633_6,addr_2633_6);

wire[3:0] wires_2634_6;

wire[31:0] addr_2634_6;

Selector_2 s2634_6(wires_658_5[2], addr_658_5, wires_2634_6,addr_2634_6);

wire[3:0] wires_2635_6;

wire[31:0] addr_2635_6;

Selector_2 s2635_6(wires_658_5[3], addr_658_5, wires_2635_6,addr_2635_6);

wire[3:0] wires_2636_6;

wire[31:0] addr_2636_6;

Selector_2 s2636_6(wires_659_5[0], addr_659_5, wires_2636_6,addr_2636_6);

wire[3:0] wires_2637_6;

wire[31:0] addr_2637_6;

Selector_2 s2637_6(wires_659_5[1], addr_659_5, wires_2637_6,addr_2637_6);

wire[3:0] wires_2638_6;

wire[31:0] addr_2638_6;

Selector_2 s2638_6(wires_659_5[2], addr_659_5, wires_2638_6,addr_2638_6);

wire[3:0] wires_2639_6;

wire[31:0] addr_2639_6;

Selector_2 s2639_6(wires_659_5[3], addr_659_5, wires_2639_6,addr_2639_6);

wire[3:0] wires_2640_6;

wire[31:0] addr_2640_6;

Selector_2 s2640_6(wires_660_5[0], addr_660_5, wires_2640_6,addr_2640_6);

wire[3:0] wires_2641_6;

wire[31:0] addr_2641_6;

Selector_2 s2641_6(wires_660_5[1], addr_660_5, wires_2641_6,addr_2641_6);

wire[3:0] wires_2642_6;

wire[31:0] addr_2642_6;

Selector_2 s2642_6(wires_660_5[2], addr_660_5, wires_2642_6,addr_2642_6);

wire[3:0] wires_2643_6;

wire[31:0] addr_2643_6;

Selector_2 s2643_6(wires_660_5[3], addr_660_5, wires_2643_6,addr_2643_6);

wire[3:0] wires_2644_6;

wire[31:0] addr_2644_6;

Selector_2 s2644_6(wires_661_5[0], addr_661_5, wires_2644_6,addr_2644_6);

wire[3:0] wires_2645_6;

wire[31:0] addr_2645_6;

Selector_2 s2645_6(wires_661_5[1], addr_661_5, wires_2645_6,addr_2645_6);

wire[3:0] wires_2646_6;

wire[31:0] addr_2646_6;

Selector_2 s2646_6(wires_661_5[2], addr_661_5, wires_2646_6,addr_2646_6);

wire[3:0] wires_2647_6;

wire[31:0] addr_2647_6;

Selector_2 s2647_6(wires_661_5[3], addr_661_5, wires_2647_6,addr_2647_6);

wire[3:0] wires_2648_6;

wire[31:0] addr_2648_6;

Selector_2 s2648_6(wires_662_5[0], addr_662_5, wires_2648_6,addr_2648_6);

wire[3:0] wires_2649_6;

wire[31:0] addr_2649_6;

Selector_2 s2649_6(wires_662_5[1], addr_662_5, wires_2649_6,addr_2649_6);

wire[3:0] wires_2650_6;

wire[31:0] addr_2650_6;

Selector_2 s2650_6(wires_662_5[2], addr_662_5, wires_2650_6,addr_2650_6);

wire[3:0] wires_2651_6;

wire[31:0] addr_2651_6;

Selector_2 s2651_6(wires_662_5[3], addr_662_5, wires_2651_6,addr_2651_6);

wire[3:0] wires_2652_6;

wire[31:0] addr_2652_6;

Selector_2 s2652_6(wires_663_5[0], addr_663_5, wires_2652_6,addr_2652_6);

wire[3:0] wires_2653_6;

wire[31:0] addr_2653_6;

Selector_2 s2653_6(wires_663_5[1], addr_663_5, wires_2653_6,addr_2653_6);

wire[3:0] wires_2654_6;

wire[31:0] addr_2654_6;

Selector_2 s2654_6(wires_663_5[2], addr_663_5, wires_2654_6,addr_2654_6);

wire[3:0] wires_2655_6;

wire[31:0] addr_2655_6;

Selector_2 s2655_6(wires_663_5[3], addr_663_5, wires_2655_6,addr_2655_6);

wire[3:0] wires_2656_6;

wire[31:0] addr_2656_6;

Selector_2 s2656_6(wires_664_5[0], addr_664_5, wires_2656_6,addr_2656_6);

wire[3:0] wires_2657_6;

wire[31:0] addr_2657_6;

Selector_2 s2657_6(wires_664_5[1], addr_664_5, wires_2657_6,addr_2657_6);

wire[3:0] wires_2658_6;

wire[31:0] addr_2658_6;

Selector_2 s2658_6(wires_664_5[2], addr_664_5, wires_2658_6,addr_2658_6);

wire[3:0] wires_2659_6;

wire[31:0] addr_2659_6;

Selector_2 s2659_6(wires_664_5[3], addr_664_5, wires_2659_6,addr_2659_6);

wire[3:0] wires_2660_6;

wire[31:0] addr_2660_6;

Selector_2 s2660_6(wires_665_5[0], addr_665_5, wires_2660_6,addr_2660_6);

wire[3:0] wires_2661_6;

wire[31:0] addr_2661_6;

Selector_2 s2661_6(wires_665_5[1], addr_665_5, wires_2661_6,addr_2661_6);

wire[3:0] wires_2662_6;

wire[31:0] addr_2662_6;

Selector_2 s2662_6(wires_665_5[2], addr_665_5, wires_2662_6,addr_2662_6);

wire[3:0] wires_2663_6;

wire[31:0] addr_2663_6;

Selector_2 s2663_6(wires_665_5[3], addr_665_5, wires_2663_6,addr_2663_6);

wire[3:0] wires_2664_6;

wire[31:0] addr_2664_6;

Selector_2 s2664_6(wires_666_5[0], addr_666_5, wires_2664_6,addr_2664_6);

wire[3:0] wires_2665_6;

wire[31:0] addr_2665_6;

Selector_2 s2665_6(wires_666_5[1], addr_666_5, wires_2665_6,addr_2665_6);

wire[3:0] wires_2666_6;

wire[31:0] addr_2666_6;

Selector_2 s2666_6(wires_666_5[2], addr_666_5, wires_2666_6,addr_2666_6);

wire[3:0] wires_2667_6;

wire[31:0] addr_2667_6;

Selector_2 s2667_6(wires_666_5[3], addr_666_5, wires_2667_6,addr_2667_6);

wire[3:0] wires_2668_6;

wire[31:0] addr_2668_6;

Selector_2 s2668_6(wires_667_5[0], addr_667_5, wires_2668_6,addr_2668_6);

wire[3:0] wires_2669_6;

wire[31:0] addr_2669_6;

Selector_2 s2669_6(wires_667_5[1], addr_667_5, wires_2669_6,addr_2669_6);

wire[3:0] wires_2670_6;

wire[31:0] addr_2670_6;

Selector_2 s2670_6(wires_667_5[2], addr_667_5, wires_2670_6,addr_2670_6);

wire[3:0] wires_2671_6;

wire[31:0] addr_2671_6;

Selector_2 s2671_6(wires_667_5[3], addr_667_5, wires_2671_6,addr_2671_6);

wire[3:0] wires_2672_6;

wire[31:0] addr_2672_6;

Selector_2 s2672_6(wires_668_5[0], addr_668_5, wires_2672_6,addr_2672_6);

wire[3:0] wires_2673_6;

wire[31:0] addr_2673_6;

Selector_2 s2673_6(wires_668_5[1], addr_668_5, wires_2673_6,addr_2673_6);

wire[3:0] wires_2674_6;

wire[31:0] addr_2674_6;

Selector_2 s2674_6(wires_668_5[2], addr_668_5, wires_2674_6,addr_2674_6);

wire[3:0] wires_2675_6;

wire[31:0] addr_2675_6;

Selector_2 s2675_6(wires_668_5[3], addr_668_5, wires_2675_6,addr_2675_6);

wire[3:0] wires_2676_6;

wire[31:0] addr_2676_6;

Selector_2 s2676_6(wires_669_5[0], addr_669_5, wires_2676_6,addr_2676_6);

wire[3:0] wires_2677_6;

wire[31:0] addr_2677_6;

Selector_2 s2677_6(wires_669_5[1], addr_669_5, wires_2677_6,addr_2677_6);

wire[3:0] wires_2678_6;

wire[31:0] addr_2678_6;

Selector_2 s2678_6(wires_669_5[2], addr_669_5, wires_2678_6,addr_2678_6);

wire[3:0] wires_2679_6;

wire[31:0] addr_2679_6;

Selector_2 s2679_6(wires_669_5[3], addr_669_5, wires_2679_6,addr_2679_6);

wire[3:0] wires_2680_6;

wire[31:0] addr_2680_6;

Selector_2 s2680_6(wires_670_5[0], addr_670_5, wires_2680_6,addr_2680_6);

wire[3:0] wires_2681_6;

wire[31:0] addr_2681_6;

Selector_2 s2681_6(wires_670_5[1], addr_670_5, wires_2681_6,addr_2681_6);

wire[3:0] wires_2682_6;

wire[31:0] addr_2682_6;

Selector_2 s2682_6(wires_670_5[2], addr_670_5, wires_2682_6,addr_2682_6);

wire[3:0] wires_2683_6;

wire[31:0] addr_2683_6;

Selector_2 s2683_6(wires_670_5[3], addr_670_5, wires_2683_6,addr_2683_6);

wire[3:0] wires_2684_6;

wire[31:0] addr_2684_6;

Selector_2 s2684_6(wires_671_5[0], addr_671_5, wires_2684_6,addr_2684_6);

wire[3:0] wires_2685_6;

wire[31:0] addr_2685_6;

Selector_2 s2685_6(wires_671_5[1], addr_671_5, wires_2685_6,addr_2685_6);

wire[3:0] wires_2686_6;

wire[31:0] addr_2686_6;

Selector_2 s2686_6(wires_671_5[2], addr_671_5, wires_2686_6,addr_2686_6);

wire[3:0] wires_2687_6;

wire[31:0] addr_2687_6;

Selector_2 s2687_6(wires_671_5[3], addr_671_5, wires_2687_6,addr_2687_6);

wire[3:0] wires_2688_6;

wire[31:0] addr_2688_6;

Selector_2 s2688_6(wires_672_5[0], addr_672_5, wires_2688_6,addr_2688_6);

wire[3:0] wires_2689_6;

wire[31:0] addr_2689_6;

Selector_2 s2689_6(wires_672_5[1], addr_672_5, wires_2689_6,addr_2689_6);

wire[3:0] wires_2690_6;

wire[31:0] addr_2690_6;

Selector_2 s2690_6(wires_672_5[2], addr_672_5, wires_2690_6,addr_2690_6);

wire[3:0] wires_2691_6;

wire[31:0] addr_2691_6;

Selector_2 s2691_6(wires_672_5[3], addr_672_5, wires_2691_6,addr_2691_6);

wire[3:0] wires_2692_6;

wire[31:0] addr_2692_6;

Selector_2 s2692_6(wires_673_5[0], addr_673_5, wires_2692_6,addr_2692_6);

wire[3:0] wires_2693_6;

wire[31:0] addr_2693_6;

Selector_2 s2693_6(wires_673_5[1], addr_673_5, wires_2693_6,addr_2693_6);

wire[3:0] wires_2694_6;

wire[31:0] addr_2694_6;

Selector_2 s2694_6(wires_673_5[2], addr_673_5, wires_2694_6,addr_2694_6);

wire[3:0] wires_2695_6;

wire[31:0] addr_2695_6;

Selector_2 s2695_6(wires_673_5[3], addr_673_5, wires_2695_6,addr_2695_6);

wire[3:0] wires_2696_6;

wire[31:0] addr_2696_6;

Selector_2 s2696_6(wires_674_5[0], addr_674_5, wires_2696_6,addr_2696_6);

wire[3:0] wires_2697_6;

wire[31:0] addr_2697_6;

Selector_2 s2697_6(wires_674_5[1], addr_674_5, wires_2697_6,addr_2697_6);

wire[3:0] wires_2698_6;

wire[31:0] addr_2698_6;

Selector_2 s2698_6(wires_674_5[2], addr_674_5, wires_2698_6,addr_2698_6);

wire[3:0] wires_2699_6;

wire[31:0] addr_2699_6;

Selector_2 s2699_6(wires_674_5[3], addr_674_5, wires_2699_6,addr_2699_6);

wire[3:0] wires_2700_6;

wire[31:0] addr_2700_6;

Selector_2 s2700_6(wires_675_5[0], addr_675_5, wires_2700_6,addr_2700_6);

wire[3:0] wires_2701_6;

wire[31:0] addr_2701_6;

Selector_2 s2701_6(wires_675_5[1], addr_675_5, wires_2701_6,addr_2701_6);

wire[3:0] wires_2702_6;

wire[31:0] addr_2702_6;

Selector_2 s2702_6(wires_675_5[2], addr_675_5, wires_2702_6,addr_2702_6);

wire[3:0] wires_2703_6;

wire[31:0] addr_2703_6;

Selector_2 s2703_6(wires_675_5[3], addr_675_5, wires_2703_6,addr_2703_6);

wire[3:0] wires_2704_6;

wire[31:0] addr_2704_6;

Selector_2 s2704_6(wires_676_5[0], addr_676_5, wires_2704_6,addr_2704_6);

wire[3:0] wires_2705_6;

wire[31:0] addr_2705_6;

Selector_2 s2705_6(wires_676_5[1], addr_676_5, wires_2705_6,addr_2705_6);

wire[3:0] wires_2706_6;

wire[31:0] addr_2706_6;

Selector_2 s2706_6(wires_676_5[2], addr_676_5, wires_2706_6,addr_2706_6);

wire[3:0] wires_2707_6;

wire[31:0] addr_2707_6;

Selector_2 s2707_6(wires_676_5[3], addr_676_5, wires_2707_6,addr_2707_6);

wire[3:0] wires_2708_6;

wire[31:0] addr_2708_6;

Selector_2 s2708_6(wires_677_5[0], addr_677_5, wires_2708_6,addr_2708_6);

wire[3:0] wires_2709_6;

wire[31:0] addr_2709_6;

Selector_2 s2709_6(wires_677_5[1], addr_677_5, wires_2709_6,addr_2709_6);

wire[3:0] wires_2710_6;

wire[31:0] addr_2710_6;

Selector_2 s2710_6(wires_677_5[2], addr_677_5, wires_2710_6,addr_2710_6);

wire[3:0] wires_2711_6;

wire[31:0] addr_2711_6;

Selector_2 s2711_6(wires_677_5[3], addr_677_5, wires_2711_6,addr_2711_6);

wire[3:0] wires_2712_6;

wire[31:0] addr_2712_6;

Selector_2 s2712_6(wires_678_5[0], addr_678_5, wires_2712_6,addr_2712_6);

wire[3:0] wires_2713_6;

wire[31:0] addr_2713_6;

Selector_2 s2713_6(wires_678_5[1], addr_678_5, wires_2713_6,addr_2713_6);

wire[3:0] wires_2714_6;

wire[31:0] addr_2714_6;

Selector_2 s2714_6(wires_678_5[2], addr_678_5, wires_2714_6,addr_2714_6);

wire[3:0] wires_2715_6;

wire[31:0] addr_2715_6;

Selector_2 s2715_6(wires_678_5[3], addr_678_5, wires_2715_6,addr_2715_6);

wire[3:0] wires_2716_6;

wire[31:0] addr_2716_6;

Selector_2 s2716_6(wires_679_5[0], addr_679_5, wires_2716_6,addr_2716_6);

wire[3:0] wires_2717_6;

wire[31:0] addr_2717_6;

Selector_2 s2717_6(wires_679_5[1], addr_679_5, wires_2717_6,addr_2717_6);

wire[3:0] wires_2718_6;

wire[31:0] addr_2718_6;

Selector_2 s2718_6(wires_679_5[2], addr_679_5, wires_2718_6,addr_2718_6);

wire[3:0] wires_2719_6;

wire[31:0] addr_2719_6;

Selector_2 s2719_6(wires_679_5[3], addr_679_5, wires_2719_6,addr_2719_6);

wire[3:0] wires_2720_6;

wire[31:0] addr_2720_6;

Selector_2 s2720_6(wires_680_5[0], addr_680_5, wires_2720_6,addr_2720_6);

wire[3:0] wires_2721_6;

wire[31:0] addr_2721_6;

Selector_2 s2721_6(wires_680_5[1], addr_680_5, wires_2721_6,addr_2721_6);

wire[3:0] wires_2722_6;

wire[31:0] addr_2722_6;

Selector_2 s2722_6(wires_680_5[2], addr_680_5, wires_2722_6,addr_2722_6);

wire[3:0] wires_2723_6;

wire[31:0] addr_2723_6;

Selector_2 s2723_6(wires_680_5[3], addr_680_5, wires_2723_6,addr_2723_6);

wire[3:0] wires_2724_6;

wire[31:0] addr_2724_6;

Selector_2 s2724_6(wires_681_5[0], addr_681_5, wires_2724_6,addr_2724_6);

wire[3:0] wires_2725_6;

wire[31:0] addr_2725_6;

Selector_2 s2725_6(wires_681_5[1], addr_681_5, wires_2725_6,addr_2725_6);

wire[3:0] wires_2726_6;

wire[31:0] addr_2726_6;

Selector_2 s2726_6(wires_681_5[2], addr_681_5, wires_2726_6,addr_2726_6);

wire[3:0] wires_2727_6;

wire[31:0] addr_2727_6;

Selector_2 s2727_6(wires_681_5[3], addr_681_5, wires_2727_6,addr_2727_6);

wire[3:0] wires_2728_6;

wire[31:0] addr_2728_6;

Selector_2 s2728_6(wires_682_5[0], addr_682_5, wires_2728_6,addr_2728_6);

wire[3:0] wires_2729_6;

wire[31:0] addr_2729_6;

Selector_2 s2729_6(wires_682_5[1], addr_682_5, wires_2729_6,addr_2729_6);

wire[3:0] wires_2730_6;

wire[31:0] addr_2730_6;

Selector_2 s2730_6(wires_682_5[2], addr_682_5, wires_2730_6,addr_2730_6);

wire[3:0] wires_2731_6;

wire[31:0] addr_2731_6;

Selector_2 s2731_6(wires_682_5[3], addr_682_5, wires_2731_6,addr_2731_6);

wire[3:0] wires_2732_6;

wire[31:0] addr_2732_6;

Selector_2 s2732_6(wires_683_5[0], addr_683_5, wires_2732_6,addr_2732_6);

wire[3:0] wires_2733_6;

wire[31:0] addr_2733_6;

Selector_2 s2733_6(wires_683_5[1], addr_683_5, wires_2733_6,addr_2733_6);

wire[3:0] wires_2734_6;

wire[31:0] addr_2734_6;

Selector_2 s2734_6(wires_683_5[2], addr_683_5, wires_2734_6,addr_2734_6);

wire[3:0] wires_2735_6;

wire[31:0] addr_2735_6;

Selector_2 s2735_6(wires_683_5[3], addr_683_5, wires_2735_6,addr_2735_6);

wire[3:0] wires_2736_6;

wire[31:0] addr_2736_6;

Selector_2 s2736_6(wires_684_5[0], addr_684_5, wires_2736_6,addr_2736_6);

wire[3:0] wires_2737_6;

wire[31:0] addr_2737_6;

Selector_2 s2737_6(wires_684_5[1], addr_684_5, wires_2737_6,addr_2737_6);

wire[3:0] wires_2738_6;

wire[31:0] addr_2738_6;

Selector_2 s2738_6(wires_684_5[2], addr_684_5, wires_2738_6,addr_2738_6);

wire[3:0] wires_2739_6;

wire[31:0] addr_2739_6;

Selector_2 s2739_6(wires_684_5[3], addr_684_5, wires_2739_6,addr_2739_6);

wire[3:0] wires_2740_6;

wire[31:0] addr_2740_6;

Selector_2 s2740_6(wires_685_5[0], addr_685_5, wires_2740_6,addr_2740_6);

wire[3:0] wires_2741_6;

wire[31:0] addr_2741_6;

Selector_2 s2741_6(wires_685_5[1], addr_685_5, wires_2741_6,addr_2741_6);

wire[3:0] wires_2742_6;

wire[31:0] addr_2742_6;

Selector_2 s2742_6(wires_685_5[2], addr_685_5, wires_2742_6,addr_2742_6);

wire[3:0] wires_2743_6;

wire[31:0] addr_2743_6;

Selector_2 s2743_6(wires_685_5[3], addr_685_5, wires_2743_6,addr_2743_6);

wire[3:0] wires_2744_6;

wire[31:0] addr_2744_6;

Selector_2 s2744_6(wires_686_5[0], addr_686_5, wires_2744_6,addr_2744_6);

wire[3:0] wires_2745_6;

wire[31:0] addr_2745_6;

Selector_2 s2745_6(wires_686_5[1], addr_686_5, wires_2745_6,addr_2745_6);

wire[3:0] wires_2746_6;

wire[31:0] addr_2746_6;

Selector_2 s2746_6(wires_686_5[2], addr_686_5, wires_2746_6,addr_2746_6);

wire[3:0] wires_2747_6;

wire[31:0] addr_2747_6;

Selector_2 s2747_6(wires_686_5[3], addr_686_5, wires_2747_6,addr_2747_6);

wire[3:0] wires_2748_6;

wire[31:0] addr_2748_6;

Selector_2 s2748_6(wires_687_5[0], addr_687_5, wires_2748_6,addr_2748_6);

wire[3:0] wires_2749_6;

wire[31:0] addr_2749_6;

Selector_2 s2749_6(wires_687_5[1], addr_687_5, wires_2749_6,addr_2749_6);

wire[3:0] wires_2750_6;

wire[31:0] addr_2750_6;

Selector_2 s2750_6(wires_687_5[2], addr_687_5, wires_2750_6,addr_2750_6);

wire[3:0] wires_2751_6;

wire[31:0] addr_2751_6;

Selector_2 s2751_6(wires_687_5[3], addr_687_5, wires_2751_6,addr_2751_6);

wire[3:0] wires_2752_6;

wire[31:0] addr_2752_6;

Selector_2 s2752_6(wires_688_5[0], addr_688_5, wires_2752_6,addr_2752_6);

wire[3:0] wires_2753_6;

wire[31:0] addr_2753_6;

Selector_2 s2753_6(wires_688_5[1], addr_688_5, wires_2753_6,addr_2753_6);

wire[3:0] wires_2754_6;

wire[31:0] addr_2754_6;

Selector_2 s2754_6(wires_688_5[2], addr_688_5, wires_2754_6,addr_2754_6);

wire[3:0] wires_2755_6;

wire[31:0] addr_2755_6;

Selector_2 s2755_6(wires_688_5[3], addr_688_5, wires_2755_6,addr_2755_6);

wire[3:0] wires_2756_6;

wire[31:0] addr_2756_6;

Selector_2 s2756_6(wires_689_5[0], addr_689_5, wires_2756_6,addr_2756_6);

wire[3:0] wires_2757_6;

wire[31:0] addr_2757_6;

Selector_2 s2757_6(wires_689_5[1], addr_689_5, wires_2757_6,addr_2757_6);

wire[3:0] wires_2758_6;

wire[31:0] addr_2758_6;

Selector_2 s2758_6(wires_689_5[2], addr_689_5, wires_2758_6,addr_2758_6);

wire[3:0] wires_2759_6;

wire[31:0] addr_2759_6;

Selector_2 s2759_6(wires_689_5[3], addr_689_5, wires_2759_6,addr_2759_6);

wire[3:0] wires_2760_6;

wire[31:0] addr_2760_6;

Selector_2 s2760_6(wires_690_5[0], addr_690_5, wires_2760_6,addr_2760_6);

wire[3:0] wires_2761_6;

wire[31:0] addr_2761_6;

Selector_2 s2761_6(wires_690_5[1], addr_690_5, wires_2761_6,addr_2761_6);

wire[3:0] wires_2762_6;

wire[31:0] addr_2762_6;

Selector_2 s2762_6(wires_690_5[2], addr_690_5, wires_2762_6,addr_2762_6);

wire[3:0] wires_2763_6;

wire[31:0] addr_2763_6;

Selector_2 s2763_6(wires_690_5[3], addr_690_5, wires_2763_6,addr_2763_6);

wire[3:0] wires_2764_6;

wire[31:0] addr_2764_6;

Selector_2 s2764_6(wires_691_5[0], addr_691_5, wires_2764_6,addr_2764_6);

wire[3:0] wires_2765_6;

wire[31:0] addr_2765_6;

Selector_2 s2765_6(wires_691_5[1], addr_691_5, wires_2765_6,addr_2765_6);

wire[3:0] wires_2766_6;

wire[31:0] addr_2766_6;

Selector_2 s2766_6(wires_691_5[2], addr_691_5, wires_2766_6,addr_2766_6);

wire[3:0] wires_2767_6;

wire[31:0] addr_2767_6;

Selector_2 s2767_6(wires_691_5[3], addr_691_5, wires_2767_6,addr_2767_6);

wire[3:0] wires_2768_6;

wire[31:0] addr_2768_6;

Selector_2 s2768_6(wires_692_5[0], addr_692_5, wires_2768_6,addr_2768_6);

wire[3:0] wires_2769_6;

wire[31:0] addr_2769_6;

Selector_2 s2769_6(wires_692_5[1], addr_692_5, wires_2769_6,addr_2769_6);

wire[3:0] wires_2770_6;

wire[31:0] addr_2770_6;

Selector_2 s2770_6(wires_692_5[2], addr_692_5, wires_2770_6,addr_2770_6);

wire[3:0] wires_2771_6;

wire[31:0] addr_2771_6;

Selector_2 s2771_6(wires_692_5[3], addr_692_5, wires_2771_6,addr_2771_6);

wire[3:0] wires_2772_6;

wire[31:0] addr_2772_6;

Selector_2 s2772_6(wires_693_5[0], addr_693_5, wires_2772_6,addr_2772_6);

wire[3:0] wires_2773_6;

wire[31:0] addr_2773_6;

Selector_2 s2773_6(wires_693_5[1], addr_693_5, wires_2773_6,addr_2773_6);

wire[3:0] wires_2774_6;

wire[31:0] addr_2774_6;

Selector_2 s2774_6(wires_693_5[2], addr_693_5, wires_2774_6,addr_2774_6);

wire[3:0] wires_2775_6;

wire[31:0] addr_2775_6;

Selector_2 s2775_6(wires_693_5[3], addr_693_5, wires_2775_6,addr_2775_6);

wire[3:0] wires_2776_6;

wire[31:0] addr_2776_6;

Selector_2 s2776_6(wires_694_5[0], addr_694_5, wires_2776_6,addr_2776_6);

wire[3:0] wires_2777_6;

wire[31:0] addr_2777_6;

Selector_2 s2777_6(wires_694_5[1], addr_694_5, wires_2777_6,addr_2777_6);

wire[3:0] wires_2778_6;

wire[31:0] addr_2778_6;

Selector_2 s2778_6(wires_694_5[2], addr_694_5, wires_2778_6,addr_2778_6);

wire[3:0] wires_2779_6;

wire[31:0] addr_2779_6;

Selector_2 s2779_6(wires_694_5[3], addr_694_5, wires_2779_6,addr_2779_6);

wire[3:0] wires_2780_6;

wire[31:0] addr_2780_6;

Selector_2 s2780_6(wires_695_5[0], addr_695_5, wires_2780_6,addr_2780_6);

wire[3:0] wires_2781_6;

wire[31:0] addr_2781_6;

Selector_2 s2781_6(wires_695_5[1], addr_695_5, wires_2781_6,addr_2781_6);

wire[3:0] wires_2782_6;

wire[31:0] addr_2782_6;

Selector_2 s2782_6(wires_695_5[2], addr_695_5, wires_2782_6,addr_2782_6);

wire[3:0] wires_2783_6;

wire[31:0] addr_2783_6;

Selector_2 s2783_6(wires_695_5[3], addr_695_5, wires_2783_6,addr_2783_6);

wire[3:0] wires_2784_6;

wire[31:0] addr_2784_6;

Selector_2 s2784_6(wires_696_5[0], addr_696_5, wires_2784_6,addr_2784_6);

wire[3:0] wires_2785_6;

wire[31:0] addr_2785_6;

Selector_2 s2785_6(wires_696_5[1], addr_696_5, wires_2785_6,addr_2785_6);

wire[3:0] wires_2786_6;

wire[31:0] addr_2786_6;

Selector_2 s2786_6(wires_696_5[2], addr_696_5, wires_2786_6,addr_2786_6);

wire[3:0] wires_2787_6;

wire[31:0] addr_2787_6;

Selector_2 s2787_6(wires_696_5[3], addr_696_5, wires_2787_6,addr_2787_6);

wire[3:0] wires_2788_6;

wire[31:0] addr_2788_6;

Selector_2 s2788_6(wires_697_5[0], addr_697_5, wires_2788_6,addr_2788_6);

wire[3:0] wires_2789_6;

wire[31:0] addr_2789_6;

Selector_2 s2789_6(wires_697_5[1], addr_697_5, wires_2789_6,addr_2789_6);

wire[3:0] wires_2790_6;

wire[31:0] addr_2790_6;

Selector_2 s2790_6(wires_697_5[2], addr_697_5, wires_2790_6,addr_2790_6);

wire[3:0] wires_2791_6;

wire[31:0] addr_2791_6;

Selector_2 s2791_6(wires_697_5[3], addr_697_5, wires_2791_6,addr_2791_6);

wire[3:0] wires_2792_6;

wire[31:0] addr_2792_6;

Selector_2 s2792_6(wires_698_5[0], addr_698_5, wires_2792_6,addr_2792_6);

wire[3:0] wires_2793_6;

wire[31:0] addr_2793_6;

Selector_2 s2793_6(wires_698_5[1], addr_698_5, wires_2793_6,addr_2793_6);

wire[3:0] wires_2794_6;

wire[31:0] addr_2794_6;

Selector_2 s2794_6(wires_698_5[2], addr_698_5, wires_2794_6,addr_2794_6);

wire[3:0] wires_2795_6;

wire[31:0] addr_2795_6;

Selector_2 s2795_6(wires_698_5[3], addr_698_5, wires_2795_6,addr_2795_6);

wire[3:0] wires_2796_6;

wire[31:0] addr_2796_6;

Selector_2 s2796_6(wires_699_5[0], addr_699_5, wires_2796_6,addr_2796_6);

wire[3:0] wires_2797_6;

wire[31:0] addr_2797_6;

Selector_2 s2797_6(wires_699_5[1], addr_699_5, wires_2797_6,addr_2797_6);

wire[3:0] wires_2798_6;

wire[31:0] addr_2798_6;

Selector_2 s2798_6(wires_699_5[2], addr_699_5, wires_2798_6,addr_2798_6);

wire[3:0] wires_2799_6;

wire[31:0] addr_2799_6;

Selector_2 s2799_6(wires_699_5[3], addr_699_5, wires_2799_6,addr_2799_6);

wire[3:0] wires_2800_6;

wire[31:0] addr_2800_6;

Selector_2 s2800_6(wires_700_5[0], addr_700_5, wires_2800_6,addr_2800_6);

wire[3:0] wires_2801_6;

wire[31:0] addr_2801_6;

Selector_2 s2801_6(wires_700_5[1], addr_700_5, wires_2801_6,addr_2801_6);

wire[3:0] wires_2802_6;

wire[31:0] addr_2802_6;

Selector_2 s2802_6(wires_700_5[2], addr_700_5, wires_2802_6,addr_2802_6);

wire[3:0] wires_2803_6;

wire[31:0] addr_2803_6;

Selector_2 s2803_6(wires_700_5[3], addr_700_5, wires_2803_6,addr_2803_6);

wire[3:0] wires_2804_6;

wire[31:0] addr_2804_6;

Selector_2 s2804_6(wires_701_5[0], addr_701_5, wires_2804_6,addr_2804_6);

wire[3:0] wires_2805_6;

wire[31:0] addr_2805_6;

Selector_2 s2805_6(wires_701_5[1], addr_701_5, wires_2805_6,addr_2805_6);

wire[3:0] wires_2806_6;

wire[31:0] addr_2806_6;

Selector_2 s2806_6(wires_701_5[2], addr_701_5, wires_2806_6,addr_2806_6);

wire[3:0] wires_2807_6;

wire[31:0] addr_2807_6;

Selector_2 s2807_6(wires_701_5[3], addr_701_5, wires_2807_6,addr_2807_6);

wire[3:0] wires_2808_6;

wire[31:0] addr_2808_6;

Selector_2 s2808_6(wires_702_5[0], addr_702_5, wires_2808_6,addr_2808_6);

wire[3:0] wires_2809_6;

wire[31:0] addr_2809_6;

Selector_2 s2809_6(wires_702_5[1], addr_702_5, wires_2809_6,addr_2809_6);

wire[3:0] wires_2810_6;

wire[31:0] addr_2810_6;

Selector_2 s2810_6(wires_702_5[2], addr_702_5, wires_2810_6,addr_2810_6);

wire[3:0] wires_2811_6;

wire[31:0] addr_2811_6;

Selector_2 s2811_6(wires_702_5[3], addr_702_5, wires_2811_6,addr_2811_6);

wire[3:0] wires_2812_6;

wire[31:0] addr_2812_6;

Selector_2 s2812_6(wires_703_5[0], addr_703_5, wires_2812_6,addr_2812_6);

wire[3:0] wires_2813_6;

wire[31:0] addr_2813_6;

Selector_2 s2813_6(wires_703_5[1], addr_703_5, wires_2813_6,addr_2813_6);

wire[3:0] wires_2814_6;

wire[31:0] addr_2814_6;

Selector_2 s2814_6(wires_703_5[2], addr_703_5, wires_2814_6,addr_2814_6);

wire[3:0] wires_2815_6;

wire[31:0] addr_2815_6;

Selector_2 s2815_6(wires_703_5[3], addr_703_5, wires_2815_6,addr_2815_6);

wire[3:0] wires_2816_6;

wire[31:0] addr_2816_6;

Selector_2 s2816_6(wires_704_5[0], addr_704_5, wires_2816_6,addr_2816_6);

wire[3:0] wires_2817_6;

wire[31:0] addr_2817_6;

Selector_2 s2817_6(wires_704_5[1], addr_704_5, wires_2817_6,addr_2817_6);

wire[3:0] wires_2818_6;

wire[31:0] addr_2818_6;

Selector_2 s2818_6(wires_704_5[2], addr_704_5, wires_2818_6,addr_2818_6);

wire[3:0] wires_2819_6;

wire[31:0] addr_2819_6;

Selector_2 s2819_6(wires_704_5[3], addr_704_5, wires_2819_6,addr_2819_6);

wire[3:0] wires_2820_6;

wire[31:0] addr_2820_6;

Selector_2 s2820_6(wires_705_5[0], addr_705_5, wires_2820_6,addr_2820_6);

wire[3:0] wires_2821_6;

wire[31:0] addr_2821_6;

Selector_2 s2821_6(wires_705_5[1], addr_705_5, wires_2821_6,addr_2821_6);

wire[3:0] wires_2822_6;

wire[31:0] addr_2822_6;

Selector_2 s2822_6(wires_705_5[2], addr_705_5, wires_2822_6,addr_2822_6);

wire[3:0] wires_2823_6;

wire[31:0] addr_2823_6;

Selector_2 s2823_6(wires_705_5[3], addr_705_5, wires_2823_6,addr_2823_6);

wire[3:0] wires_2824_6;

wire[31:0] addr_2824_6;

Selector_2 s2824_6(wires_706_5[0], addr_706_5, wires_2824_6,addr_2824_6);

wire[3:0] wires_2825_6;

wire[31:0] addr_2825_6;

Selector_2 s2825_6(wires_706_5[1], addr_706_5, wires_2825_6,addr_2825_6);

wire[3:0] wires_2826_6;

wire[31:0] addr_2826_6;

Selector_2 s2826_6(wires_706_5[2], addr_706_5, wires_2826_6,addr_2826_6);

wire[3:0] wires_2827_6;

wire[31:0] addr_2827_6;

Selector_2 s2827_6(wires_706_5[3], addr_706_5, wires_2827_6,addr_2827_6);

wire[3:0] wires_2828_6;

wire[31:0] addr_2828_6;

Selector_2 s2828_6(wires_707_5[0], addr_707_5, wires_2828_6,addr_2828_6);

wire[3:0] wires_2829_6;

wire[31:0] addr_2829_6;

Selector_2 s2829_6(wires_707_5[1], addr_707_5, wires_2829_6,addr_2829_6);

wire[3:0] wires_2830_6;

wire[31:0] addr_2830_6;

Selector_2 s2830_6(wires_707_5[2], addr_707_5, wires_2830_6,addr_2830_6);

wire[3:0] wires_2831_6;

wire[31:0] addr_2831_6;

Selector_2 s2831_6(wires_707_5[3], addr_707_5, wires_2831_6,addr_2831_6);

wire[3:0] wires_2832_6;

wire[31:0] addr_2832_6;

Selector_2 s2832_6(wires_708_5[0], addr_708_5, wires_2832_6,addr_2832_6);

wire[3:0] wires_2833_6;

wire[31:0] addr_2833_6;

Selector_2 s2833_6(wires_708_5[1], addr_708_5, wires_2833_6,addr_2833_6);

wire[3:0] wires_2834_6;

wire[31:0] addr_2834_6;

Selector_2 s2834_6(wires_708_5[2], addr_708_5, wires_2834_6,addr_2834_6);

wire[3:0] wires_2835_6;

wire[31:0] addr_2835_6;

Selector_2 s2835_6(wires_708_5[3], addr_708_5, wires_2835_6,addr_2835_6);

wire[3:0] wires_2836_6;

wire[31:0] addr_2836_6;

Selector_2 s2836_6(wires_709_5[0], addr_709_5, wires_2836_6,addr_2836_6);

wire[3:0] wires_2837_6;

wire[31:0] addr_2837_6;

Selector_2 s2837_6(wires_709_5[1], addr_709_5, wires_2837_6,addr_2837_6);

wire[3:0] wires_2838_6;

wire[31:0] addr_2838_6;

Selector_2 s2838_6(wires_709_5[2], addr_709_5, wires_2838_6,addr_2838_6);

wire[3:0] wires_2839_6;

wire[31:0] addr_2839_6;

Selector_2 s2839_6(wires_709_5[3], addr_709_5, wires_2839_6,addr_2839_6);

wire[3:0] wires_2840_6;

wire[31:0] addr_2840_6;

Selector_2 s2840_6(wires_710_5[0], addr_710_5, wires_2840_6,addr_2840_6);

wire[3:0] wires_2841_6;

wire[31:0] addr_2841_6;

Selector_2 s2841_6(wires_710_5[1], addr_710_5, wires_2841_6,addr_2841_6);

wire[3:0] wires_2842_6;

wire[31:0] addr_2842_6;

Selector_2 s2842_6(wires_710_5[2], addr_710_5, wires_2842_6,addr_2842_6);

wire[3:0] wires_2843_6;

wire[31:0] addr_2843_6;

Selector_2 s2843_6(wires_710_5[3], addr_710_5, wires_2843_6,addr_2843_6);

wire[3:0] wires_2844_6;

wire[31:0] addr_2844_6;

Selector_2 s2844_6(wires_711_5[0], addr_711_5, wires_2844_6,addr_2844_6);

wire[3:0] wires_2845_6;

wire[31:0] addr_2845_6;

Selector_2 s2845_6(wires_711_5[1], addr_711_5, wires_2845_6,addr_2845_6);

wire[3:0] wires_2846_6;

wire[31:0] addr_2846_6;

Selector_2 s2846_6(wires_711_5[2], addr_711_5, wires_2846_6,addr_2846_6);

wire[3:0] wires_2847_6;

wire[31:0] addr_2847_6;

Selector_2 s2847_6(wires_711_5[3], addr_711_5, wires_2847_6,addr_2847_6);

wire[3:0] wires_2848_6;

wire[31:0] addr_2848_6;

Selector_2 s2848_6(wires_712_5[0], addr_712_5, wires_2848_6,addr_2848_6);

wire[3:0] wires_2849_6;

wire[31:0] addr_2849_6;

Selector_2 s2849_6(wires_712_5[1], addr_712_5, wires_2849_6,addr_2849_6);

wire[3:0] wires_2850_6;

wire[31:0] addr_2850_6;

Selector_2 s2850_6(wires_712_5[2], addr_712_5, wires_2850_6,addr_2850_6);

wire[3:0] wires_2851_6;

wire[31:0] addr_2851_6;

Selector_2 s2851_6(wires_712_5[3], addr_712_5, wires_2851_6,addr_2851_6);

wire[3:0] wires_2852_6;

wire[31:0] addr_2852_6;

Selector_2 s2852_6(wires_713_5[0], addr_713_5, wires_2852_6,addr_2852_6);

wire[3:0] wires_2853_6;

wire[31:0] addr_2853_6;

Selector_2 s2853_6(wires_713_5[1], addr_713_5, wires_2853_6,addr_2853_6);

wire[3:0] wires_2854_6;

wire[31:0] addr_2854_6;

Selector_2 s2854_6(wires_713_5[2], addr_713_5, wires_2854_6,addr_2854_6);

wire[3:0] wires_2855_6;

wire[31:0] addr_2855_6;

Selector_2 s2855_6(wires_713_5[3], addr_713_5, wires_2855_6,addr_2855_6);

wire[3:0] wires_2856_6;

wire[31:0] addr_2856_6;

Selector_2 s2856_6(wires_714_5[0], addr_714_5, wires_2856_6,addr_2856_6);

wire[3:0] wires_2857_6;

wire[31:0] addr_2857_6;

Selector_2 s2857_6(wires_714_5[1], addr_714_5, wires_2857_6,addr_2857_6);

wire[3:0] wires_2858_6;

wire[31:0] addr_2858_6;

Selector_2 s2858_6(wires_714_5[2], addr_714_5, wires_2858_6,addr_2858_6);

wire[3:0] wires_2859_6;

wire[31:0] addr_2859_6;

Selector_2 s2859_6(wires_714_5[3], addr_714_5, wires_2859_6,addr_2859_6);

wire[3:0] wires_2860_6;

wire[31:0] addr_2860_6;

Selector_2 s2860_6(wires_715_5[0], addr_715_5, wires_2860_6,addr_2860_6);

wire[3:0] wires_2861_6;

wire[31:0] addr_2861_6;

Selector_2 s2861_6(wires_715_5[1], addr_715_5, wires_2861_6,addr_2861_6);

wire[3:0] wires_2862_6;

wire[31:0] addr_2862_6;

Selector_2 s2862_6(wires_715_5[2], addr_715_5, wires_2862_6,addr_2862_6);

wire[3:0] wires_2863_6;

wire[31:0] addr_2863_6;

Selector_2 s2863_6(wires_715_5[3], addr_715_5, wires_2863_6,addr_2863_6);

wire[3:0] wires_2864_6;

wire[31:0] addr_2864_6;

Selector_2 s2864_6(wires_716_5[0], addr_716_5, wires_2864_6,addr_2864_6);

wire[3:0] wires_2865_6;

wire[31:0] addr_2865_6;

Selector_2 s2865_6(wires_716_5[1], addr_716_5, wires_2865_6,addr_2865_6);

wire[3:0] wires_2866_6;

wire[31:0] addr_2866_6;

Selector_2 s2866_6(wires_716_5[2], addr_716_5, wires_2866_6,addr_2866_6);

wire[3:0] wires_2867_6;

wire[31:0] addr_2867_6;

Selector_2 s2867_6(wires_716_5[3], addr_716_5, wires_2867_6,addr_2867_6);

wire[3:0] wires_2868_6;

wire[31:0] addr_2868_6;

Selector_2 s2868_6(wires_717_5[0], addr_717_5, wires_2868_6,addr_2868_6);

wire[3:0] wires_2869_6;

wire[31:0] addr_2869_6;

Selector_2 s2869_6(wires_717_5[1], addr_717_5, wires_2869_6,addr_2869_6);

wire[3:0] wires_2870_6;

wire[31:0] addr_2870_6;

Selector_2 s2870_6(wires_717_5[2], addr_717_5, wires_2870_6,addr_2870_6);

wire[3:0] wires_2871_6;

wire[31:0] addr_2871_6;

Selector_2 s2871_6(wires_717_5[3], addr_717_5, wires_2871_6,addr_2871_6);

wire[3:0] wires_2872_6;

wire[31:0] addr_2872_6;

Selector_2 s2872_6(wires_718_5[0], addr_718_5, wires_2872_6,addr_2872_6);

wire[3:0] wires_2873_6;

wire[31:0] addr_2873_6;

Selector_2 s2873_6(wires_718_5[1], addr_718_5, wires_2873_6,addr_2873_6);

wire[3:0] wires_2874_6;

wire[31:0] addr_2874_6;

Selector_2 s2874_6(wires_718_5[2], addr_718_5, wires_2874_6,addr_2874_6);

wire[3:0] wires_2875_6;

wire[31:0] addr_2875_6;

Selector_2 s2875_6(wires_718_5[3], addr_718_5, wires_2875_6,addr_2875_6);

wire[3:0] wires_2876_6;

wire[31:0] addr_2876_6;

Selector_2 s2876_6(wires_719_5[0], addr_719_5, wires_2876_6,addr_2876_6);

wire[3:0] wires_2877_6;

wire[31:0] addr_2877_6;

Selector_2 s2877_6(wires_719_5[1], addr_719_5, wires_2877_6,addr_2877_6);

wire[3:0] wires_2878_6;

wire[31:0] addr_2878_6;

Selector_2 s2878_6(wires_719_5[2], addr_719_5, wires_2878_6,addr_2878_6);

wire[3:0] wires_2879_6;

wire[31:0] addr_2879_6;

Selector_2 s2879_6(wires_719_5[3], addr_719_5, wires_2879_6,addr_2879_6);

wire[3:0] wires_2880_6;

wire[31:0] addr_2880_6;

Selector_2 s2880_6(wires_720_5[0], addr_720_5, wires_2880_6,addr_2880_6);

wire[3:0] wires_2881_6;

wire[31:0] addr_2881_6;

Selector_2 s2881_6(wires_720_5[1], addr_720_5, wires_2881_6,addr_2881_6);

wire[3:0] wires_2882_6;

wire[31:0] addr_2882_6;

Selector_2 s2882_6(wires_720_5[2], addr_720_5, wires_2882_6,addr_2882_6);

wire[3:0] wires_2883_6;

wire[31:0] addr_2883_6;

Selector_2 s2883_6(wires_720_5[3], addr_720_5, wires_2883_6,addr_2883_6);

wire[3:0] wires_2884_6;

wire[31:0] addr_2884_6;

Selector_2 s2884_6(wires_721_5[0], addr_721_5, wires_2884_6,addr_2884_6);

wire[3:0] wires_2885_6;

wire[31:0] addr_2885_6;

Selector_2 s2885_6(wires_721_5[1], addr_721_5, wires_2885_6,addr_2885_6);

wire[3:0] wires_2886_6;

wire[31:0] addr_2886_6;

Selector_2 s2886_6(wires_721_5[2], addr_721_5, wires_2886_6,addr_2886_6);

wire[3:0] wires_2887_6;

wire[31:0] addr_2887_6;

Selector_2 s2887_6(wires_721_5[3], addr_721_5, wires_2887_6,addr_2887_6);

wire[3:0] wires_2888_6;

wire[31:0] addr_2888_6;

Selector_2 s2888_6(wires_722_5[0], addr_722_5, wires_2888_6,addr_2888_6);

wire[3:0] wires_2889_6;

wire[31:0] addr_2889_6;

Selector_2 s2889_6(wires_722_5[1], addr_722_5, wires_2889_6,addr_2889_6);

wire[3:0] wires_2890_6;

wire[31:0] addr_2890_6;

Selector_2 s2890_6(wires_722_5[2], addr_722_5, wires_2890_6,addr_2890_6);

wire[3:0] wires_2891_6;

wire[31:0] addr_2891_6;

Selector_2 s2891_6(wires_722_5[3], addr_722_5, wires_2891_6,addr_2891_6);

wire[3:0] wires_2892_6;

wire[31:0] addr_2892_6;

Selector_2 s2892_6(wires_723_5[0], addr_723_5, wires_2892_6,addr_2892_6);

wire[3:0] wires_2893_6;

wire[31:0] addr_2893_6;

Selector_2 s2893_6(wires_723_5[1], addr_723_5, wires_2893_6,addr_2893_6);

wire[3:0] wires_2894_6;

wire[31:0] addr_2894_6;

Selector_2 s2894_6(wires_723_5[2], addr_723_5, wires_2894_6,addr_2894_6);

wire[3:0] wires_2895_6;

wire[31:0] addr_2895_6;

Selector_2 s2895_6(wires_723_5[3], addr_723_5, wires_2895_6,addr_2895_6);

wire[3:0] wires_2896_6;

wire[31:0] addr_2896_6;

Selector_2 s2896_6(wires_724_5[0], addr_724_5, wires_2896_6,addr_2896_6);

wire[3:0] wires_2897_6;

wire[31:0] addr_2897_6;

Selector_2 s2897_6(wires_724_5[1], addr_724_5, wires_2897_6,addr_2897_6);

wire[3:0] wires_2898_6;

wire[31:0] addr_2898_6;

Selector_2 s2898_6(wires_724_5[2], addr_724_5, wires_2898_6,addr_2898_6);

wire[3:0] wires_2899_6;

wire[31:0] addr_2899_6;

Selector_2 s2899_6(wires_724_5[3], addr_724_5, wires_2899_6,addr_2899_6);

wire[3:0] wires_2900_6;

wire[31:0] addr_2900_6;

Selector_2 s2900_6(wires_725_5[0], addr_725_5, wires_2900_6,addr_2900_6);

wire[3:0] wires_2901_6;

wire[31:0] addr_2901_6;

Selector_2 s2901_6(wires_725_5[1], addr_725_5, wires_2901_6,addr_2901_6);

wire[3:0] wires_2902_6;

wire[31:0] addr_2902_6;

Selector_2 s2902_6(wires_725_5[2], addr_725_5, wires_2902_6,addr_2902_6);

wire[3:0] wires_2903_6;

wire[31:0] addr_2903_6;

Selector_2 s2903_6(wires_725_5[3], addr_725_5, wires_2903_6,addr_2903_6);

wire[3:0] wires_2904_6;

wire[31:0] addr_2904_6;

Selector_2 s2904_6(wires_726_5[0], addr_726_5, wires_2904_6,addr_2904_6);

wire[3:0] wires_2905_6;

wire[31:0] addr_2905_6;

Selector_2 s2905_6(wires_726_5[1], addr_726_5, wires_2905_6,addr_2905_6);

wire[3:0] wires_2906_6;

wire[31:0] addr_2906_6;

Selector_2 s2906_6(wires_726_5[2], addr_726_5, wires_2906_6,addr_2906_6);

wire[3:0] wires_2907_6;

wire[31:0] addr_2907_6;

Selector_2 s2907_6(wires_726_5[3], addr_726_5, wires_2907_6,addr_2907_6);

wire[3:0] wires_2908_6;

wire[31:0] addr_2908_6;

Selector_2 s2908_6(wires_727_5[0], addr_727_5, wires_2908_6,addr_2908_6);

wire[3:0] wires_2909_6;

wire[31:0] addr_2909_6;

Selector_2 s2909_6(wires_727_5[1], addr_727_5, wires_2909_6,addr_2909_6);

wire[3:0] wires_2910_6;

wire[31:0] addr_2910_6;

Selector_2 s2910_6(wires_727_5[2], addr_727_5, wires_2910_6,addr_2910_6);

wire[3:0] wires_2911_6;

wire[31:0] addr_2911_6;

Selector_2 s2911_6(wires_727_5[3], addr_727_5, wires_2911_6,addr_2911_6);

wire[3:0] wires_2912_6;

wire[31:0] addr_2912_6;

Selector_2 s2912_6(wires_728_5[0], addr_728_5, wires_2912_6,addr_2912_6);

wire[3:0] wires_2913_6;

wire[31:0] addr_2913_6;

Selector_2 s2913_6(wires_728_5[1], addr_728_5, wires_2913_6,addr_2913_6);

wire[3:0] wires_2914_6;

wire[31:0] addr_2914_6;

Selector_2 s2914_6(wires_728_5[2], addr_728_5, wires_2914_6,addr_2914_6);

wire[3:0] wires_2915_6;

wire[31:0] addr_2915_6;

Selector_2 s2915_6(wires_728_5[3], addr_728_5, wires_2915_6,addr_2915_6);

wire[3:0] wires_2916_6;

wire[31:0] addr_2916_6;

Selector_2 s2916_6(wires_729_5[0], addr_729_5, wires_2916_6,addr_2916_6);

wire[3:0] wires_2917_6;

wire[31:0] addr_2917_6;

Selector_2 s2917_6(wires_729_5[1], addr_729_5, wires_2917_6,addr_2917_6);

wire[3:0] wires_2918_6;

wire[31:0] addr_2918_6;

Selector_2 s2918_6(wires_729_5[2], addr_729_5, wires_2918_6,addr_2918_6);

wire[3:0] wires_2919_6;

wire[31:0] addr_2919_6;

Selector_2 s2919_6(wires_729_5[3], addr_729_5, wires_2919_6,addr_2919_6);

wire[3:0] wires_2920_6;

wire[31:0] addr_2920_6;

Selector_2 s2920_6(wires_730_5[0], addr_730_5, wires_2920_6,addr_2920_6);

wire[3:0] wires_2921_6;

wire[31:0] addr_2921_6;

Selector_2 s2921_6(wires_730_5[1], addr_730_5, wires_2921_6,addr_2921_6);

wire[3:0] wires_2922_6;

wire[31:0] addr_2922_6;

Selector_2 s2922_6(wires_730_5[2], addr_730_5, wires_2922_6,addr_2922_6);

wire[3:0] wires_2923_6;

wire[31:0] addr_2923_6;

Selector_2 s2923_6(wires_730_5[3], addr_730_5, wires_2923_6,addr_2923_6);

wire[3:0] wires_2924_6;

wire[31:0] addr_2924_6;

Selector_2 s2924_6(wires_731_5[0], addr_731_5, wires_2924_6,addr_2924_6);

wire[3:0] wires_2925_6;

wire[31:0] addr_2925_6;

Selector_2 s2925_6(wires_731_5[1], addr_731_5, wires_2925_6,addr_2925_6);

wire[3:0] wires_2926_6;

wire[31:0] addr_2926_6;

Selector_2 s2926_6(wires_731_5[2], addr_731_5, wires_2926_6,addr_2926_6);

wire[3:0] wires_2927_6;

wire[31:0] addr_2927_6;

Selector_2 s2927_6(wires_731_5[3], addr_731_5, wires_2927_6,addr_2927_6);

wire[3:0] wires_2928_6;

wire[31:0] addr_2928_6;

Selector_2 s2928_6(wires_732_5[0], addr_732_5, wires_2928_6,addr_2928_6);

wire[3:0] wires_2929_6;

wire[31:0] addr_2929_6;

Selector_2 s2929_6(wires_732_5[1], addr_732_5, wires_2929_6,addr_2929_6);

wire[3:0] wires_2930_6;

wire[31:0] addr_2930_6;

Selector_2 s2930_6(wires_732_5[2], addr_732_5, wires_2930_6,addr_2930_6);

wire[3:0] wires_2931_6;

wire[31:0] addr_2931_6;

Selector_2 s2931_6(wires_732_5[3], addr_732_5, wires_2931_6,addr_2931_6);

wire[3:0] wires_2932_6;

wire[31:0] addr_2932_6;

Selector_2 s2932_6(wires_733_5[0], addr_733_5, wires_2932_6,addr_2932_6);

wire[3:0] wires_2933_6;

wire[31:0] addr_2933_6;

Selector_2 s2933_6(wires_733_5[1], addr_733_5, wires_2933_6,addr_2933_6);

wire[3:0] wires_2934_6;

wire[31:0] addr_2934_6;

Selector_2 s2934_6(wires_733_5[2], addr_733_5, wires_2934_6,addr_2934_6);

wire[3:0] wires_2935_6;

wire[31:0] addr_2935_6;

Selector_2 s2935_6(wires_733_5[3], addr_733_5, wires_2935_6,addr_2935_6);

wire[3:0] wires_2936_6;

wire[31:0] addr_2936_6;

Selector_2 s2936_6(wires_734_5[0], addr_734_5, wires_2936_6,addr_2936_6);

wire[3:0] wires_2937_6;

wire[31:0] addr_2937_6;

Selector_2 s2937_6(wires_734_5[1], addr_734_5, wires_2937_6,addr_2937_6);

wire[3:0] wires_2938_6;

wire[31:0] addr_2938_6;

Selector_2 s2938_6(wires_734_5[2], addr_734_5, wires_2938_6,addr_2938_6);

wire[3:0] wires_2939_6;

wire[31:0] addr_2939_6;

Selector_2 s2939_6(wires_734_5[3], addr_734_5, wires_2939_6,addr_2939_6);

wire[3:0] wires_2940_6;

wire[31:0] addr_2940_6;

Selector_2 s2940_6(wires_735_5[0], addr_735_5, wires_2940_6,addr_2940_6);

wire[3:0] wires_2941_6;

wire[31:0] addr_2941_6;

Selector_2 s2941_6(wires_735_5[1], addr_735_5, wires_2941_6,addr_2941_6);

wire[3:0] wires_2942_6;

wire[31:0] addr_2942_6;

Selector_2 s2942_6(wires_735_5[2], addr_735_5, wires_2942_6,addr_2942_6);

wire[3:0] wires_2943_6;

wire[31:0] addr_2943_6;

Selector_2 s2943_6(wires_735_5[3], addr_735_5, wires_2943_6,addr_2943_6);

wire[3:0] wires_2944_6;

wire[31:0] addr_2944_6;

Selector_2 s2944_6(wires_736_5[0], addr_736_5, wires_2944_6,addr_2944_6);

wire[3:0] wires_2945_6;

wire[31:0] addr_2945_6;

Selector_2 s2945_6(wires_736_5[1], addr_736_5, wires_2945_6,addr_2945_6);

wire[3:0] wires_2946_6;

wire[31:0] addr_2946_6;

Selector_2 s2946_6(wires_736_5[2], addr_736_5, wires_2946_6,addr_2946_6);

wire[3:0] wires_2947_6;

wire[31:0] addr_2947_6;

Selector_2 s2947_6(wires_736_5[3], addr_736_5, wires_2947_6,addr_2947_6);

wire[3:0] wires_2948_6;

wire[31:0] addr_2948_6;

Selector_2 s2948_6(wires_737_5[0], addr_737_5, wires_2948_6,addr_2948_6);

wire[3:0] wires_2949_6;

wire[31:0] addr_2949_6;

Selector_2 s2949_6(wires_737_5[1], addr_737_5, wires_2949_6,addr_2949_6);

wire[3:0] wires_2950_6;

wire[31:0] addr_2950_6;

Selector_2 s2950_6(wires_737_5[2], addr_737_5, wires_2950_6,addr_2950_6);

wire[3:0] wires_2951_6;

wire[31:0] addr_2951_6;

Selector_2 s2951_6(wires_737_5[3], addr_737_5, wires_2951_6,addr_2951_6);

wire[3:0] wires_2952_6;

wire[31:0] addr_2952_6;

Selector_2 s2952_6(wires_738_5[0], addr_738_5, wires_2952_6,addr_2952_6);

wire[3:0] wires_2953_6;

wire[31:0] addr_2953_6;

Selector_2 s2953_6(wires_738_5[1], addr_738_5, wires_2953_6,addr_2953_6);

wire[3:0] wires_2954_6;

wire[31:0] addr_2954_6;

Selector_2 s2954_6(wires_738_5[2], addr_738_5, wires_2954_6,addr_2954_6);

wire[3:0] wires_2955_6;

wire[31:0] addr_2955_6;

Selector_2 s2955_6(wires_738_5[3], addr_738_5, wires_2955_6,addr_2955_6);

wire[3:0] wires_2956_6;

wire[31:0] addr_2956_6;

Selector_2 s2956_6(wires_739_5[0], addr_739_5, wires_2956_6,addr_2956_6);

wire[3:0] wires_2957_6;

wire[31:0] addr_2957_6;

Selector_2 s2957_6(wires_739_5[1], addr_739_5, wires_2957_6,addr_2957_6);

wire[3:0] wires_2958_6;

wire[31:0] addr_2958_6;

Selector_2 s2958_6(wires_739_5[2], addr_739_5, wires_2958_6,addr_2958_6);

wire[3:0] wires_2959_6;

wire[31:0] addr_2959_6;

Selector_2 s2959_6(wires_739_5[3], addr_739_5, wires_2959_6,addr_2959_6);

wire[3:0] wires_2960_6;

wire[31:0] addr_2960_6;

Selector_2 s2960_6(wires_740_5[0], addr_740_5, wires_2960_6,addr_2960_6);

wire[3:0] wires_2961_6;

wire[31:0] addr_2961_6;

Selector_2 s2961_6(wires_740_5[1], addr_740_5, wires_2961_6,addr_2961_6);

wire[3:0] wires_2962_6;

wire[31:0] addr_2962_6;

Selector_2 s2962_6(wires_740_5[2], addr_740_5, wires_2962_6,addr_2962_6);

wire[3:0] wires_2963_6;

wire[31:0] addr_2963_6;

Selector_2 s2963_6(wires_740_5[3], addr_740_5, wires_2963_6,addr_2963_6);

wire[3:0] wires_2964_6;

wire[31:0] addr_2964_6;

Selector_2 s2964_6(wires_741_5[0], addr_741_5, wires_2964_6,addr_2964_6);

wire[3:0] wires_2965_6;

wire[31:0] addr_2965_6;

Selector_2 s2965_6(wires_741_5[1], addr_741_5, wires_2965_6,addr_2965_6);

wire[3:0] wires_2966_6;

wire[31:0] addr_2966_6;

Selector_2 s2966_6(wires_741_5[2], addr_741_5, wires_2966_6,addr_2966_6);

wire[3:0] wires_2967_6;

wire[31:0] addr_2967_6;

Selector_2 s2967_6(wires_741_5[3], addr_741_5, wires_2967_6,addr_2967_6);

wire[3:0] wires_2968_6;

wire[31:0] addr_2968_6;

Selector_2 s2968_6(wires_742_5[0], addr_742_5, wires_2968_6,addr_2968_6);

wire[3:0] wires_2969_6;

wire[31:0] addr_2969_6;

Selector_2 s2969_6(wires_742_5[1], addr_742_5, wires_2969_6,addr_2969_6);

wire[3:0] wires_2970_6;

wire[31:0] addr_2970_6;

Selector_2 s2970_6(wires_742_5[2], addr_742_5, wires_2970_6,addr_2970_6);

wire[3:0] wires_2971_6;

wire[31:0] addr_2971_6;

Selector_2 s2971_6(wires_742_5[3], addr_742_5, wires_2971_6,addr_2971_6);

wire[3:0] wires_2972_6;

wire[31:0] addr_2972_6;

Selector_2 s2972_6(wires_743_5[0], addr_743_5, wires_2972_6,addr_2972_6);

wire[3:0] wires_2973_6;

wire[31:0] addr_2973_6;

Selector_2 s2973_6(wires_743_5[1], addr_743_5, wires_2973_6,addr_2973_6);

wire[3:0] wires_2974_6;

wire[31:0] addr_2974_6;

Selector_2 s2974_6(wires_743_5[2], addr_743_5, wires_2974_6,addr_2974_6);

wire[3:0] wires_2975_6;

wire[31:0] addr_2975_6;

Selector_2 s2975_6(wires_743_5[3], addr_743_5, wires_2975_6,addr_2975_6);

wire[3:0] wires_2976_6;

wire[31:0] addr_2976_6;

Selector_2 s2976_6(wires_744_5[0], addr_744_5, wires_2976_6,addr_2976_6);

wire[3:0] wires_2977_6;

wire[31:0] addr_2977_6;

Selector_2 s2977_6(wires_744_5[1], addr_744_5, wires_2977_6,addr_2977_6);

wire[3:0] wires_2978_6;

wire[31:0] addr_2978_6;

Selector_2 s2978_6(wires_744_5[2], addr_744_5, wires_2978_6,addr_2978_6);

wire[3:0] wires_2979_6;

wire[31:0] addr_2979_6;

Selector_2 s2979_6(wires_744_5[3], addr_744_5, wires_2979_6,addr_2979_6);

wire[3:0] wires_2980_6;

wire[31:0] addr_2980_6;

Selector_2 s2980_6(wires_745_5[0], addr_745_5, wires_2980_6,addr_2980_6);

wire[3:0] wires_2981_6;

wire[31:0] addr_2981_6;

Selector_2 s2981_6(wires_745_5[1], addr_745_5, wires_2981_6,addr_2981_6);

wire[3:0] wires_2982_6;

wire[31:0] addr_2982_6;

Selector_2 s2982_6(wires_745_5[2], addr_745_5, wires_2982_6,addr_2982_6);

wire[3:0] wires_2983_6;

wire[31:0] addr_2983_6;

Selector_2 s2983_6(wires_745_5[3], addr_745_5, wires_2983_6,addr_2983_6);

wire[3:0] wires_2984_6;

wire[31:0] addr_2984_6;

Selector_2 s2984_6(wires_746_5[0], addr_746_5, wires_2984_6,addr_2984_6);

wire[3:0] wires_2985_6;

wire[31:0] addr_2985_6;

Selector_2 s2985_6(wires_746_5[1], addr_746_5, wires_2985_6,addr_2985_6);

wire[3:0] wires_2986_6;

wire[31:0] addr_2986_6;

Selector_2 s2986_6(wires_746_5[2], addr_746_5, wires_2986_6,addr_2986_6);

wire[3:0] wires_2987_6;

wire[31:0] addr_2987_6;

Selector_2 s2987_6(wires_746_5[3], addr_746_5, wires_2987_6,addr_2987_6);

wire[3:0] wires_2988_6;

wire[31:0] addr_2988_6;

Selector_2 s2988_6(wires_747_5[0], addr_747_5, wires_2988_6,addr_2988_6);

wire[3:0] wires_2989_6;

wire[31:0] addr_2989_6;

Selector_2 s2989_6(wires_747_5[1], addr_747_5, wires_2989_6,addr_2989_6);

wire[3:0] wires_2990_6;

wire[31:0] addr_2990_6;

Selector_2 s2990_6(wires_747_5[2], addr_747_5, wires_2990_6,addr_2990_6);

wire[3:0] wires_2991_6;

wire[31:0] addr_2991_6;

Selector_2 s2991_6(wires_747_5[3], addr_747_5, wires_2991_6,addr_2991_6);

wire[3:0] wires_2992_6;

wire[31:0] addr_2992_6;

Selector_2 s2992_6(wires_748_5[0], addr_748_5, wires_2992_6,addr_2992_6);

wire[3:0] wires_2993_6;

wire[31:0] addr_2993_6;

Selector_2 s2993_6(wires_748_5[1], addr_748_5, wires_2993_6,addr_2993_6);

wire[3:0] wires_2994_6;

wire[31:0] addr_2994_6;

Selector_2 s2994_6(wires_748_5[2], addr_748_5, wires_2994_6,addr_2994_6);

wire[3:0] wires_2995_6;

wire[31:0] addr_2995_6;

Selector_2 s2995_6(wires_748_5[3], addr_748_5, wires_2995_6,addr_2995_6);

wire[3:0] wires_2996_6;

wire[31:0] addr_2996_6;

Selector_2 s2996_6(wires_749_5[0], addr_749_5, wires_2996_6,addr_2996_6);

wire[3:0] wires_2997_6;

wire[31:0] addr_2997_6;

Selector_2 s2997_6(wires_749_5[1], addr_749_5, wires_2997_6,addr_2997_6);

wire[3:0] wires_2998_6;

wire[31:0] addr_2998_6;

Selector_2 s2998_6(wires_749_5[2], addr_749_5, wires_2998_6,addr_2998_6);

wire[3:0] wires_2999_6;

wire[31:0] addr_2999_6;

Selector_2 s2999_6(wires_749_5[3], addr_749_5, wires_2999_6,addr_2999_6);

wire[3:0] wires_3000_6;

wire[31:0] addr_3000_6;

Selector_2 s3000_6(wires_750_5[0], addr_750_5, wires_3000_6,addr_3000_6);

wire[3:0] wires_3001_6;

wire[31:0] addr_3001_6;

Selector_2 s3001_6(wires_750_5[1], addr_750_5, wires_3001_6,addr_3001_6);

wire[3:0] wires_3002_6;

wire[31:0] addr_3002_6;

Selector_2 s3002_6(wires_750_5[2], addr_750_5, wires_3002_6,addr_3002_6);

wire[3:0] wires_3003_6;

wire[31:0] addr_3003_6;

Selector_2 s3003_6(wires_750_5[3], addr_750_5, wires_3003_6,addr_3003_6);

wire[3:0] wires_3004_6;

wire[31:0] addr_3004_6;

Selector_2 s3004_6(wires_751_5[0], addr_751_5, wires_3004_6,addr_3004_6);

wire[3:0] wires_3005_6;

wire[31:0] addr_3005_6;

Selector_2 s3005_6(wires_751_5[1], addr_751_5, wires_3005_6,addr_3005_6);

wire[3:0] wires_3006_6;

wire[31:0] addr_3006_6;

Selector_2 s3006_6(wires_751_5[2], addr_751_5, wires_3006_6,addr_3006_6);

wire[3:0] wires_3007_6;

wire[31:0] addr_3007_6;

Selector_2 s3007_6(wires_751_5[3], addr_751_5, wires_3007_6,addr_3007_6);

wire[3:0] wires_3008_6;

wire[31:0] addr_3008_6;

Selector_2 s3008_6(wires_752_5[0], addr_752_5, wires_3008_6,addr_3008_6);

wire[3:0] wires_3009_6;

wire[31:0] addr_3009_6;

Selector_2 s3009_6(wires_752_5[1], addr_752_5, wires_3009_6,addr_3009_6);

wire[3:0] wires_3010_6;

wire[31:0] addr_3010_6;

Selector_2 s3010_6(wires_752_5[2], addr_752_5, wires_3010_6,addr_3010_6);

wire[3:0] wires_3011_6;

wire[31:0] addr_3011_6;

Selector_2 s3011_6(wires_752_5[3], addr_752_5, wires_3011_6,addr_3011_6);

wire[3:0] wires_3012_6;

wire[31:0] addr_3012_6;

Selector_2 s3012_6(wires_753_5[0], addr_753_5, wires_3012_6,addr_3012_6);

wire[3:0] wires_3013_6;

wire[31:0] addr_3013_6;

Selector_2 s3013_6(wires_753_5[1], addr_753_5, wires_3013_6,addr_3013_6);

wire[3:0] wires_3014_6;

wire[31:0] addr_3014_6;

Selector_2 s3014_6(wires_753_5[2], addr_753_5, wires_3014_6,addr_3014_6);

wire[3:0] wires_3015_6;

wire[31:0] addr_3015_6;

Selector_2 s3015_6(wires_753_5[3], addr_753_5, wires_3015_6,addr_3015_6);

wire[3:0] wires_3016_6;

wire[31:0] addr_3016_6;

Selector_2 s3016_6(wires_754_5[0], addr_754_5, wires_3016_6,addr_3016_6);

wire[3:0] wires_3017_6;

wire[31:0] addr_3017_6;

Selector_2 s3017_6(wires_754_5[1], addr_754_5, wires_3017_6,addr_3017_6);

wire[3:0] wires_3018_6;

wire[31:0] addr_3018_6;

Selector_2 s3018_6(wires_754_5[2], addr_754_5, wires_3018_6,addr_3018_6);

wire[3:0] wires_3019_6;

wire[31:0] addr_3019_6;

Selector_2 s3019_6(wires_754_5[3], addr_754_5, wires_3019_6,addr_3019_6);

wire[3:0] wires_3020_6;

wire[31:0] addr_3020_6;

Selector_2 s3020_6(wires_755_5[0], addr_755_5, wires_3020_6,addr_3020_6);

wire[3:0] wires_3021_6;

wire[31:0] addr_3021_6;

Selector_2 s3021_6(wires_755_5[1], addr_755_5, wires_3021_6,addr_3021_6);

wire[3:0] wires_3022_6;

wire[31:0] addr_3022_6;

Selector_2 s3022_6(wires_755_5[2], addr_755_5, wires_3022_6,addr_3022_6);

wire[3:0] wires_3023_6;

wire[31:0] addr_3023_6;

Selector_2 s3023_6(wires_755_5[3], addr_755_5, wires_3023_6,addr_3023_6);

wire[3:0] wires_3024_6;

wire[31:0] addr_3024_6;

Selector_2 s3024_6(wires_756_5[0], addr_756_5, wires_3024_6,addr_3024_6);

wire[3:0] wires_3025_6;

wire[31:0] addr_3025_6;

Selector_2 s3025_6(wires_756_5[1], addr_756_5, wires_3025_6,addr_3025_6);

wire[3:0] wires_3026_6;

wire[31:0] addr_3026_6;

Selector_2 s3026_6(wires_756_5[2], addr_756_5, wires_3026_6,addr_3026_6);

wire[3:0] wires_3027_6;

wire[31:0] addr_3027_6;

Selector_2 s3027_6(wires_756_5[3], addr_756_5, wires_3027_6,addr_3027_6);

wire[3:0] wires_3028_6;

wire[31:0] addr_3028_6;

Selector_2 s3028_6(wires_757_5[0], addr_757_5, wires_3028_6,addr_3028_6);

wire[3:0] wires_3029_6;

wire[31:0] addr_3029_6;

Selector_2 s3029_6(wires_757_5[1], addr_757_5, wires_3029_6,addr_3029_6);

wire[3:0] wires_3030_6;

wire[31:0] addr_3030_6;

Selector_2 s3030_6(wires_757_5[2], addr_757_5, wires_3030_6,addr_3030_6);

wire[3:0] wires_3031_6;

wire[31:0] addr_3031_6;

Selector_2 s3031_6(wires_757_5[3], addr_757_5, wires_3031_6,addr_3031_6);

wire[3:0] wires_3032_6;

wire[31:0] addr_3032_6;

Selector_2 s3032_6(wires_758_5[0], addr_758_5, wires_3032_6,addr_3032_6);

wire[3:0] wires_3033_6;

wire[31:0] addr_3033_6;

Selector_2 s3033_6(wires_758_5[1], addr_758_5, wires_3033_6,addr_3033_6);

wire[3:0] wires_3034_6;

wire[31:0] addr_3034_6;

Selector_2 s3034_6(wires_758_5[2], addr_758_5, wires_3034_6,addr_3034_6);

wire[3:0] wires_3035_6;

wire[31:0] addr_3035_6;

Selector_2 s3035_6(wires_758_5[3], addr_758_5, wires_3035_6,addr_3035_6);

wire[3:0] wires_3036_6;

wire[31:0] addr_3036_6;

Selector_2 s3036_6(wires_759_5[0], addr_759_5, wires_3036_6,addr_3036_6);

wire[3:0] wires_3037_6;

wire[31:0] addr_3037_6;

Selector_2 s3037_6(wires_759_5[1], addr_759_5, wires_3037_6,addr_3037_6);

wire[3:0] wires_3038_6;

wire[31:0] addr_3038_6;

Selector_2 s3038_6(wires_759_5[2], addr_759_5, wires_3038_6,addr_3038_6);

wire[3:0] wires_3039_6;

wire[31:0] addr_3039_6;

Selector_2 s3039_6(wires_759_5[3], addr_759_5, wires_3039_6,addr_3039_6);

wire[3:0] wires_3040_6;

wire[31:0] addr_3040_6;

Selector_2 s3040_6(wires_760_5[0], addr_760_5, wires_3040_6,addr_3040_6);

wire[3:0] wires_3041_6;

wire[31:0] addr_3041_6;

Selector_2 s3041_6(wires_760_5[1], addr_760_5, wires_3041_6,addr_3041_6);

wire[3:0] wires_3042_6;

wire[31:0] addr_3042_6;

Selector_2 s3042_6(wires_760_5[2], addr_760_5, wires_3042_6,addr_3042_6);

wire[3:0] wires_3043_6;

wire[31:0] addr_3043_6;

Selector_2 s3043_6(wires_760_5[3], addr_760_5, wires_3043_6,addr_3043_6);

wire[3:0] wires_3044_6;

wire[31:0] addr_3044_6;

Selector_2 s3044_6(wires_761_5[0], addr_761_5, wires_3044_6,addr_3044_6);

wire[3:0] wires_3045_6;

wire[31:0] addr_3045_6;

Selector_2 s3045_6(wires_761_5[1], addr_761_5, wires_3045_6,addr_3045_6);

wire[3:0] wires_3046_6;

wire[31:0] addr_3046_6;

Selector_2 s3046_6(wires_761_5[2], addr_761_5, wires_3046_6,addr_3046_6);

wire[3:0] wires_3047_6;

wire[31:0] addr_3047_6;

Selector_2 s3047_6(wires_761_5[3], addr_761_5, wires_3047_6,addr_3047_6);

wire[3:0] wires_3048_6;

wire[31:0] addr_3048_6;

Selector_2 s3048_6(wires_762_5[0], addr_762_5, wires_3048_6,addr_3048_6);

wire[3:0] wires_3049_6;

wire[31:0] addr_3049_6;

Selector_2 s3049_6(wires_762_5[1], addr_762_5, wires_3049_6,addr_3049_6);

wire[3:0] wires_3050_6;

wire[31:0] addr_3050_6;

Selector_2 s3050_6(wires_762_5[2], addr_762_5, wires_3050_6,addr_3050_6);

wire[3:0] wires_3051_6;

wire[31:0] addr_3051_6;

Selector_2 s3051_6(wires_762_5[3], addr_762_5, wires_3051_6,addr_3051_6);

wire[3:0] wires_3052_6;

wire[31:0] addr_3052_6;

Selector_2 s3052_6(wires_763_5[0], addr_763_5, wires_3052_6,addr_3052_6);

wire[3:0] wires_3053_6;

wire[31:0] addr_3053_6;

Selector_2 s3053_6(wires_763_5[1], addr_763_5, wires_3053_6,addr_3053_6);

wire[3:0] wires_3054_6;

wire[31:0] addr_3054_6;

Selector_2 s3054_6(wires_763_5[2], addr_763_5, wires_3054_6,addr_3054_6);

wire[3:0] wires_3055_6;

wire[31:0] addr_3055_6;

Selector_2 s3055_6(wires_763_5[3], addr_763_5, wires_3055_6,addr_3055_6);

wire[3:0] wires_3056_6;

wire[31:0] addr_3056_6;

Selector_2 s3056_6(wires_764_5[0], addr_764_5, wires_3056_6,addr_3056_6);

wire[3:0] wires_3057_6;

wire[31:0] addr_3057_6;

Selector_2 s3057_6(wires_764_5[1], addr_764_5, wires_3057_6,addr_3057_6);

wire[3:0] wires_3058_6;

wire[31:0] addr_3058_6;

Selector_2 s3058_6(wires_764_5[2], addr_764_5, wires_3058_6,addr_3058_6);

wire[3:0] wires_3059_6;

wire[31:0] addr_3059_6;

Selector_2 s3059_6(wires_764_5[3], addr_764_5, wires_3059_6,addr_3059_6);

wire[3:0] wires_3060_6;

wire[31:0] addr_3060_6;

Selector_2 s3060_6(wires_765_5[0], addr_765_5, wires_3060_6,addr_3060_6);

wire[3:0] wires_3061_6;

wire[31:0] addr_3061_6;

Selector_2 s3061_6(wires_765_5[1], addr_765_5, wires_3061_6,addr_3061_6);

wire[3:0] wires_3062_6;

wire[31:0] addr_3062_6;

Selector_2 s3062_6(wires_765_5[2], addr_765_5, wires_3062_6,addr_3062_6);

wire[3:0] wires_3063_6;

wire[31:0] addr_3063_6;

Selector_2 s3063_6(wires_765_5[3], addr_765_5, wires_3063_6,addr_3063_6);

wire[3:0] wires_3064_6;

wire[31:0] addr_3064_6;

Selector_2 s3064_6(wires_766_5[0], addr_766_5, wires_3064_6,addr_3064_6);

wire[3:0] wires_3065_6;

wire[31:0] addr_3065_6;

Selector_2 s3065_6(wires_766_5[1], addr_766_5, wires_3065_6,addr_3065_6);

wire[3:0] wires_3066_6;

wire[31:0] addr_3066_6;

Selector_2 s3066_6(wires_766_5[2], addr_766_5, wires_3066_6,addr_3066_6);

wire[3:0] wires_3067_6;

wire[31:0] addr_3067_6;

Selector_2 s3067_6(wires_766_5[3], addr_766_5, wires_3067_6,addr_3067_6);

wire[3:0] wires_3068_6;

wire[31:0] addr_3068_6;

Selector_2 s3068_6(wires_767_5[0], addr_767_5, wires_3068_6,addr_3068_6);

wire[3:0] wires_3069_6;

wire[31:0] addr_3069_6;

Selector_2 s3069_6(wires_767_5[1], addr_767_5, wires_3069_6,addr_3069_6);

wire[3:0] wires_3070_6;

wire[31:0] addr_3070_6;

Selector_2 s3070_6(wires_767_5[2], addr_767_5, wires_3070_6,addr_3070_6);

wire[3:0] wires_3071_6;

wire[31:0] addr_3071_6;

Selector_2 s3071_6(wires_767_5[3], addr_767_5, wires_3071_6,addr_3071_6);

wire[3:0] wires_3072_6;

wire[31:0] addr_3072_6;

Selector_2 s3072_6(wires_768_5[0], addr_768_5, wires_3072_6,addr_3072_6);

wire[3:0] wires_3073_6;

wire[31:0] addr_3073_6;

Selector_2 s3073_6(wires_768_5[1], addr_768_5, wires_3073_6,addr_3073_6);

wire[3:0] wires_3074_6;

wire[31:0] addr_3074_6;

Selector_2 s3074_6(wires_768_5[2], addr_768_5, wires_3074_6,addr_3074_6);

wire[3:0] wires_3075_6;

wire[31:0] addr_3075_6;

Selector_2 s3075_6(wires_768_5[3], addr_768_5, wires_3075_6,addr_3075_6);

wire[3:0] wires_3076_6;

wire[31:0] addr_3076_6;

Selector_2 s3076_6(wires_769_5[0], addr_769_5, wires_3076_6,addr_3076_6);

wire[3:0] wires_3077_6;

wire[31:0] addr_3077_6;

Selector_2 s3077_6(wires_769_5[1], addr_769_5, wires_3077_6,addr_3077_6);

wire[3:0] wires_3078_6;

wire[31:0] addr_3078_6;

Selector_2 s3078_6(wires_769_5[2], addr_769_5, wires_3078_6,addr_3078_6);

wire[3:0] wires_3079_6;

wire[31:0] addr_3079_6;

Selector_2 s3079_6(wires_769_5[3], addr_769_5, wires_3079_6,addr_3079_6);

wire[3:0] wires_3080_6;

wire[31:0] addr_3080_6;

Selector_2 s3080_6(wires_770_5[0], addr_770_5, wires_3080_6,addr_3080_6);

wire[3:0] wires_3081_6;

wire[31:0] addr_3081_6;

Selector_2 s3081_6(wires_770_5[1], addr_770_5, wires_3081_6,addr_3081_6);

wire[3:0] wires_3082_6;

wire[31:0] addr_3082_6;

Selector_2 s3082_6(wires_770_5[2], addr_770_5, wires_3082_6,addr_3082_6);

wire[3:0] wires_3083_6;

wire[31:0] addr_3083_6;

Selector_2 s3083_6(wires_770_5[3], addr_770_5, wires_3083_6,addr_3083_6);

wire[3:0] wires_3084_6;

wire[31:0] addr_3084_6;

Selector_2 s3084_6(wires_771_5[0], addr_771_5, wires_3084_6,addr_3084_6);

wire[3:0] wires_3085_6;

wire[31:0] addr_3085_6;

Selector_2 s3085_6(wires_771_5[1], addr_771_5, wires_3085_6,addr_3085_6);

wire[3:0] wires_3086_6;

wire[31:0] addr_3086_6;

Selector_2 s3086_6(wires_771_5[2], addr_771_5, wires_3086_6,addr_3086_6);

wire[3:0] wires_3087_6;

wire[31:0] addr_3087_6;

Selector_2 s3087_6(wires_771_5[3], addr_771_5, wires_3087_6,addr_3087_6);

wire[3:0] wires_3088_6;

wire[31:0] addr_3088_6;

Selector_2 s3088_6(wires_772_5[0], addr_772_5, wires_3088_6,addr_3088_6);

wire[3:0] wires_3089_6;

wire[31:0] addr_3089_6;

Selector_2 s3089_6(wires_772_5[1], addr_772_5, wires_3089_6,addr_3089_6);

wire[3:0] wires_3090_6;

wire[31:0] addr_3090_6;

Selector_2 s3090_6(wires_772_5[2], addr_772_5, wires_3090_6,addr_3090_6);

wire[3:0] wires_3091_6;

wire[31:0] addr_3091_6;

Selector_2 s3091_6(wires_772_5[3], addr_772_5, wires_3091_6,addr_3091_6);

wire[3:0] wires_3092_6;

wire[31:0] addr_3092_6;

Selector_2 s3092_6(wires_773_5[0], addr_773_5, wires_3092_6,addr_3092_6);

wire[3:0] wires_3093_6;

wire[31:0] addr_3093_6;

Selector_2 s3093_6(wires_773_5[1], addr_773_5, wires_3093_6,addr_3093_6);

wire[3:0] wires_3094_6;

wire[31:0] addr_3094_6;

Selector_2 s3094_6(wires_773_5[2], addr_773_5, wires_3094_6,addr_3094_6);

wire[3:0] wires_3095_6;

wire[31:0] addr_3095_6;

Selector_2 s3095_6(wires_773_5[3], addr_773_5, wires_3095_6,addr_3095_6);

wire[3:0] wires_3096_6;

wire[31:0] addr_3096_6;

Selector_2 s3096_6(wires_774_5[0], addr_774_5, wires_3096_6,addr_3096_6);

wire[3:0] wires_3097_6;

wire[31:0] addr_3097_6;

Selector_2 s3097_6(wires_774_5[1], addr_774_5, wires_3097_6,addr_3097_6);

wire[3:0] wires_3098_6;

wire[31:0] addr_3098_6;

Selector_2 s3098_6(wires_774_5[2], addr_774_5, wires_3098_6,addr_3098_6);

wire[3:0] wires_3099_6;

wire[31:0] addr_3099_6;

Selector_2 s3099_6(wires_774_5[3], addr_774_5, wires_3099_6,addr_3099_6);

wire[3:0] wires_3100_6;

wire[31:0] addr_3100_6;

Selector_2 s3100_6(wires_775_5[0], addr_775_5, wires_3100_6,addr_3100_6);

wire[3:0] wires_3101_6;

wire[31:0] addr_3101_6;

Selector_2 s3101_6(wires_775_5[1], addr_775_5, wires_3101_6,addr_3101_6);

wire[3:0] wires_3102_6;

wire[31:0] addr_3102_6;

Selector_2 s3102_6(wires_775_5[2], addr_775_5, wires_3102_6,addr_3102_6);

wire[3:0] wires_3103_6;

wire[31:0] addr_3103_6;

Selector_2 s3103_6(wires_775_5[3], addr_775_5, wires_3103_6,addr_3103_6);

wire[3:0] wires_3104_6;

wire[31:0] addr_3104_6;

Selector_2 s3104_6(wires_776_5[0], addr_776_5, wires_3104_6,addr_3104_6);

wire[3:0] wires_3105_6;

wire[31:0] addr_3105_6;

Selector_2 s3105_6(wires_776_5[1], addr_776_5, wires_3105_6,addr_3105_6);

wire[3:0] wires_3106_6;

wire[31:0] addr_3106_6;

Selector_2 s3106_6(wires_776_5[2], addr_776_5, wires_3106_6,addr_3106_6);

wire[3:0] wires_3107_6;

wire[31:0] addr_3107_6;

Selector_2 s3107_6(wires_776_5[3], addr_776_5, wires_3107_6,addr_3107_6);

wire[3:0] wires_3108_6;

wire[31:0] addr_3108_6;

Selector_2 s3108_6(wires_777_5[0], addr_777_5, wires_3108_6,addr_3108_6);

wire[3:0] wires_3109_6;

wire[31:0] addr_3109_6;

Selector_2 s3109_6(wires_777_5[1], addr_777_5, wires_3109_6,addr_3109_6);

wire[3:0] wires_3110_6;

wire[31:0] addr_3110_6;

Selector_2 s3110_6(wires_777_5[2], addr_777_5, wires_3110_6,addr_3110_6);

wire[3:0] wires_3111_6;

wire[31:0] addr_3111_6;

Selector_2 s3111_6(wires_777_5[3], addr_777_5, wires_3111_6,addr_3111_6);

wire[3:0] wires_3112_6;

wire[31:0] addr_3112_6;

Selector_2 s3112_6(wires_778_5[0], addr_778_5, wires_3112_6,addr_3112_6);

wire[3:0] wires_3113_6;

wire[31:0] addr_3113_6;

Selector_2 s3113_6(wires_778_5[1], addr_778_5, wires_3113_6,addr_3113_6);

wire[3:0] wires_3114_6;

wire[31:0] addr_3114_6;

Selector_2 s3114_6(wires_778_5[2], addr_778_5, wires_3114_6,addr_3114_6);

wire[3:0] wires_3115_6;

wire[31:0] addr_3115_6;

Selector_2 s3115_6(wires_778_5[3], addr_778_5, wires_3115_6,addr_3115_6);

wire[3:0] wires_3116_6;

wire[31:0] addr_3116_6;

Selector_2 s3116_6(wires_779_5[0], addr_779_5, wires_3116_6,addr_3116_6);

wire[3:0] wires_3117_6;

wire[31:0] addr_3117_6;

Selector_2 s3117_6(wires_779_5[1], addr_779_5, wires_3117_6,addr_3117_6);

wire[3:0] wires_3118_6;

wire[31:0] addr_3118_6;

Selector_2 s3118_6(wires_779_5[2], addr_779_5, wires_3118_6,addr_3118_6);

wire[3:0] wires_3119_6;

wire[31:0] addr_3119_6;

Selector_2 s3119_6(wires_779_5[3], addr_779_5, wires_3119_6,addr_3119_6);

wire[3:0] wires_3120_6;

wire[31:0] addr_3120_6;

Selector_2 s3120_6(wires_780_5[0], addr_780_5, wires_3120_6,addr_3120_6);

wire[3:0] wires_3121_6;

wire[31:0] addr_3121_6;

Selector_2 s3121_6(wires_780_5[1], addr_780_5, wires_3121_6,addr_3121_6);

wire[3:0] wires_3122_6;

wire[31:0] addr_3122_6;

Selector_2 s3122_6(wires_780_5[2], addr_780_5, wires_3122_6,addr_3122_6);

wire[3:0] wires_3123_6;

wire[31:0] addr_3123_6;

Selector_2 s3123_6(wires_780_5[3], addr_780_5, wires_3123_6,addr_3123_6);

wire[3:0] wires_3124_6;

wire[31:0] addr_3124_6;

Selector_2 s3124_6(wires_781_5[0], addr_781_5, wires_3124_6,addr_3124_6);

wire[3:0] wires_3125_6;

wire[31:0] addr_3125_6;

Selector_2 s3125_6(wires_781_5[1], addr_781_5, wires_3125_6,addr_3125_6);

wire[3:0] wires_3126_6;

wire[31:0] addr_3126_6;

Selector_2 s3126_6(wires_781_5[2], addr_781_5, wires_3126_6,addr_3126_6);

wire[3:0] wires_3127_6;

wire[31:0] addr_3127_6;

Selector_2 s3127_6(wires_781_5[3], addr_781_5, wires_3127_6,addr_3127_6);

wire[3:0] wires_3128_6;

wire[31:0] addr_3128_6;

Selector_2 s3128_6(wires_782_5[0], addr_782_5, wires_3128_6,addr_3128_6);

wire[3:0] wires_3129_6;

wire[31:0] addr_3129_6;

Selector_2 s3129_6(wires_782_5[1], addr_782_5, wires_3129_6,addr_3129_6);

wire[3:0] wires_3130_6;

wire[31:0] addr_3130_6;

Selector_2 s3130_6(wires_782_5[2], addr_782_5, wires_3130_6,addr_3130_6);

wire[3:0] wires_3131_6;

wire[31:0] addr_3131_6;

Selector_2 s3131_6(wires_782_5[3], addr_782_5, wires_3131_6,addr_3131_6);

wire[3:0] wires_3132_6;

wire[31:0] addr_3132_6;

Selector_2 s3132_6(wires_783_5[0], addr_783_5, wires_3132_6,addr_3132_6);

wire[3:0] wires_3133_6;

wire[31:0] addr_3133_6;

Selector_2 s3133_6(wires_783_5[1], addr_783_5, wires_3133_6,addr_3133_6);

wire[3:0] wires_3134_6;

wire[31:0] addr_3134_6;

Selector_2 s3134_6(wires_783_5[2], addr_783_5, wires_3134_6,addr_3134_6);

wire[3:0] wires_3135_6;

wire[31:0] addr_3135_6;

Selector_2 s3135_6(wires_783_5[3], addr_783_5, wires_3135_6,addr_3135_6);

wire[3:0] wires_3136_6;

wire[31:0] addr_3136_6;

Selector_2 s3136_6(wires_784_5[0], addr_784_5, wires_3136_6,addr_3136_6);

wire[3:0] wires_3137_6;

wire[31:0] addr_3137_6;

Selector_2 s3137_6(wires_784_5[1], addr_784_5, wires_3137_6,addr_3137_6);

wire[3:0] wires_3138_6;

wire[31:0] addr_3138_6;

Selector_2 s3138_6(wires_784_5[2], addr_784_5, wires_3138_6,addr_3138_6);

wire[3:0] wires_3139_6;

wire[31:0] addr_3139_6;

Selector_2 s3139_6(wires_784_5[3], addr_784_5, wires_3139_6,addr_3139_6);

wire[3:0] wires_3140_6;

wire[31:0] addr_3140_6;

Selector_2 s3140_6(wires_785_5[0], addr_785_5, wires_3140_6,addr_3140_6);

wire[3:0] wires_3141_6;

wire[31:0] addr_3141_6;

Selector_2 s3141_6(wires_785_5[1], addr_785_5, wires_3141_6,addr_3141_6);

wire[3:0] wires_3142_6;

wire[31:0] addr_3142_6;

Selector_2 s3142_6(wires_785_5[2], addr_785_5, wires_3142_6,addr_3142_6);

wire[3:0] wires_3143_6;

wire[31:0] addr_3143_6;

Selector_2 s3143_6(wires_785_5[3], addr_785_5, wires_3143_6,addr_3143_6);

wire[3:0] wires_3144_6;

wire[31:0] addr_3144_6;

Selector_2 s3144_6(wires_786_5[0], addr_786_5, wires_3144_6,addr_3144_6);

wire[3:0] wires_3145_6;

wire[31:0] addr_3145_6;

Selector_2 s3145_6(wires_786_5[1], addr_786_5, wires_3145_6,addr_3145_6);

wire[3:0] wires_3146_6;

wire[31:0] addr_3146_6;

Selector_2 s3146_6(wires_786_5[2], addr_786_5, wires_3146_6,addr_3146_6);

wire[3:0] wires_3147_6;

wire[31:0] addr_3147_6;

Selector_2 s3147_6(wires_786_5[3], addr_786_5, wires_3147_6,addr_3147_6);

wire[3:0] wires_3148_6;

wire[31:0] addr_3148_6;

Selector_2 s3148_6(wires_787_5[0], addr_787_5, wires_3148_6,addr_3148_6);

wire[3:0] wires_3149_6;

wire[31:0] addr_3149_6;

Selector_2 s3149_6(wires_787_5[1], addr_787_5, wires_3149_6,addr_3149_6);

wire[3:0] wires_3150_6;

wire[31:0] addr_3150_6;

Selector_2 s3150_6(wires_787_5[2], addr_787_5, wires_3150_6,addr_3150_6);

wire[3:0] wires_3151_6;

wire[31:0] addr_3151_6;

Selector_2 s3151_6(wires_787_5[3], addr_787_5, wires_3151_6,addr_3151_6);

wire[3:0] wires_3152_6;

wire[31:0] addr_3152_6;

Selector_2 s3152_6(wires_788_5[0], addr_788_5, wires_3152_6,addr_3152_6);

wire[3:0] wires_3153_6;

wire[31:0] addr_3153_6;

Selector_2 s3153_6(wires_788_5[1], addr_788_5, wires_3153_6,addr_3153_6);

wire[3:0] wires_3154_6;

wire[31:0] addr_3154_6;

Selector_2 s3154_6(wires_788_5[2], addr_788_5, wires_3154_6,addr_3154_6);

wire[3:0] wires_3155_6;

wire[31:0] addr_3155_6;

Selector_2 s3155_6(wires_788_5[3], addr_788_5, wires_3155_6,addr_3155_6);

wire[3:0] wires_3156_6;

wire[31:0] addr_3156_6;

Selector_2 s3156_6(wires_789_5[0], addr_789_5, wires_3156_6,addr_3156_6);

wire[3:0] wires_3157_6;

wire[31:0] addr_3157_6;

Selector_2 s3157_6(wires_789_5[1], addr_789_5, wires_3157_6,addr_3157_6);

wire[3:0] wires_3158_6;

wire[31:0] addr_3158_6;

Selector_2 s3158_6(wires_789_5[2], addr_789_5, wires_3158_6,addr_3158_6);

wire[3:0] wires_3159_6;

wire[31:0] addr_3159_6;

Selector_2 s3159_6(wires_789_5[3], addr_789_5, wires_3159_6,addr_3159_6);

wire[3:0] wires_3160_6;

wire[31:0] addr_3160_6;

Selector_2 s3160_6(wires_790_5[0], addr_790_5, wires_3160_6,addr_3160_6);

wire[3:0] wires_3161_6;

wire[31:0] addr_3161_6;

Selector_2 s3161_6(wires_790_5[1], addr_790_5, wires_3161_6,addr_3161_6);

wire[3:0] wires_3162_6;

wire[31:0] addr_3162_6;

Selector_2 s3162_6(wires_790_5[2], addr_790_5, wires_3162_6,addr_3162_6);

wire[3:0] wires_3163_6;

wire[31:0] addr_3163_6;

Selector_2 s3163_6(wires_790_5[3], addr_790_5, wires_3163_6,addr_3163_6);

wire[3:0] wires_3164_6;

wire[31:0] addr_3164_6;

Selector_2 s3164_6(wires_791_5[0], addr_791_5, wires_3164_6,addr_3164_6);

wire[3:0] wires_3165_6;

wire[31:0] addr_3165_6;

Selector_2 s3165_6(wires_791_5[1], addr_791_5, wires_3165_6,addr_3165_6);

wire[3:0] wires_3166_6;

wire[31:0] addr_3166_6;

Selector_2 s3166_6(wires_791_5[2], addr_791_5, wires_3166_6,addr_3166_6);

wire[3:0] wires_3167_6;

wire[31:0] addr_3167_6;

Selector_2 s3167_6(wires_791_5[3], addr_791_5, wires_3167_6,addr_3167_6);

wire[3:0] wires_3168_6;

wire[31:0] addr_3168_6;

Selector_2 s3168_6(wires_792_5[0], addr_792_5, wires_3168_6,addr_3168_6);

wire[3:0] wires_3169_6;

wire[31:0] addr_3169_6;

Selector_2 s3169_6(wires_792_5[1], addr_792_5, wires_3169_6,addr_3169_6);

wire[3:0] wires_3170_6;

wire[31:0] addr_3170_6;

Selector_2 s3170_6(wires_792_5[2], addr_792_5, wires_3170_6,addr_3170_6);

wire[3:0] wires_3171_6;

wire[31:0] addr_3171_6;

Selector_2 s3171_6(wires_792_5[3], addr_792_5, wires_3171_6,addr_3171_6);

wire[3:0] wires_3172_6;

wire[31:0] addr_3172_6;

Selector_2 s3172_6(wires_793_5[0], addr_793_5, wires_3172_6,addr_3172_6);

wire[3:0] wires_3173_6;

wire[31:0] addr_3173_6;

Selector_2 s3173_6(wires_793_5[1], addr_793_5, wires_3173_6,addr_3173_6);

wire[3:0] wires_3174_6;

wire[31:0] addr_3174_6;

Selector_2 s3174_6(wires_793_5[2], addr_793_5, wires_3174_6,addr_3174_6);

wire[3:0] wires_3175_6;

wire[31:0] addr_3175_6;

Selector_2 s3175_6(wires_793_5[3], addr_793_5, wires_3175_6,addr_3175_6);

wire[3:0] wires_3176_6;

wire[31:0] addr_3176_6;

Selector_2 s3176_6(wires_794_5[0], addr_794_5, wires_3176_6,addr_3176_6);

wire[3:0] wires_3177_6;

wire[31:0] addr_3177_6;

Selector_2 s3177_6(wires_794_5[1], addr_794_5, wires_3177_6,addr_3177_6);

wire[3:0] wires_3178_6;

wire[31:0] addr_3178_6;

Selector_2 s3178_6(wires_794_5[2], addr_794_5, wires_3178_6,addr_3178_6);

wire[3:0] wires_3179_6;

wire[31:0] addr_3179_6;

Selector_2 s3179_6(wires_794_5[3], addr_794_5, wires_3179_6,addr_3179_6);

wire[3:0] wires_3180_6;

wire[31:0] addr_3180_6;

Selector_2 s3180_6(wires_795_5[0], addr_795_5, wires_3180_6,addr_3180_6);

wire[3:0] wires_3181_6;

wire[31:0] addr_3181_6;

Selector_2 s3181_6(wires_795_5[1], addr_795_5, wires_3181_6,addr_3181_6);

wire[3:0] wires_3182_6;

wire[31:0] addr_3182_6;

Selector_2 s3182_6(wires_795_5[2], addr_795_5, wires_3182_6,addr_3182_6);

wire[3:0] wires_3183_6;

wire[31:0] addr_3183_6;

Selector_2 s3183_6(wires_795_5[3], addr_795_5, wires_3183_6,addr_3183_6);

wire[3:0] wires_3184_6;

wire[31:0] addr_3184_6;

Selector_2 s3184_6(wires_796_5[0], addr_796_5, wires_3184_6,addr_3184_6);

wire[3:0] wires_3185_6;

wire[31:0] addr_3185_6;

Selector_2 s3185_6(wires_796_5[1], addr_796_5, wires_3185_6,addr_3185_6);

wire[3:0] wires_3186_6;

wire[31:0] addr_3186_6;

Selector_2 s3186_6(wires_796_5[2], addr_796_5, wires_3186_6,addr_3186_6);

wire[3:0] wires_3187_6;

wire[31:0] addr_3187_6;

Selector_2 s3187_6(wires_796_5[3], addr_796_5, wires_3187_6,addr_3187_6);

wire[3:0] wires_3188_6;

wire[31:0] addr_3188_6;

Selector_2 s3188_6(wires_797_5[0], addr_797_5, wires_3188_6,addr_3188_6);

wire[3:0] wires_3189_6;

wire[31:0] addr_3189_6;

Selector_2 s3189_6(wires_797_5[1], addr_797_5, wires_3189_6,addr_3189_6);

wire[3:0] wires_3190_6;

wire[31:0] addr_3190_6;

Selector_2 s3190_6(wires_797_5[2], addr_797_5, wires_3190_6,addr_3190_6);

wire[3:0] wires_3191_6;

wire[31:0] addr_3191_6;

Selector_2 s3191_6(wires_797_5[3], addr_797_5, wires_3191_6,addr_3191_6);

wire[3:0] wires_3192_6;

wire[31:0] addr_3192_6;

Selector_2 s3192_6(wires_798_5[0], addr_798_5, wires_3192_6,addr_3192_6);

wire[3:0] wires_3193_6;

wire[31:0] addr_3193_6;

Selector_2 s3193_6(wires_798_5[1], addr_798_5, wires_3193_6,addr_3193_6);

wire[3:0] wires_3194_6;

wire[31:0] addr_3194_6;

Selector_2 s3194_6(wires_798_5[2], addr_798_5, wires_3194_6,addr_3194_6);

wire[3:0] wires_3195_6;

wire[31:0] addr_3195_6;

Selector_2 s3195_6(wires_798_5[3], addr_798_5, wires_3195_6,addr_3195_6);

wire[3:0] wires_3196_6;

wire[31:0] addr_3196_6;

Selector_2 s3196_6(wires_799_5[0], addr_799_5, wires_3196_6,addr_3196_6);

wire[3:0] wires_3197_6;

wire[31:0] addr_3197_6;

Selector_2 s3197_6(wires_799_5[1], addr_799_5, wires_3197_6,addr_3197_6);

wire[3:0] wires_3198_6;

wire[31:0] addr_3198_6;

Selector_2 s3198_6(wires_799_5[2], addr_799_5, wires_3198_6,addr_3198_6);

wire[3:0] wires_3199_6;

wire[31:0] addr_3199_6;

Selector_2 s3199_6(wires_799_5[3], addr_799_5, wires_3199_6,addr_3199_6);

wire[3:0] wires_3200_6;

wire[31:0] addr_3200_6;

Selector_2 s3200_6(wires_800_5[0], addr_800_5, wires_3200_6,addr_3200_6);

wire[3:0] wires_3201_6;

wire[31:0] addr_3201_6;

Selector_2 s3201_6(wires_800_5[1], addr_800_5, wires_3201_6,addr_3201_6);

wire[3:0] wires_3202_6;

wire[31:0] addr_3202_6;

Selector_2 s3202_6(wires_800_5[2], addr_800_5, wires_3202_6,addr_3202_6);

wire[3:0] wires_3203_6;

wire[31:0] addr_3203_6;

Selector_2 s3203_6(wires_800_5[3], addr_800_5, wires_3203_6,addr_3203_6);

wire[3:0] wires_3204_6;

wire[31:0] addr_3204_6;

Selector_2 s3204_6(wires_801_5[0], addr_801_5, wires_3204_6,addr_3204_6);

wire[3:0] wires_3205_6;

wire[31:0] addr_3205_6;

Selector_2 s3205_6(wires_801_5[1], addr_801_5, wires_3205_6,addr_3205_6);

wire[3:0] wires_3206_6;

wire[31:0] addr_3206_6;

Selector_2 s3206_6(wires_801_5[2], addr_801_5, wires_3206_6,addr_3206_6);

wire[3:0] wires_3207_6;

wire[31:0] addr_3207_6;

Selector_2 s3207_6(wires_801_5[3], addr_801_5, wires_3207_6,addr_3207_6);

wire[3:0] wires_3208_6;

wire[31:0] addr_3208_6;

Selector_2 s3208_6(wires_802_5[0], addr_802_5, wires_3208_6,addr_3208_6);

wire[3:0] wires_3209_6;

wire[31:0] addr_3209_6;

Selector_2 s3209_6(wires_802_5[1], addr_802_5, wires_3209_6,addr_3209_6);

wire[3:0] wires_3210_6;

wire[31:0] addr_3210_6;

Selector_2 s3210_6(wires_802_5[2], addr_802_5, wires_3210_6,addr_3210_6);

wire[3:0] wires_3211_6;

wire[31:0] addr_3211_6;

Selector_2 s3211_6(wires_802_5[3], addr_802_5, wires_3211_6,addr_3211_6);

wire[3:0] wires_3212_6;

wire[31:0] addr_3212_6;

Selector_2 s3212_6(wires_803_5[0], addr_803_5, wires_3212_6,addr_3212_6);

wire[3:0] wires_3213_6;

wire[31:0] addr_3213_6;

Selector_2 s3213_6(wires_803_5[1], addr_803_5, wires_3213_6,addr_3213_6);

wire[3:0] wires_3214_6;

wire[31:0] addr_3214_6;

Selector_2 s3214_6(wires_803_5[2], addr_803_5, wires_3214_6,addr_3214_6);

wire[3:0] wires_3215_6;

wire[31:0] addr_3215_6;

Selector_2 s3215_6(wires_803_5[3], addr_803_5, wires_3215_6,addr_3215_6);

wire[3:0] wires_3216_6;

wire[31:0] addr_3216_6;

Selector_2 s3216_6(wires_804_5[0], addr_804_5, wires_3216_6,addr_3216_6);

wire[3:0] wires_3217_6;

wire[31:0] addr_3217_6;

Selector_2 s3217_6(wires_804_5[1], addr_804_5, wires_3217_6,addr_3217_6);

wire[3:0] wires_3218_6;

wire[31:0] addr_3218_6;

Selector_2 s3218_6(wires_804_5[2], addr_804_5, wires_3218_6,addr_3218_6);

wire[3:0] wires_3219_6;

wire[31:0] addr_3219_6;

Selector_2 s3219_6(wires_804_5[3], addr_804_5, wires_3219_6,addr_3219_6);

wire[3:0] wires_3220_6;

wire[31:0] addr_3220_6;

Selector_2 s3220_6(wires_805_5[0], addr_805_5, wires_3220_6,addr_3220_6);

wire[3:0] wires_3221_6;

wire[31:0] addr_3221_6;

Selector_2 s3221_6(wires_805_5[1], addr_805_5, wires_3221_6,addr_3221_6);

wire[3:0] wires_3222_6;

wire[31:0] addr_3222_6;

Selector_2 s3222_6(wires_805_5[2], addr_805_5, wires_3222_6,addr_3222_6);

wire[3:0] wires_3223_6;

wire[31:0] addr_3223_6;

Selector_2 s3223_6(wires_805_5[3], addr_805_5, wires_3223_6,addr_3223_6);

wire[3:0] wires_3224_6;

wire[31:0] addr_3224_6;

Selector_2 s3224_6(wires_806_5[0], addr_806_5, wires_3224_6,addr_3224_6);

wire[3:0] wires_3225_6;

wire[31:0] addr_3225_6;

Selector_2 s3225_6(wires_806_5[1], addr_806_5, wires_3225_6,addr_3225_6);

wire[3:0] wires_3226_6;

wire[31:0] addr_3226_6;

Selector_2 s3226_6(wires_806_5[2], addr_806_5, wires_3226_6,addr_3226_6);

wire[3:0] wires_3227_6;

wire[31:0] addr_3227_6;

Selector_2 s3227_6(wires_806_5[3], addr_806_5, wires_3227_6,addr_3227_6);

wire[3:0] wires_3228_6;

wire[31:0] addr_3228_6;

Selector_2 s3228_6(wires_807_5[0], addr_807_5, wires_3228_6,addr_3228_6);

wire[3:0] wires_3229_6;

wire[31:0] addr_3229_6;

Selector_2 s3229_6(wires_807_5[1], addr_807_5, wires_3229_6,addr_3229_6);

wire[3:0] wires_3230_6;

wire[31:0] addr_3230_6;

Selector_2 s3230_6(wires_807_5[2], addr_807_5, wires_3230_6,addr_3230_6);

wire[3:0] wires_3231_6;

wire[31:0] addr_3231_6;

Selector_2 s3231_6(wires_807_5[3], addr_807_5, wires_3231_6,addr_3231_6);

wire[3:0] wires_3232_6;

wire[31:0] addr_3232_6;

Selector_2 s3232_6(wires_808_5[0], addr_808_5, wires_3232_6,addr_3232_6);

wire[3:0] wires_3233_6;

wire[31:0] addr_3233_6;

Selector_2 s3233_6(wires_808_5[1], addr_808_5, wires_3233_6,addr_3233_6);

wire[3:0] wires_3234_6;

wire[31:0] addr_3234_6;

Selector_2 s3234_6(wires_808_5[2], addr_808_5, wires_3234_6,addr_3234_6);

wire[3:0] wires_3235_6;

wire[31:0] addr_3235_6;

Selector_2 s3235_6(wires_808_5[3], addr_808_5, wires_3235_6,addr_3235_6);

wire[3:0] wires_3236_6;

wire[31:0] addr_3236_6;

Selector_2 s3236_6(wires_809_5[0], addr_809_5, wires_3236_6,addr_3236_6);

wire[3:0] wires_3237_6;

wire[31:0] addr_3237_6;

Selector_2 s3237_6(wires_809_5[1], addr_809_5, wires_3237_6,addr_3237_6);

wire[3:0] wires_3238_6;

wire[31:0] addr_3238_6;

Selector_2 s3238_6(wires_809_5[2], addr_809_5, wires_3238_6,addr_3238_6);

wire[3:0] wires_3239_6;

wire[31:0] addr_3239_6;

Selector_2 s3239_6(wires_809_5[3], addr_809_5, wires_3239_6,addr_3239_6);

wire[3:0] wires_3240_6;

wire[31:0] addr_3240_6;

Selector_2 s3240_6(wires_810_5[0], addr_810_5, wires_3240_6,addr_3240_6);

wire[3:0] wires_3241_6;

wire[31:0] addr_3241_6;

Selector_2 s3241_6(wires_810_5[1], addr_810_5, wires_3241_6,addr_3241_6);

wire[3:0] wires_3242_6;

wire[31:0] addr_3242_6;

Selector_2 s3242_6(wires_810_5[2], addr_810_5, wires_3242_6,addr_3242_6);

wire[3:0] wires_3243_6;

wire[31:0] addr_3243_6;

Selector_2 s3243_6(wires_810_5[3], addr_810_5, wires_3243_6,addr_3243_6);

wire[3:0] wires_3244_6;

wire[31:0] addr_3244_6;

Selector_2 s3244_6(wires_811_5[0], addr_811_5, wires_3244_6,addr_3244_6);

wire[3:0] wires_3245_6;

wire[31:0] addr_3245_6;

Selector_2 s3245_6(wires_811_5[1], addr_811_5, wires_3245_6,addr_3245_6);

wire[3:0] wires_3246_6;

wire[31:0] addr_3246_6;

Selector_2 s3246_6(wires_811_5[2], addr_811_5, wires_3246_6,addr_3246_6);

wire[3:0] wires_3247_6;

wire[31:0] addr_3247_6;

Selector_2 s3247_6(wires_811_5[3], addr_811_5, wires_3247_6,addr_3247_6);

wire[3:0] wires_3248_6;

wire[31:0] addr_3248_6;

Selector_2 s3248_6(wires_812_5[0], addr_812_5, wires_3248_6,addr_3248_6);

wire[3:0] wires_3249_6;

wire[31:0] addr_3249_6;

Selector_2 s3249_6(wires_812_5[1], addr_812_5, wires_3249_6,addr_3249_6);

wire[3:0] wires_3250_6;

wire[31:0] addr_3250_6;

Selector_2 s3250_6(wires_812_5[2], addr_812_5, wires_3250_6,addr_3250_6);

wire[3:0] wires_3251_6;

wire[31:0] addr_3251_6;

Selector_2 s3251_6(wires_812_5[3], addr_812_5, wires_3251_6,addr_3251_6);

wire[3:0] wires_3252_6;

wire[31:0] addr_3252_6;

Selector_2 s3252_6(wires_813_5[0], addr_813_5, wires_3252_6,addr_3252_6);

wire[3:0] wires_3253_6;

wire[31:0] addr_3253_6;

Selector_2 s3253_6(wires_813_5[1], addr_813_5, wires_3253_6,addr_3253_6);

wire[3:0] wires_3254_6;

wire[31:0] addr_3254_6;

Selector_2 s3254_6(wires_813_5[2], addr_813_5, wires_3254_6,addr_3254_6);

wire[3:0] wires_3255_6;

wire[31:0] addr_3255_6;

Selector_2 s3255_6(wires_813_5[3], addr_813_5, wires_3255_6,addr_3255_6);

wire[3:0] wires_3256_6;

wire[31:0] addr_3256_6;

Selector_2 s3256_6(wires_814_5[0], addr_814_5, wires_3256_6,addr_3256_6);

wire[3:0] wires_3257_6;

wire[31:0] addr_3257_6;

Selector_2 s3257_6(wires_814_5[1], addr_814_5, wires_3257_6,addr_3257_6);

wire[3:0] wires_3258_6;

wire[31:0] addr_3258_6;

Selector_2 s3258_6(wires_814_5[2], addr_814_5, wires_3258_6,addr_3258_6);

wire[3:0] wires_3259_6;

wire[31:0] addr_3259_6;

Selector_2 s3259_6(wires_814_5[3], addr_814_5, wires_3259_6,addr_3259_6);

wire[3:0] wires_3260_6;

wire[31:0] addr_3260_6;

Selector_2 s3260_6(wires_815_5[0], addr_815_5, wires_3260_6,addr_3260_6);

wire[3:0] wires_3261_6;

wire[31:0] addr_3261_6;

Selector_2 s3261_6(wires_815_5[1], addr_815_5, wires_3261_6,addr_3261_6);

wire[3:0] wires_3262_6;

wire[31:0] addr_3262_6;

Selector_2 s3262_6(wires_815_5[2], addr_815_5, wires_3262_6,addr_3262_6);

wire[3:0] wires_3263_6;

wire[31:0] addr_3263_6;

Selector_2 s3263_6(wires_815_5[3], addr_815_5, wires_3263_6,addr_3263_6);

wire[3:0] wires_3264_6;

wire[31:0] addr_3264_6;

Selector_2 s3264_6(wires_816_5[0], addr_816_5, wires_3264_6,addr_3264_6);

wire[3:0] wires_3265_6;

wire[31:0] addr_3265_6;

Selector_2 s3265_6(wires_816_5[1], addr_816_5, wires_3265_6,addr_3265_6);

wire[3:0] wires_3266_6;

wire[31:0] addr_3266_6;

Selector_2 s3266_6(wires_816_5[2], addr_816_5, wires_3266_6,addr_3266_6);

wire[3:0] wires_3267_6;

wire[31:0] addr_3267_6;

Selector_2 s3267_6(wires_816_5[3], addr_816_5, wires_3267_6,addr_3267_6);

wire[3:0] wires_3268_6;

wire[31:0] addr_3268_6;

Selector_2 s3268_6(wires_817_5[0], addr_817_5, wires_3268_6,addr_3268_6);

wire[3:0] wires_3269_6;

wire[31:0] addr_3269_6;

Selector_2 s3269_6(wires_817_5[1], addr_817_5, wires_3269_6,addr_3269_6);

wire[3:0] wires_3270_6;

wire[31:0] addr_3270_6;

Selector_2 s3270_6(wires_817_5[2], addr_817_5, wires_3270_6,addr_3270_6);

wire[3:0] wires_3271_6;

wire[31:0] addr_3271_6;

Selector_2 s3271_6(wires_817_5[3], addr_817_5, wires_3271_6,addr_3271_6);

wire[3:0] wires_3272_6;

wire[31:0] addr_3272_6;

Selector_2 s3272_6(wires_818_5[0], addr_818_5, wires_3272_6,addr_3272_6);

wire[3:0] wires_3273_6;

wire[31:0] addr_3273_6;

Selector_2 s3273_6(wires_818_5[1], addr_818_5, wires_3273_6,addr_3273_6);

wire[3:0] wires_3274_6;

wire[31:0] addr_3274_6;

Selector_2 s3274_6(wires_818_5[2], addr_818_5, wires_3274_6,addr_3274_6);

wire[3:0] wires_3275_6;

wire[31:0] addr_3275_6;

Selector_2 s3275_6(wires_818_5[3], addr_818_5, wires_3275_6,addr_3275_6);

wire[3:0] wires_3276_6;

wire[31:0] addr_3276_6;

Selector_2 s3276_6(wires_819_5[0], addr_819_5, wires_3276_6,addr_3276_6);

wire[3:0] wires_3277_6;

wire[31:0] addr_3277_6;

Selector_2 s3277_6(wires_819_5[1], addr_819_5, wires_3277_6,addr_3277_6);

wire[3:0] wires_3278_6;

wire[31:0] addr_3278_6;

Selector_2 s3278_6(wires_819_5[2], addr_819_5, wires_3278_6,addr_3278_6);

wire[3:0] wires_3279_6;

wire[31:0] addr_3279_6;

Selector_2 s3279_6(wires_819_5[3], addr_819_5, wires_3279_6,addr_3279_6);

wire[3:0] wires_3280_6;

wire[31:0] addr_3280_6;

Selector_2 s3280_6(wires_820_5[0], addr_820_5, wires_3280_6,addr_3280_6);

wire[3:0] wires_3281_6;

wire[31:0] addr_3281_6;

Selector_2 s3281_6(wires_820_5[1], addr_820_5, wires_3281_6,addr_3281_6);

wire[3:0] wires_3282_6;

wire[31:0] addr_3282_6;

Selector_2 s3282_6(wires_820_5[2], addr_820_5, wires_3282_6,addr_3282_6);

wire[3:0] wires_3283_6;

wire[31:0] addr_3283_6;

Selector_2 s3283_6(wires_820_5[3], addr_820_5, wires_3283_6,addr_3283_6);

wire[3:0] wires_3284_6;

wire[31:0] addr_3284_6;

Selector_2 s3284_6(wires_821_5[0], addr_821_5, wires_3284_6,addr_3284_6);

wire[3:0] wires_3285_6;

wire[31:0] addr_3285_6;

Selector_2 s3285_6(wires_821_5[1], addr_821_5, wires_3285_6,addr_3285_6);

wire[3:0] wires_3286_6;

wire[31:0] addr_3286_6;

Selector_2 s3286_6(wires_821_5[2], addr_821_5, wires_3286_6,addr_3286_6);

wire[3:0] wires_3287_6;

wire[31:0] addr_3287_6;

Selector_2 s3287_6(wires_821_5[3], addr_821_5, wires_3287_6,addr_3287_6);

wire[3:0] wires_3288_6;

wire[31:0] addr_3288_6;

Selector_2 s3288_6(wires_822_5[0], addr_822_5, wires_3288_6,addr_3288_6);

wire[3:0] wires_3289_6;

wire[31:0] addr_3289_6;

Selector_2 s3289_6(wires_822_5[1], addr_822_5, wires_3289_6,addr_3289_6);

wire[3:0] wires_3290_6;

wire[31:0] addr_3290_6;

Selector_2 s3290_6(wires_822_5[2], addr_822_5, wires_3290_6,addr_3290_6);

wire[3:0] wires_3291_6;

wire[31:0] addr_3291_6;

Selector_2 s3291_6(wires_822_5[3], addr_822_5, wires_3291_6,addr_3291_6);

wire[3:0] wires_3292_6;

wire[31:0] addr_3292_6;

Selector_2 s3292_6(wires_823_5[0], addr_823_5, wires_3292_6,addr_3292_6);

wire[3:0] wires_3293_6;

wire[31:0] addr_3293_6;

Selector_2 s3293_6(wires_823_5[1], addr_823_5, wires_3293_6,addr_3293_6);

wire[3:0] wires_3294_6;

wire[31:0] addr_3294_6;

Selector_2 s3294_6(wires_823_5[2], addr_823_5, wires_3294_6,addr_3294_6);

wire[3:0] wires_3295_6;

wire[31:0] addr_3295_6;

Selector_2 s3295_6(wires_823_5[3], addr_823_5, wires_3295_6,addr_3295_6);

wire[3:0] wires_3296_6;

wire[31:0] addr_3296_6;

Selector_2 s3296_6(wires_824_5[0], addr_824_5, wires_3296_6,addr_3296_6);

wire[3:0] wires_3297_6;

wire[31:0] addr_3297_6;

Selector_2 s3297_6(wires_824_5[1], addr_824_5, wires_3297_6,addr_3297_6);

wire[3:0] wires_3298_6;

wire[31:0] addr_3298_6;

Selector_2 s3298_6(wires_824_5[2], addr_824_5, wires_3298_6,addr_3298_6);

wire[3:0] wires_3299_6;

wire[31:0] addr_3299_6;

Selector_2 s3299_6(wires_824_5[3], addr_824_5, wires_3299_6,addr_3299_6);

wire[3:0] wires_3300_6;

wire[31:0] addr_3300_6;

Selector_2 s3300_6(wires_825_5[0], addr_825_5, wires_3300_6,addr_3300_6);

wire[3:0] wires_3301_6;

wire[31:0] addr_3301_6;

Selector_2 s3301_6(wires_825_5[1], addr_825_5, wires_3301_6,addr_3301_6);

wire[3:0] wires_3302_6;

wire[31:0] addr_3302_6;

Selector_2 s3302_6(wires_825_5[2], addr_825_5, wires_3302_6,addr_3302_6);

wire[3:0] wires_3303_6;

wire[31:0] addr_3303_6;

Selector_2 s3303_6(wires_825_5[3], addr_825_5, wires_3303_6,addr_3303_6);

wire[3:0] wires_3304_6;

wire[31:0] addr_3304_6;

Selector_2 s3304_6(wires_826_5[0], addr_826_5, wires_3304_6,addr_3304_6);

wire[3:0] wires_3305_6;

wire[31:0] addr_3305_6;

Selector_2 s3305_6(wires_826_5[1], addr_826_5, wires_3305_6,addr_3305_6);

wire[3:0] wires_3306_6;

wire[31:0] addr_3306_6;

Selector_2 s3306_6(wires_826_5[2], addr_826_5, wires_3306_6,addr_3306_6);

wire[3:0] wires_3307_6;

wire[31:0] addr_3307_6;

Selector_2 s3307_6(wires_826_5[3], addr_826_5, wires_3307_6,addr_3307_6);

wire[3:0] wires_3308_6;

wire[31:0] addr_3308_6;

Selector_2 s3308_6(wires_827_5[0], addr_827_5, wires_3308_6,addr_3308_6);

wire[3:0] wires_3309_6;

wire[31:0] addr_3309_6;

Selector_2 s3309_6(wires_827_5[1], addr_827_5, wires_3309_6,addr_3309_6);

wire[3:0] wires_3310_6;

wire[31:0] addr_3310_6;

Selector_2 s3310_6(wires_827_5[2], addr_827_5, wires_3310_6,addr_3310_6);

wire[3:0] wires_3311_6;

wire[31:0] addr_3311_6;

Selector_2 s3311_6(wires_827_5[3], addr_827_5, wires_3311_6,addr_3311_6);

wire[3:0] wires_3312_6;

wire[31:0] addr_3312_6;

Selector_2 s3312_6(wires_828_5[0], addr_828_5, wires_3312_6,addr_3312_6);

wire[3:0] wires_3313_6;

wire[31:0] addr_3313_6;

Selector_2 s3313_6(wires_828_5[1], addr_828_5, wires_3313_6,addr_3313_6);

wire[3:0] wires_3314_6;

wire[31:0] addr_3314_6;

Selector_2 s3314_6(wires_828_5[2], addr_828_5, wires_3314_6,addr_3314_6);

wire[3:0] wires_3315_6;

wire[31:0] addr_3315_6;

Selector_2 s3315_6(wires_828_5[3], addr_828_5, wires_3315_6,addr_3315_6);

wire[3:0] wires_3316_6;

wire[31:0] addr_3316_6;

Selector_2 s3316_6(wires_829_5[0], addr_829_5, wires_3316_6,addr_3316_6);

wire[3:0] wires_3317_6;

wire[31:0] addr_3317_6;

Selector_2 s3317_6(wires_829_5[1], addr_829_5, wires_3317_6,addr_3317_6);

wire[3:0] wires_3318_6;

wire[31:0] addr_3318_6;

Selector_2 s3318_6(wires_829_5[2], addr_829_5, wires_3318_6,addr_3318_6);

wire[3:0] wires_3319_6;

wire[31:0] addr_3319_6;

Selector_2 s3319_6(wires_829_5[3], addr_829_5, wires_3319_6,addr_3319_6);

wire[3:0] wires_3320_6;

wire[31:0] addr_3320_6;

Selector_2 s3320_6(wires_830_5[0], addr_830_5, wires_3320_6,addr_3320_6);

wire[3:0] wires_3321_6;

wire[31:0] addr_3321_6;

Selector_2 s3321_6(wires_830_5[1], addr_830_5, wires_3321_6,addr_3321_6);

wire[3:0] wires_3322_6;

wire[31:0] addr_3322_6;

Selector_2 s3322_6(wires_830_5[2], addr_830_5, wires_3322_6,addr_3322_6);

wire[3:0] wires_3323_6;

wire[31:0] addr_3323_6;

Selector_2 s3323_6(wires_830_5[3], addr_830_5, wires_3323_6,addr_3323_6);

wire[3:0] wires_3324_6;

wire[31:0] addr_3324_6;

Selector_2 s3324_6(wires_831_5[0], addr_831_5, wires_3324_6,addr_3324_6);

wire[3:0] wires_3325_6;

wire[31:0] addr_3325_6;

Selector_2 s3325_6(wires_831_5[1], addr_831_5, wires_3325_6,addr_3325_6);

wire[3:0] wires_3326_6;

wire[31:0] addr_3326_6;

Selector_2 s3326_6(wires_831_5[2], addr_831_5, wires_3326_6,addr_3326_6);

wire[3:0] wires_3327_6;

wire[31:0] addr_3327_6;

Selector_2 s3327_6(wires_831_5[3], addr_831_5, wires_3327_6,addr_3327_6);

wire[3:0] wires_3328_6;

wire[31:0] addr_3328_6;

Selector_2 s3328_6(wires_832_5[0], addr_832_5, wires_3328_6,addr_3328_6);

wire[3:0] wires_3329_6;

wire[31:0] addr_3329_6;

Selector_2 s3329_6(wires_832_5[1], addr_832_5, wires_3329_6,addr_3329_6);

wire[3:0] wires_3330_6;

wire[31:0] addr_3330_6;

Selector_2 s3330_6(wires_832_5[2], addr_832_5, wires_3330_6,addr_3330_6);

wire[3:0] wires_3331_6;

wire[31:0] addr_3331_6;

Selector_2 s3331_6(wires_832_5[3], addr_832_5, wires_3331_6,addr_3331_6);

wire[3:0] wires_3332_6;

wire[31:0] addr_3332_6;

Selector_2 s3332_6(wires_833_5[0], addr_833_5, wires_3332_6,addr_3332_6);

wire[3:0] wires_3333_6;

wire[31:0] addr_3333_6;

Selector_2 s3333_6(wires_833_5[1], addr_833_5, wires_3333_6,addr_3333_6);

wire[3:0] wires_3334_6;

wire[31:0] addr_3334_6;

Selector_2 s3334_6(wires_833_5[2], addr_833_5, wires_3334_6,addr_3334_6);

wire[3:0] wires_3335_6;

wire[31:0] addr_3335_6;

Selector_2 s3335_6(wires_833_5[3], addr_833_5, wires_3335_6,addr_3335_6);

wire[3:0] wires_3336_6;

wire[31:0] addr_3336_6;

Selector_2 s3336_6(wires_834_5[0], addr_834_5, wires_3336_6,addr_3336_6);

wire[3:0] wires_3337_6;

wire[31:0] addr_3337_6;

Selector_2 s3337_6(wires_834_5[1], addr_834_5, wires_3337_6,addr_3337_6);

wire[3:0] wires_3338_6;

wire[31:0] addr_3338_6;

Selector_2 s3338_6(wires_834_5[2], addr_834_5, wires_3338_6,addr_3338_6);

wire[3:0] wires_3339_6;

wire[31:0] addr_3339_6;

Selector_2 s3339_6(wires_834_5[3], addr_834_5, wires_3339_6,addr_3339_6);

wire[3:0] wires_3340_6;

wire[31:0] addr_3340_6;

Selector_2 s3340_6(wires_835_5[0], addr_835_5, wires_3340_6,addr_3340_6);

wire[3:0] wires_3341_6;

wire[31:0] addr_3341_6;

Selector_2 s3341_6(wires_835_5[1], addr_835_5, wires_3341_6,addr_3341_6);

wire[3:0] wires_3342_6;

wire[31:0] addr_3342_6;

Selector_2 s3342_6(wires_835_5[2], addr_835_5, wires_3342_6,addr_3342_6);

wire[3:0] wires_3343_6;

wire[31:0] addr_3343_6;

Selector_2 s3343_6(wires_835_5[3], addr_835_5, wires_3343_6,addr_3343_6);

wire[3:0] wires_3344_6;

wire[31:0] addr_3344_6;

Selector_2 s3344_6(wires_836_5[0], addr_836_5, wires_3344_6,addr_3344_6);

wire[3:0] wires_3345_6;

wire[31:0] addr_3345_6;

Selector_2 s3345_6(wires_836_5[1], addr_836_5, wires_3345_6,addr_3345_6);

wire[3:0] wires_3346_6;

wire[31:0] addr_3346_6;

Selector_2 s3346_6(wires_836_5[2], addr_836_5, wires_3346_6,addr_3346_6);

wire[3:0] wires_3347_6;

wire[31:0] addr_3347_6;

Selector_2 s3347_6(wires_836_5[3], addr_836_5, wires_3347_6,addr_3347_6);

wire[3:0] wires_3348_6;

wire[31:0] addr_3348_6;

Selector_2 s3348_6(wires_837_5[0], addr_837_5, wires_3348_6,addr_3348_6);

wire[3:0] wires_3349_6;

wire[31:0] addr_3349_6;

Selector_2 s3349_6(wires_837_5[1], addr_837_5, wires_3349_6,addr_3349_6);

wire[3:0] wires_3350_6;

wire[31:0] addr_3350_6;

Selector_2 s3350_6(wires_837_5[2], addr_837_5, wires_3350_6,addr_3350_6);

wire[3:0] wires_3351_6;

wire[31:0] addr_3351_6;

Selector_2 s3351_6(wires_837_5[3], addr_837_5, wires_3351_6,addr_3351_6);

wire[3:0] wires_3352_6;

wire[31:0] addr_3352_6;

Selector_2 s3352_6(wires_838_5[0], addr_838_5, wires_3352_6,addr_3352_6);

wire[3:0] wires_3353_6;

wire[31:0] addr_3353_6;

Selector_2 s3353_6(wires_838_5[1], addr_838_5, wires_3353_6,addr_3353_6);

wire[3:0] wires_3354_6;

wire[31:0] addr_3354_6;

Selector_2 s3354_6(wires_838_5[2], addr_838_5, wires_3354_6,addr_3354_6);

wire[3:0] wires_3355_6;

wire[31:0] addr_3355_6;

Selector_2 s3355_6(wires_838_5[3], addr_838_5, wires_3355_6,addr_3355_6);

wire[3:0] wires_3356_6;

wire[31:0] addr_3356_6;

Selector_2 s3356_6(wires_839_5[0], addr_839_5, wires_3356_6,addr_3356_6);

wire[3:0] wires_3357_6;

wire[31:0] addr_3357_6;

Selector_2 s3357_6(wires_839_5[1], addr_839_5, wires_3357_6,addr_3357_6);

wire[3:0] wires_3358_6;

wire[31:0] addr_3358_6;

Selector_2 s3358_6(wires_839_5[2], addr_839_5, wires_3358_6,addr_3358_6);

wire[3:0] wires_3359_6;

wire[31:0] addr_3359_6;

Selector_2 s3359_6(wires_839_5[3], addr_839_5, wires_3359_6,addr_3359_6);

wire[3:0] wires_3360_6;

wire[31:0] addr_3360_6;

Selector_2 s3360_6(wires_840_5[0], addr_840_5, wires_3360_6,addr_3360_6);

wire[3:0] wires_3361_6;

wire[31:0] addr_3361_6;

Selector_2 s3361_6(wires_840_5[1], addr_840_5, wires_3361_6,addr_3361_6);

wire[3:0] wires_3362_6;

wire[31:0] addr_3362_6;

Selector_2 s3362_6(wires_840_5[2], addr_840_5, wires_3362_6,addr_3362_6);

wire[3:0] wires_3363_6;

wire[31:0] addr_3363_6;

Selector_2 s3363_6(wires_840_5[3], addr_840_5, wires_3363_6,addr_3363_6);

wire[3:0] wires_3364_6;

wire[31:0] addr_3364_6;

Selector_2 s3364_6(wires_841_5[0], addr_841_5, wires_3364_6,addr_3364_6);

wire[3:0] wires_3365_6;

wire[31:0] addr_3365_6;

Selector_2 s3365_6(wires_841_5[1], addr_841_5, wires_3365_6,addr_3365_6);

wire[3:0] wires_3366_6;

wire[31:0] addr_3366_6;

Selector_2 s3366_6(wires_841_5[2], addr_841_5, wires_3366_6,addr_3366_6);

wire[3:0] wires_3367_6;

wire[31:0] addr_3367_6;

Selector_2 s3367_6(wires_841_5[3], addr_841_5, wires_3367_6,addr_3367_6);

wire[3:0] wires_3368_6;

wire[31:0] addr_3368_6;

Selector_2 s3368_6(wires_842_5[0], addr_842_5, wires_3368_6,addr_3368_6);

wire[3:0] wires_3369_6;

wire[31:0] addr_3369_6;

Selector_2 s3369_6(wires_842_5[1], addr_842_5, wires_3369_6,addr_3369_6);

wire[3:0] wires_3370_6;

wire[31:0] addr_3370_6;

Selector_2 s3370_6(wires_842_5[2], addr_842_5, wires_3370_6,addr_3370_6);

wire[3:0] wires_3371_6;

wire[31:0] addr_3371_6;

Selector_2 s3371_6(wires_842_5[3], addr_842_5, wires_3371_6,addr_3371_6);

wire[3:0] wires_3372_6;

wire[31:0] addr_3372_6;

Selector_2 s3372_6(wires_843_5[0], addr_843_5, wires_3372_6,addr_3372_6);

wire[3:0] wires_3373_6;

wire[31:0] addr_3373_6;

Selector_2 s3373_6(wires_843_5[1], addr_843_5, wires_3373_6,addr_3373_6);

wire[3:0] wires_3374_6;

wire[31:0] addr_3374_6;

Selector_2 s3374_6(wires_843_5[2], addr_843_5, wires_3374_6,addr_3374_6);

wire[3:0] wires_3375_6;

wire[31:0] addr_3375_6;

Selector_2 s3375_6(wires_843_5[3], addr_843_5, wires_3375_6,addr_3375_6);

wire[3:0] wires_3376_6;

wire[31:0] addr_3376_6;

Selector_2 s3376_6(wires_844_5[0], addr_844_5, wires_3376_6,addr_3376_6);

wire[3:0] wires_3377_6;

wire[31:0] addr_3377_6;

Selector_2 s3377_6(wires_844_5[1], addr_844_5, wires_3377_6,addr_3377_6);

wire[3:0] wires_3378_6;

wire[31:0] addr_3378_6;

Selector_2 s3378_6(wires_844_5[2], addr_844_5, wires_3378_6,addr_3378_6);

wire[3:0] wires_3379_6;

wire[31:0] addr_3379_6;

Selector_2 s3379_6(wires_844_5[3], addr_844_5, wires_3379_6,addr_3379_6);

wire[3:0] wires_3380_6;

wire[31:0] addr_3380_6;

Selector_2 s3380_6(wires_845_5[0], addr_845_5, wires_3380_6,addr_3380_6);

wire[3:0] wires_3381_6;

wire[31:0] addr_3381_6;

Selector_2 s3381_6(wires_845_5[1], addr_845_5, wires_3381_6,addr_3381_6);

wire[3:0] wires_3382_6;

wire[31:0] addr_3382_6;

Selector_2 s3382_6(wires_845_5[2], addr_845_5, wires_3382_6,addr_3382_6);

wire[3:0] wires_3383_6;

wire[31:0] addr_3383_6;

Selector_2 s3383_6(wires_845_5[3], addr_845_5, wires_3383_6,addr_3383_6);

wire[3:0] wires_3384_6;

wire[31:0] addr_3384_6;

Selector_2 s3384_6(wires_846_5[0], addr_846_5, wires_3384_6,addr_3384_6);

wire[3:0] wires_3385_6;

wire[31:0] addr_3385_6;

Selector_2 s3385_6(wires_846_5[1], addr_846_5, wires_3385_6,addr_3385_6);

wire[3:0] wires_3386_6;

wire[31:0] addr_3386_6;

Selector_2 s3386_6(wires_846_5[2], addr_846_5, wires_3386_6,addr_3386_6);

wire[3:0] wires_3387_6;

wire[31:0] addr_3387_6;

Selector_2 s3387_6(wires_846_5[3], addr_846_5, wires_3387_6,addr_3387_6);

wire[3:0] wires_3388_6;

wire[31:0] addr_3388_6;

Selector_2 s3388_6(wires_847_5[0], addr_847_5, wires_3388_6,addr_3388_6);

wire[3:0] wires_3389_6;

wire[31:0] addr_3389_6;

Selector_2 s3389_6(wires_847_5[1], addr_847_5, wires_3389_6,addr_3389_6);

wire[3:0] wires_3390_6;

wire[31:0] addr_3390_6;

Selector_2 s3390_6(wires_847_5[2], addr_847_5, wires_3390_6,addr_3390_6);

wire[3:0] wires_3391_6;

wire[31:0] addr_3391_6;

Selector_2 s3391_6(wires_847_5[3], addr_847_5, wires_3391_6,addr_3391_6);

wire[3:0] wires_3392_6;

wire[31:0] addr_3392_6;

Selector_2 s3392_6(wires_848_5[0], addr_848_5, wires_3392_6,addr_3392_6);

wire[3:0] wires_3393_6;

wire[31:0] addr_3393_6;

Selector_2 s3393_6(wires_848_5[1], addr_848_5, wires_3393_6,addr_3393_6);

wire[3:0] wires_3394_6;

wire[31:0] addr_3394_6;

Selector_2 s3394_6(wires_848_5[2], addr_848_5, wires_3394_6,addr_3394_6);

wire[3:0] wires_3395_6;

wire[31:0] addr_3395_6;

Selector_2 s3395_6(wires_848_5[3], addr_848_5, wires_3395_6,addr_3395_6);

wire[3:0] wires_3396_6;

wire[31:0] addr_3396_6;

Selector_2 s3396_6(wires_849_5[0], addr_849_5, wires_3396_6,addr_3396_6);

wire[3:0] wires_3397_6;

wire[31:0] addr_3397_6;

Selector_2 s3397_6(wires_849_5[1], addr_849_5, wires_3397_6,addr_3397_6);

wire[3:0] wires_3398_6;

wire[31:0] addr_3398_6;

Selector_2 s3398_6(wires_849_5[2], addr_849_5, wires_3398_6,addr_3398_6);

wire[3:0] wires_3399_6;

wire[31:0] addr_3399_6;

Selector_2 s3399_6(wires_849_5[3], addr_849_5, wires_3399_6,addr_3399_6);

wire[3:0] wires_3400_6;

wire[31:0] addr_3400_6;

Selector_2 s3400_6(wires_850_5[0], addr_850_5, wires_3400_6,addr_3400_6);

wire[3:0] wires_3401_6;

wire[31:0] addr_3401_6;

Selector_2 s3401_6(wires_850_5[1], addr_850_5, wires_3401_6,addr_3401_6);

wire[3:0] wires_3402_6;

wire[31:0] addr_3402_6;

Selector_2 s3402_6(wires_850_5[2], addr_850_5, wires_3402_6,addr_3402_6);

wire[3:0] wires_3403_6;

wire[31:0] addr_3403_6;

Selector_2 s3403_6(wires_850_5[3], addr_850_5, wires_3403_6,addr_3403_6);

wire[3:0] wires_3404_6;

wire[31:0] addr_3404_6;

Selector_2 s3404_6(wires_851_5[0], addr_851_5, wires_3404_6,addr_3404_6);

wire[3:0] wires_3405_6;

wire[31:0] addr_3405_6;

Selector_2 s3405_6(wires_851_5[1], addr_851_5, wires_3405_6,addr_3405_6);

wire[3:0] wires_3406_6;

wire[31:0] addr_3406_6;

Selector_2 s3406_6(wires_851_5[2], addr_851_5, wires_3406_6,addr_3406_6);

wire[3:0] wires_3407_6;

wire[31:0] addr_3407_6;

Selector_2 s3407_6(wires_851_5[3], addr_851_5, wires_3407_6,addr_3407_6);

wire[3:0] wires_3408_6;

wire[31:0] addr_3408_6;

Selector_2 s3408_6(wires_852_5[0], addr_852_5, wires_3408_6,addr_3408_6);

wire[3:0] wires_3409_6;

wire[31:0] addr_3409_6;

Selector_2 s3409_6(wires_852_5[1], addr_852_5, wires_3409_6,addr_3409_6);

wire[3:0] wires_3410_6;

wire[31:0] addr_3410_6;

Selector_2 s3410_6(wires_852_5[2], addr_852_5, wires_3410_6,addr_3410_6);

wire[3:0] wires_3411_6;

wire[31:0] addr_3411_6;

Selector_2 s3411_6(wires_852_5[3], addr_852_5, wires_3411_6,addr_3411_6);

wire[3:0] wires_3412_6;

wire[31:0] addr_3412_6;

Selector_2 s3412_6(wires_853_5[0], addr_853_5, wires_3412_6,addr_3412_6);

wire[3:0] wires_3413_6;

wire[31:0] addr_3413_6;

Selector_2 s3413_6(wires_853_5[1], addr_853_5, wires_3413_6,addr_3413_6);

wire[3:0] wires_3414_6;

wire[31:0] addr_3414_6;

Selector_2 s3414_6(wires_853_5[2], addr_853_5, wires_3414_6,addr_3414_6);

wire[3:0] wires_3415_6;

wire[31:0] addr_3415_6;

Selector_2 s3415_6(wires_853_5[3], addr_853_5, wires_3415_6,addr_3415_6);

wire[3:0] wires_3416_6;

wire[31:0] addr_3416_6;

Selector_2 s3416_6(wires_854_5[0], addr_854_5, wires_3416_6,addr_3416_6);

wire[3:0] wires_3417_6;

wire[31:0] addr_3417_6;

Selector_2 s3417_6(wires_854_5[1], addr_854_5, wires_3417_6,addr_3417_6);

wire[3:0] wires_3418_6;

wire[31:0] addr_3418_6;

Selector_2 s3418_6(wires_854_5[2], addr_854_5, wires_3418_6,addr_3418_6);

wire[3:0] wires_3419_6;

wire[31:0] addr_3419_6;

Selector_2 s3419_6(wires_854_5[3], addr_854_5, wires_3419_6,addr_3419_6);

wire[3:0] wires_3420_6;

wire[31:0] addr_3420_6;

Selector_2 s3420_6(wires_855_5[0], addr_855_5, wires_3420_6,addr_3420_6);

wire[3:0] wires_3421_6;

wire[31:0] addr_3421_6;

Selector_2 s3421_6(wires_855_5[1], addr_855_5, wires_3421_6,addr_3421_6);

wire[3:0] wires_3422_6;

wire[31:0] addr_3422_6;

Selector_2 s3422_6(wires_855_5[2], addr_855_5, wires_3422_6,addr_3422_6);

wire[3:0] wires_3423_6;

wire[31:0] addr_3423_6;

Selector_2 s3423_6(wires_855_5[3], addr_855_5, wires_3423_6,addr_3423_6);

wire[3:0] wires_3424_6;

wire[31:0] addr_3424_6;

Selector_2 s3424_6(wires_856_5[0], addr_856_5, wires_3424_6,addr_3424_6);

wire[3:0] wires_3425_6;

wire[31:0] addr_3425_6;

Selector_2 s3425_6(wires_856_5[1], addr_856_5, wires_3425_6,addr_3425_6);

wire[3:0] wires_3426_6;

wire[31:0] addr_3426_6;

Selector_2 s3426_6(wires_856_5[2], addr_856_5, wires_3426_6,addr_3426_6);

wire[3:0] wires_3427_6;

wire[31:0] addr_3427_6;

Selector_2 s3427_6(wires_856_5[3], addr_856_5, wires_3427_6,addr_3427_6);

wire[3:0] wires_3428_6;

wire[31:0] addr_3428_6;

Selector_2 s3428_6(wires_857_5[0], addr_857_5, wires_3428_6,addr_3428_6);

wire[3:0] wires_3429_6;

wire[31:0] addr_3429_6;

Selector_2 s3429_6(wires_857_5[1], addr_857_5, wires_3429_6,addr_3429_6);

wire[3:0] wires_3430_6;

wire[31:0] addr_3430_6;

Selector_2 s3430_6(wires_857_5[2], addr_857_5, wires_3430_6,addr_3430_6);

wire[3:0] wires_3431_6;

wire[31:0] addr_3431_6;

Selector_2 s3431_6(wires_857_5[3], addr_857_5, wires_3431_6,addr_3431_6);

wire[3:0] wires_3432_6;

wire[31:0] addr_3432_6;

Selector_2 s3432_6(wires_858_5[0], addr_858_5, wires_3432_6,addr_3432_6);

wire[3:0] wires_3433_6;

wire[31:0] addr_3433_6;

Selector_2 s3433_6(wires_858_5[1], addr_858_5, wires_3433_6,addr_3433_6);

wire[3:0] wires_3434_6;

wire[31:0] addr_3434_6;

Selector_2 s3434_6(wires_858_5[2], addr_858_5, wires_3434_6,addr_3434_6);

wire[3:0] wires_3435_6;

wire[31:0] addr_3435_6;

Selector_2 s3435_6(wires_858_5[3], addr_858_5, wires_3435_6,addr_3435_6);

wire[3:0] wires_3436_6;

wire[31:0] addr_3436_6;

Selector_2 s3436_6(wires_859_5[0], addr_859_5, wires_3436_6,addr_3436_6);

wire[3:0] wires_3437_6;

wire[31:0] addr_3437_6;

Selector_2 s3437_6(wires_859_5[1], addr_859_5, wires_3437_6,addr_3437_6);

wire[3:0] wires_3438_6;

wire[31:0] addr_3438_6;

Selector_2 s3438_6(wires_859_5[2], addr_859_5, wires_3438_6,addr_3438_6);

wire[3:0] wires_3439_6;

wire[31:0] addr_3439_6;

Selector_2 s3439_6(wires_859_5[3], addr_859_5, wires_3439_6,addr_3439_6);

wire[3:0] wires_3440_6;

wire[31:0] addr_3440_6;

Selector_2 s3440_6(wires_860_5[0], addr_860_5, wires_3440_6,addr_3440_6);

wire[3:0] wires_3441_6;

wire[31:0] addr_3441_6;

Selector_2 s3441_6(wires_860_5[1], addr_860_5, wires_3441_6,addr_3441_6);

wire[3:0] wires_3442_6;

wire[31:0] addr_3442_6;

Selector_2 s3442_6(wires_860_5[2], addr_860_5, wires_3442_6,addr_3442_6);

wire[3:0] wires_3443_6;

wire[31:0] addr_3443_6;

Selector_2 s3443_6(wires_860_5[3], addr_860_5, wires_3443_6,addr_3443_6);

wire[3:0] wires_3444_6;

wire[31:0] addr_3444_6;

Selector_2 s3444_6(wires_861_5[0], addr_861_5, wires_3444_6,addr_3444_6);

wire[3:0] wires_3445_6;

wire[31:0] addr_3445_6;

Selector_2 s3445_6(wires_861_5[1], addr_861_5, wires_3445_6,addr_3445_6);

wire[3:0] wires_3446_6;

wire[31:0] addr_3446_6;

Selector_2 s3446_6(wires_861_5[2], addr_861_5, wires_3446_6,addr_3446_6);

wire[3:0] wires_3447_6;

wire[31:0] addr_3447_6;

Selector_2 s3447_6(wires_861_5[3], addr_861_5, wires_3447_6,addr_3447_6);

wire[3:0] wires_3448_6;

wire[31:0] addr_3448_6;

Selector_2 s3448_6(wires_862_5[0], addr_862_5, wires_3448_6,addr_3448_6);

wire[3:0] wires_3449_6;

wire[31:0] addr_3449_6;

Selector_2 s3449_6(wires_862_5[1], addr_862_5, wires_3449_6,addr_3449_6);

wire[3:0] wires_3450_6;

wire[31:0] addr_3450_6;

Selector_2 s3450_6(wires_862_5[2], addr_862_5, wires_3450_6,addr_3450_6);

wire[3:0] wires_3451_6;

wire[31:0] addr_3451_6;

Selector_2 s3451_6(wires_862_5[3], addr_862_5, wires_3451_6,addr_3451_6);

wire[3:0] wires_3452_6;

wire[31:0] addr_3452_6;

Selector_2 s3452_6(wires_863_5[0], addr_863_5, wires_3452_6,addr_3452_6);

wire[3:0] wires_3453_6;

wire[31:0] addr_3453_6;

Selector_2 s3453_6(wires_863_5[1], addr_863_5, wires_3453_6,addr_3453_6);

wire[3:0] wires_3454_6;

wire[31:0] addr_3454_6;

Selector_2 s3454_6(wires_863_5[2], addr_863_5, wires_3454_6,addr_3454_6);

wire[3:0] wires_3455_6;

wire[31:0] addr_3455_6;

Selector_2 s3455_6(wires_863_5[3], addr_863_5, wires_3455_6,addr_3455_6);

wire[3:0] wires_3456_6;

wire[31:0] addr_3456_6;

Selector_2 s3456_6(wires_864_5[0], addr_864_5, wires_3456_6,addr_3456_6);

wire[3:0] wires_3457_6;

wire[31:0] addr_3457_6;

Selector_2 s3457_6(wires_864_5[1], addr_864_5, wires_3457_6,addr_3457_6);

wire[3:0] wires_3458_6;

wire[31:0] addr_3458_6;

Selector_2 s3458_6(wires_864_5[2], addr_864_5, wires_3458_6,addr_3458_6);

wire[3:0] wires_3459_6;

wire[31:0] addr_3459_6;

Selector_2 s3459_6(wires_864_5[3], addr_864_5, wires_3459_6,addr_3459_6);

wire[3:0] wires_3460_6;

wire[31:0] addr_3460_6;

Selector_2 s3460_6(wires_865_5[0], addr_865_5, wires_3460_6,addr_3460_6);

wire[3:0] wires_3461_6;

wire[31:0] addr_3461_6;

Selector_2 s3461_6(wires_865_5[1], addr_865_5, wires_3461_6,addr_3461_6);

wire[3:0] wires_3462_6;

wire[31:0] addr_3462_6;

Selector_2 s3462_6(wires_865_5[2], addr_865_5, wires_3462_6,addr_3462_6);

wire[3:0] wires_3463_6;

wire[31:0] addr_3463_6;

Selector_2 s3463_6(wires_865_5[3], addr_865_5, wires_3463_6,addr_3463_6);

wire[3:0] wires_3464_6;

wire[31:0] addr_3464_6;

Selector_2 s3464_6(wires_866_5[0], addr_866_5, wires_3464_6,addr_3464_6);

wire[3:0] wires_3465_6;

wire[31:0] addr_3465_6;

Selector_2 s3465_6(wires_866_5[1], addr_866_5, wires_3465_6,addr_3465_6);

wire[3:0] wires_3466_6;

wire[31:0] addr_3466_6;

Selector_2 s3466_6(wires_866_5[2], addr_866_5, wires_3466_6,addr_3466_6);

wire[3:0] wires_3467_6;

wire[31:0] addr_3467_6;

Selector_2 s3467_6(wires_866_5[3], addr_866_5, wires_3467_6,addr_3467_6);

wire[3:0] wires_3468_6;

wire[31:0] addr_3468_6;

Selector_2 s3468_6(wires_867_5[0], addr_867_5, wires_3468_6,addr_3468_6);

wire[3:0] wires_3469_6;

wire[31:0] addr_3469_6;

Selector_2 s3469_6(wires_867_5[1], addr_867_5, wires_3469_6,addr_3469_6);

wire[3:0] wires_3470_6;

wire[31:0] addr_3470_6;

Selector_2 s3470_6(wires_867_5[2], addr_867_5, wires_3470_6,addr_3470_6);

wire[3:0] wires_3471_6;

wire[31:0] addr_3471_6;

Selector_2 s3471_6(wires_867_5[3], addr_867_5, wires_3471_6,addr_3471_6);

wire[3:0] wires_3472_6;

wire[31:0] addr_3472_6;

Selector_2 s3472_6(wires_868_5[0], addr_868_5, wires_3472_6,addr_3472_6);

wire[3:0] wires_3473_6;

wire[31:0] addr_3473_6;

Selector_2 s3473_6(wires_868_5[1], addr_868_5, wires_3473_6,addr_3473_6);

wire[3:0] wires_3474_6;

wire[31:0] addr_3474_6;

Selector_2 s3474_6(wires_868_5[2], addr_868_5, wires_3474_6,addr_3474_6);

wire[3:0] wires_3475_6;

wire[31:0] addr_3475_6;

Selector_2 s3475_6(wires_868_5[3], addr_868_5, wires_3475_6,addr_3475_6);

wire[3:0] wires_3476_6;

wire[31:0] addr_3476_6;

Selector_2 s3476_6(wires_869_5[0], addr_869_5, wires_3476_6,addr_3476_6);

wire[3:0] wires_3477_6;

wire[31:0] addr_3477_6;

Selector_2 s3477_6(wires_869_5[1], addr_869_5, wires_3477_6,addr_3477_6);

wire[3:0] wires_3478_6;

wire[31:0] addr_3478_6;

Selector_2 s3478_6(wires_869_5[2], addr_869_5, wires_3478_6,addr_3478_6);

wire[3:0] wires_3479_6;

wire[31:0] addr_3479_6;

Selector_2 s3479_6(wires_869_5[3], addr_869_5, wires_3479_6,addr_3479_6);

wire[3:0] wires_3480_6;

wire[31:0] addr_3480_6;

Selector_2 s3480_6(wires_870_5[0], addr_870_5, wires_3480_6,addr_3480_6);

wire[3:0] wires_3481_6;

wire[31:0] addr_3481_6;

Selector_2 s3481_6(wires_870_5[1], addr_870_5, wires_3481_6,addr_3481_6);

wire[3:0] wires_3482_6;

wire[31:0] addr_3482_6;

Selector_2 s3482_6(wires_870_5[2], addr_870_5, wires_3482_6,addr_3482_6);

wire[3:0] wires_3483_6;

wire[31:0] addr_3483_6;

Selector_2 s3483_6(wires_870_5[3], addr_870_5, wires_3483_6,addr_3483_6);

wire[3:0] wires_3484_6;

wire[31:0] addr_3484_6;

Selector_2 s3484_6(wires_871_5[0], addr_871_5, wires_3484_6,addr_3484_6);

wire[3:0] wires_3485_6;

wire[31:0] addr_3485_6;

Selector_2 s3485_6(wires_871_5[1], addr_871_5, wires_3485_6,addr_3485_6);

wire[3:0] wires_3486_6;

wire[31:0] addr_3486_6;

Selector_2 s3486_6(wires_871_5[2], addr_871_5, wires_3486_6,addr_3486_6);

wire[3:0] wires_3487_6;

wire[31:0] addr_3487_6;

Selector_2 s3487_6(wires_871_5[3], addr_871_5, wires_3487_6,addr_3487_6);

wire[3:0] wires_3488_6;

wire[31:0] addr_3488_6;

Selector_2 s3488_6(wires_872_5[0], addr_872_5, wires_3488_6,addr_3488_6);

wire[3:0] wires_3489_6;

wire[31:0] addr_3489_6;

Selector_2 s3489_6(wires_872_5[1], addr_872_5, wires_3489_6,addr_3489_6);

wire[3:0] wires_3490_6;

wire[31:0] addr_3490_6;

Selector_2 s3490_6(wires_872_5[2], addr_872_5, wires_3490_6,addr_3490_6);

wire[3:0] wires_3491_6;

wire[31:0] addr_3491_6;

Selector_2 s3491_6(wires_872_5[3], addr_872_5, wires_3491_6,addr_3491_6);

wire[3:0] wires_3492_6;

wire[31:0] addr_3492_6;

Selector_2 s3492_6(wires_873_5[0], addr_873_5, wires_3492_6,addr_3492_6);

wire[3:0] wires_3493_6;

wire[31:0] addr_3493_6;

Selector_2 s3493_6(wires_873_5[1], addr_873_5, wires_3493_6,addr_3493_6);

wire[3:0] wires_3494_6;

wire[31:0] addr_3494_6;

Selector_2 s3494_6(wires_873_5[2], addr_873_5, wires_3494_6,addr_3494_6);

wire[3:0] wires_3495_6;

wire[31:0] addr_3495_6;

Selector_2 s3495_6(wires_873_5[3], addr_873_5, wires_3495_6,addr_3495_6);

wire[3:0] wires_3496_6;

wire[31:0] addr_3496_6;

Selector_2 s3496_6(wires_874_5[0], addr_874_5, wires_3496_6,addr_3496_6);

wire[3:0] wires_3497_6;

wire[31:0] addr_3497_6;

Selector_2 s3497_6(wires_874_5[1], addr_874_5, wires_3497_6,addr_3497_6);

wire[3:0] wires_3498_6;

wire[31:0] addr_3498_6;

Selector_2 s3498_6(wires_874_5[2], addr_874_5, wires_3498_6,addr_3498_6);

wire[3:0] wires_3499_6;

wire[31:0] addr_3499_6;

Selector_2 s3499_6(wires_874_5[3], addr_874_5, wires_3499_6,addr_3499_6);

wire[3:0] wires_3500_6;

wire[31:0] addr_3500_6;

Selector_2 s3500_6(wires_875_5[0], addr_875_5, wires_3500_6,addr_3500_6);

wire[3:0] wires_3501_6;

wire[31:0] addr_3501_6;

Selector_2 s3501_6(wires_875_5[1], addr_875_5, wires_3501_6,addr_3501_6);

wire[3:0] wires_3502_6;

wire[31:0] addr_3502_6;

Selector_2 s3502_6(wires_875_5[2], addr_875_5, wires_3502_6,addr_3502_6);

wire[3:0] wires_3503_6;

wire[31:0] addr_3503_6;

Selector_2 s3503_6(wires_875_5[3], addr_875_5, wires_3503_6,addr_3503_6);

wire[3:0] wires_3504_6;

wire[31:0] addr_3504_6;

Selector_2 s3504_6(wires_876_5[0], addr_876_5, wires_3504_6,addr_3504_6);

wire[3:0] wires_3505_6;

wire[31:0] addr_3505_6;

Selector_2 s3505_6(wires_876_5[1], addr_876_5, wires_3505_6,addr_3505_6);

wire[3:0] wires_3506_6;

wire[31:0] addr_3506_6;

Selector_2 s3506_6(wires_876_5[2], addr_876_5, wires_3506_6,addr_3506_6);

wire[3:0] wires_3507_6;

wire[31:0] addr_3507_6;

Selector_2 s3507_6(wires_876_5[3], addr_876_5, wires_3507_6,addr_3507_6);

wire[3:0] wires_3508_6;

wire[31:0] addr_3508_6;

Selector_2 s3508_6(wires_877_5[0], addr_877_5, wires_3508_6,addr_3508_6);

wire[3:0] wires_3509_6;

wire[31:0] addr_3509_6;

Selector_2 s3509_6(wires_877_5[1], addr_877_5, wires_3509_6,addr_3509_6);

wire[3:0] wires_3510_6;

wire[31:0] addr_3510_6;

Selector_2 s3510_6(wires_877_5[2], addr_877_5, wires_3510_6,addr_3510_6);

wire[3:0] wires_3511_6;

wire[31:0] addr_3511_6;

Selector_2 s3511_6(wires_877_5[3], addr_877_5, wires_3511_6,addr_3511_6);

wire[3:0] wires_3512_6;

wire[31:0] addr_3512_6;

Selector_2 s3512_6(wires_878_5[0], addr_878_5, wires_3512_6,addr_3512_6);

wire[3:0] wires_3513_6;

wire[31:0] addr_3513_6;

Selector_2 s3513_6(wires_878_5[1], addr_878_5, wires_3513_6,addr_3513_6);

wire[3:0] wires_3514_6;

wire[31:0] addr_3514_6;

Selector_2 s3514_6(wires_878_5[2], addr_878_5, wires_3514_6,addr_3514_6);

wire[3:0] wires_3515_6;

wire[31:0] addr_3515_6;

Selector_2 s3515_6(wires_878_5[3], addr_878_5, wires_3515_6,addr_3515_6);

wire[3:0] wires_3516_6;

wire[31:0] addr_3516_6;

Selector_2 s3516_6(wires_879_5[0], addr_879_5, wires_3516_6,addr_3516_6);

wire[3:0] wires_3517_6;

wire[31:0] addr_3517_6;

Selector_2 s3517_6(wires_879_5[1], addr_879_5, wires_3517_6,addr_3517_6);

wire[3:0] wires_3518_6;

wire[31:0] addr_3518_6;

Selector_2 s3518_6(wires_879_5[2], addr_879_5, wires_3518_6,addr_3518_6);

wire[3:0] wires_3519_6;

wire[31:0] addr_3519_6;

Selector_2 s3519_6(wires_879_5[3], addr_879_5, wires_3519_6,addr_3519_6);

wire[3:0] wires_3520_6;

wire[31:0] addr_3520_6;

Selector_2 s3520_6(wires_880_5[0], addr_880_5, wires_3520_6,addr_3520_6);

wire[3:0] wires_3521_6;

wire[31:0] addr_3521_6;

Selector_2 s3521_6(wires_880_5[1], addr_880_5, wires_3521_6,addr_3521_6);

wire[3:0] wires_3522_6;

wire[31:0] addr_3522_6;

Selector_2 s3522_6(wires_880_5[2], addr_880_5, wires_3522_6,addr_3522_6);

wire[3:0] wires_3523_6;

wire[31:0] addr_3523_6;

Selector_2 s3523_6(wires_880_5[3], addr_880_5, wires_3523_6,addr_3523_6);

wire[3:0] wires_3524_6;

wire[31:0] addr_3524_6;

Selector_2 s3524_6(wires_881_5[0], addr_881_5, wires_3524_6,addr_3524_6);

wire[3:0] wires_3525_6;

wire[31:0] addr_3525_6;

Selector_2 s3525_6(wires_881_5[1], addr_881_5, wires_3525_6,addr_3525_6);

wire[3:0] wires_3526_6;

wire[31:0] addr_3526_6;

Selector_2 s3526_6(wires_881_5[2], addr_881_5, wires_3526_6,addr_3526_6);

wire[3:0] wires_3527_6;

wire[31:0] addr_3527_6;

Selector_2 s3527_6(wires_881_5[3], addr_881_5, wires_3527_6,addr_3527_6);

wire[3:0] wires_3528_6;

wire[31:0] addr_3528_6;

Selector_2 s3528_6(wires_882_5[0], addr_882_5, wires_3528_6,addr_3528_6);

wire[3:0] wires_3529_6;

wire[31:0] addr_3529_6;

Selector_2 s3529_6(wires_882_5[1], addr_882_5, wires_3529_6,addr_3529_6);

wire[3:0] wires_3530_6;

wire[31:0] addr_3530_6;

Selector_2 s3530_6(wires_882_5[2], addr_882_5, wires_3530_6,addr_3530_6);

wire[3:0] wires_3531_6;

wire[31:0] addr_3531_6;

Selector_2 s3531_6(wires_882_5[3], addr_882_5, wires_3531_6,addr_3531_6);

wire[3:0] wires_3532_6;

wire[31:0] addr_3532_6;

Selector_2 s3532_6(wires_883_5[0], addr_883_5, wires_3532_6,addr_3532_6);

wire[3:0] wires_3533_6;

wire[31:0] addr_3533_6;

Selector_2 s3533_6(wires_883_5[1], addr_883_5, wires_3533_6,addr_3533_6);

wire[3:0] wires_3534_6;

wire[31:0] addr_3534_6;

Selector_2 s3534_6(wires_883_5[2], addr_883_5, wires_3534_6,addr_3534_6);

wire[3:0] wires_3535_6;

wire[31:0] addr_3535_6;

Selector_2 s3535_6(wires_883_5[3], addr_883_5, wires_3535_6,addr_3535_6);

wire[3:0] wires_3536_6;

wire[31:0] addr_3536_6;

Selector_2 s3536_6(wires_884_5[0], addr_884_5, wires_3536_6,addr_3536_6);

wire[3:0] wires_3537_6;

wire[31:0] addr_3537_6;

Selector_2 s3537_6(wires_884_5[1], addr_884_5, wires_3537_6,addr_3537_6);

wire[3:0] wires_3538_6;

wire[31:0] addr_3538_6;

Selector_2 s3538_6(wires_884_5[2], addr_884_5, wires_3538_6,addr_3538_6);

wire[3:0] wires_3539_6;

wire[31:0] addr_3539_6;

Selector_2 s3539_6(wires_884_5[3], addr_884_5, wires_3539_6,addr_3539_6);

wire[3:0] wires_3540_6;

wire[31:0] addr_3540_6;

Selector_2 s3540_6(wires_885_5[0], addr_885_5, wires_3540_6,addr_3540_6);

wire[3:0] wires_3541_6;

wire[31:0] addr_3541_6;

Selector_2 s3541_6(wires_885_5[1], addr_885_5, wires_3541_6,addr_3541_6);

wire[3:0] wires_3542_6;

wire[31:0] addr_3542_6;

Selector_2 s3542_6(wires_885_5[2], addr_885_5, wires_3542_6,addr_3542_6);

wire[3:0] wires_3543_6;

wire[31:0] addr_3543_6;

Selector_2 s3543_6(wires_885_5[3], addr_885_5, wires_3543_6,addr_3543_6);

wire[3:0] wires_3544_6;

wire[31:0] addr_3544_6;

Selector_2 s3544_6(wires_886_5[0], addr_886_5, wires_3544_6,addr_3544_6);

wire[3:0] wires_3545_6;

wire[31:0] addr_3545_6;

Selector_2 s3545_6(wires_886_5[1], addr_886_5, wires_3545_6,addr_3545_6);

wire[3:0] wires_3546_6;

wire[31:0] addr_3546_6;

Selector_2 s3546_6(wires_886_5[2], addr_886_5, wires_3546_6,addr_3546_6);

wire[3:0] wires_3547_6;

wire[31:0] addr_3547_6;

Selector_2 s3547_6(wires_886_5[3], addr_886_5, wires_3547_6,addr_3547_6);

wire[3:0] wires_3548_6;

wire[31:0] addr_3548_6;

Selector_2 s3548_6(wires_887_5[0], addr_887_5, wires_3548_6,addr_3548_6);

wire[3:0] wires_3549_6;

wire[31:0] addr_3549_6;

Selector_2 s3549_6(wires_887_5[1], addr_887_5, wires_3549_6,addr_3549_6);

wire[3:0] wires_3550_6;

wire[31:0] addr_3550_6;

Selector_2 s3550_6(wires_887_5[2], addr_887_5, wires_3550_6,addr_3550_6);

wire[3:0] wires_3551_6;

wire[31:0] addr_3551_6;

Selector_2 s3551_6(wires_887_5[3], addr_887_5, wires_3551_6,addr_3551_6);

wire[3:0] wires_3552_6;

wire[31:0] addr_3552_6;

Selector_2 s3552_6(wires_888_5[0], addr_888_5, wires_3552_6,addr_3552_6);

wire[3:0] wires_3553_6;

wire[31:0] addr_3553_6;

Selector_2 s3553_6(wires_888_5[1], addr_888_5, wires_3553_6,addr_3553_6);

wire[3:0] wires_3554_6;

wire[31:0] addr_3554_6;

Selector_2 s3554_6(wires_888_5[2], addr_888_5, wires_3554_6,addr_3554_6);

wire[3:0] wires_3555_6;

wire[31:0] addr_3555_6;

Selector_2 s3555_6(wires_888_5[3], addr_888_5, wires_3555_6,addr_3555_6);

wire[3:0] wires_3556_6;

wire[31:0] addr_3556_6;

Selector_2 s3556_6(wires_889_5[0], addr_889_5, wires_3556_6,addr_3556_6);

wire[3:0] wires_3557_6;

wire[31:0] addr_3557_6;

Selector_2 s3557_6(wires_889_5[1], addr_889_5, wires_3557_6,addr_3557_6);

wire[3:0] wires_3558_6;

wire[31:0] addr_3558_6;

Selector_2 s3558_6(wires_889_5[2], addr_889_5, wires_3558_6,addr_3558_6);

wire[3:0] wires_3559_6;

wire[31:0] addr_3559_6;

Selector_2 s3559_6(wires_889_5[3], addr_889_5, wires_3559_6,addr_3559_6);

wire[3:0] wires_3560_6;

wire[31:0] addr_3560_6;

Selector_2 s3560_6(wires_890_5[0], addr_890_5, wires_3560_6,addr_3560_6);

wire[3:0] wires_3561_6;

wire[31:0] addr_3561_6;

Selector_2 s3561_6(wires_890_5[1], addr_890_5, wires_3561_6,addr_3561_6);

wire[3:0] wires_3562_6;

wire[31:0] addr_3562_6;

Selector_2 s3562_6(wires_890_5[2], addr_890_5, wires_3562_6,addr_3562_6);

wire[3:0] wires_3563_6;

wire[31:0] addr_3563_6;

Selector_2 s3563_6(wires_890_5[3], addr_890_5, wires_3563_6,addr_3563_6);

wire[3:0] wires_3564_6;

wire[31:0] addr_3564_6;

Selector_2 s3564_6(wires_891_5[0], addr_891_5, wires_3564_6,addr_3564_6);

wire[3:0] wires_3565_6;

wire[31:0] addr_3565_6;

Selector_2 s3565_6(wires_891_5[1], addr_891_5, wires_3565_6,addr_3565_6);

wire[3:0] wires_3566_6;

wire[31:0] addr_3566_6;

Selector_2 s3566_6(wires_891_5[2], addr_891_5, wires_3566_6,addr_3566_6);

wire[3:0] wires_3567_6;

wire[31:0] addr_3567_6;

Selector_2 s3567_6(wires_891_5[3], addr_891_5, wires_3567_6,addr_3567_6);

wire[3:0] wires_3568_6;

wire[31:0] addr_3568_6;

Selector_2 s3568_6(wires_892_5[0], addr_892_5, wires_3568_6,addr_3568_6);

wire[3:0] wires_3569_6;

wire[31:0] addr_3569_6;

Selector_2 s3569_6(wires_892_5[1], addr_892_5, wires_3569_6,addr_3569_6);

wire[3:0] wires_3570_6;

wire[31:0] addr_3570_6;

Selector_2 s3570_6(wires_892_5[2], addr_892_5, wires_3570_6,addr_3570_6);

wire[3:0] wires_3571_6;

wire[31:0] addr_3571_6;

Selector_2 s3571_6(wires_892_5[3], addr_892_5, wires_3571_6,addr_3571_6);

wire[3:0] wires_3572_6;

wire[31:0] addr_3572_6;

Selector_2 s3572_6(wires_893_5[0], addr_893_5, wires_3572_6,addr_3572_6);

wire[3:0] wires_3573_6;

wire[31:0] addr_3573_6;

Selector_2 s3573_6(wires_893_5[1], addr_893_5, wires_3573_6,addr_3573_6);

wire[3:0] wires_3574_6;

wire[31:0] addr_3574_6;

Selector_2 s3574_6(wires_893_5[2], addr_893_5, wires_3574_6,addr_3574_6);

wire[3:0] wires_3575_6;

wire[31:0] addr_3575_6;

Selector_2 s3575_6(wires_893_5[3], addr_893_5, wires_3575_6,addr_3575_6);

wire[3:0] wires_3576_6;

wire[31:0] addr_3576_6;

Selector_2 s3576_6(wires_894_5[0], addr_894_5, wires_3576_6,addr_3576_6);

wire[3:0] wires_3577_6;

wire[31:0] addr_3577_6;

Selector_2 s3577_6(wires_894_5[1], addr_894_5, wires_3577_6,addr_3577_6);

wire[3:0] wires_3578_6;

wire[31:0] addr_3578_6;

Selector_2 s3578_6(wires_894_5[2], addr_894_5, wires_3578_6,addr_3578_6);

wire[3:0] wires_3579_6;

wire[31:0] addr_3579_6;

Selector_2 s3579_6(wires_894_5[3], addr_894_5, wires_3579_6,addr_3579_6);

wire[3:0] wires_3580_6;

wire[31:0] addr_3580_6;

Selector_2 s3580_6(wires_895_5[0], addr_895_5, wires_3580_6,addr_3580_6);

wire[3:0] wires_3581_6;

wire[31:0] addr_3581_6;

Selector_2 s3581_6(wires_895_5[1], addr_895_5, wires_3581_6,addr_3581_6);

wire[3:0] wires_3582_6;

wire[31:0] addr_3582_6;

Selector_2 s3582_6(wires_895_5[2], addr_895_5, wires_3582_6,addr_3582_6);

wire[3:0] wires_3583_6;

wire[31:0] addr_3583_6;

Selector_2 s3583_6(wires_895_5[3], addr_895_5, wires_3583_6,addr_3583_6);

wire[3:0] wires_3584_6;

wire[31:0] addr_3584_6;

Selector_2 s3584_6(wires_896_5[0], addr_896_5, wires_3584_6,addr_3584_6);

wire[3:0] wires_3585_6;

wire[31:0] addr_3585_6;

Selector_2 s3585_6(wires_896_5[1], addr_896_5, wires_3585_6,addr_3585_6);

wire[3:0] wires_3586_6;

wire[31:0] addr_3586_6;

Selector_2 s3586_6(wires_896_5[2], addr_896_5, wires_3586_6,addr_3586_6);

wire[3:0] wires_3587_6;

wire[31:0] addr_3587_6;

Selector_2 s3587_6(wires_896_5[3], addr_896_5, wires_3587_6,addr_3587_6);

wire[3:0] wires_3588_6;

wire[31:0] addr_3588_6;

Selector_2 s3588_6(wires_897_5[0], addr_897_5, wires_3588_6,addr_3588_6);

wire[3:0] wires_3589_6;

wire[31:0] addr_3589_6;

Selector_2 s3589_6(wires_897_5[1], addr_897_5, wires_3589_6,addr_3589_6);

wire[3:0] wires_3590_6;

wire[31:0] addr_3590_6;

Selector_2 s3590_6(wires_897_5[2], addr_897_5, wires_3590_6,addr_3590_6);

wire[3:0] wires_3591_6;

wire[31:0] addr_3591_6;

Selector_2 s3591_6(wires_897_5[3], addr_897_5, wires_3591_6,addr_3591_6);

wire[3:0] wires_3592_6;

wire[31:0] addr_3592_6;

Selector_2 s3592_6(wires_898_5[0], addr_898_5, wires_3592_6,addr_3592_6);

wire[3:0] wires_3593_6;

wire[31:0] addr_3593_6;

Selector_2 s3593_6(wires_898_5[1], addr_898_5, wires_3593_6,addr_3593_6);

wire[3:0] wires_3594_6;

wire[31:0] addr_3594_6;

Selector_2 s3594_6(wires_898_5[2], addr_898_5, wires_3594_6,addr_3594_6);

wire[3:0] wires_3595_6;

wire[31:0] addr_3595_6;

Selector_2 s3595_6(wires_898_5[3], addr_898_5, wires_3595_6,addr_3595_6);

wire[3:0] wires_3596_6;

wire[31:0] addr_3596_6;

Selector_2 s3596_6(wires_899_5[0], addr_899_5, wires_3596_6,addr_3596_6);

wire[3:0] wires_3597_6;

wire[31:0] addr_3597_6;

Selector_2 s3597_6(wires_899_5[1], addr_899_5, wires_3597_6,addr_3597_6);

wire[3:0] wires_3598_6;

wire[31:0] addr_3598_6;

Selector_2 s3598_6(wires_899_5[2], addr_899_5, wires_3598_6,addr_3598_6);

wire[3:0] wires_3599_6;

wire[31:0] addr_3599_6;

Selector_2 s3599_6(wires_899_5[3], addr_899_5, wires_3599_6,addr_3599_6);

wire[3:0] wires_3600_6;

wire[31:0] addr_3600_6;

Selector_2 s3600_6(wires_900_5[0], addr_900_5, wires_3600_6,addr_3600_6);

wire[3:0] wires_3601_6;

wire[31:0] addr_3601_6;

Selector_2 s3601_6(wires_900_5[1], addr_900_5, wires_3601_6,addr_3601_6);

wire[3:0] wires_3602_6;

wire[31:0] addr_3602_6;

Selector_2 s3602_6(wires_900_5[2], addr_900_5, wires_3602_6,addr_3602_6);

wire[3:0] wires_3603_6;

wire[31:0] addr_3603_6;

Selector_2 s3603_6(wires_900_5[3], addr_900_5, wires_3603_6,addr_3603_6);

wire[3:0] wires_3604_6;

wire[31:0] addr_3604_6;

Selector_2 s3604_6(wires_901_5[0], addr_901_5, wires_3604_6,addr_3604_6);

wire[3:0] wires_3605_6;

wire[31:0] addr_3605_6;

Selector_2 s3605_6(wires_901_5[1], addr_901_5, wires_3605_6,addr_3605_6);

wire[3:0] wires_3606_6;

wire[31:0] addr_3606_6;

Selector_2 s3606_6(wires_901_5[2], addr_901_5, wires_3606_6,addr_3606_6);

wire[3:0] wires_3607_6;

wire[31:0] addr_3607_6;

Selector_2 s3607_6(wires_901_5[3], addr_901_5, wires_3607_6,addr_3607_6);

wire[3:0] wires_3608_6;

wire[31:0] addr_3608_6;

Selector_2 s3608_6(wires_902_5[0], addr_902_5, wires_3608_6,addr_3608_6);

wire[3:0] wires_3609_6;

wire[31:0] addr_3609_6;

Selector_2 s3609_6(wires_902_5[1], addr_902_5, wires_3609_6,addr_3609_6);

wire[3:0] wires_3610_6;

wire[31:0] addr_3610_6;

Selector_2 s3610_6(wires_902_5[2], addr_902_5, wires_3610_6,addr_3610_6);

wire[3:0] wires_3611_6;

wire[31:0] addr_3611_6;

Selector_2 s3611_6(wires_902_5[3], addr_902_5, wires_3611_6,addr_3611_6);

wire[3:0] wires_3612_6;

wire[31:0] addr_3612_6;

Selector_2 s3612_6(wires_903_5[0], addr_903_5, wires_3612_6,addr_3612_6);

wire[3:0] wires_3613_6;

wire[31:0] addr_3613_6;

Selector_2 s3613_6(wires_903_5[1], addr_903_5, wires_3613_6,addr_3613_6);

wire[3:0] wires_3614_6;

wire[31:0] addr_3614_6;

Selector_2 s3614_6(wires_903_5[2], addr_903_5, wires_3614_6,addr_3614_6);

wire[3:0] wires_3615_6;

wire[31:0] addr_3615_6;

Selector_2 s3615_6(wires_903_5[3], addr_903_5, wires_3615_6,addr_3615_6);

wire[3:0] wires_3616_6;

wire[31:0] addr_3616_6;

Selector_2 s3616_6(wires_904_5[0], addr_904_5, wires_3616_6,addr_3616_6);

wire[3:0] wires_3617_6;

wire[31:0] addr_3617_6;

Selector_2 s3617_6(wires_904_5[1], addr_904_5, wires_3617_6,addr_3617_6);

wire[3:0] wires_3618_6;

wire[31:0] addr_3618_6;

Selector_2 s3618_6(wires_904_5[2], addr_904_5, wires_3618_6,addr_3618_6);

wire[3:0] wires_3619_6;

wire[31:0] addr_3619_6;

Selector_2 s3619_6(wires_904_5[3], addr_904_5, wires_3619_6,addr_3619_6);

wire[3:0] wires_3620_6;

wire[31:0] addr_3620_6;

Selector_2 s3620_6(wires_905_5[0], addr_905_5, wires_3620_6,addr_3620_6);

wire[3:0] wires_3621_6;

wire[31:0] addr_3621_6;

Selector_2 s3621_6(wires_905_5[1], addr_905_5, wires_3621_6,addr_3621_6);

wire[3:0] wires_3622_6;

wire[31:0] addr_3622_6;

Selector_2 s3622_6(wires_905_5[2], addr_905_5, wires_3622_6,addr_3622_6);

wire[3:0] wires_3623_6;

wire[31:0] addr_3623_6;

Selector_2 s3623_6(wires_905_5[3], addr_905_5, wires_3623_6,addr_3623_6);

wire[3:0] wires_3624_6;

wire[31:0] addr_3624_6;

Selector_2 s3624_6(wires_906_5[0], addr_906_5, wires_3624_6,addr_3624_6);

wire[3:0] wires_3625_6;

wire[31:0] addr_3625_6;

Selector_2 s3625_6(wires_906_5[1], addr_906_5, wires_3625_6,addr_3625_6);

wire[3:0] wires_3626_6;

wire[31:0] addr_3626_6;

Selector_2 s3626_6(wires_906_5[2], addr_906_5, wires_3626_6,addr_3626_6);

wire[3:0] wires_3627_6;

wire[31:0] addr_3627_6;

Selector_2 s3627_6(wires_906_5[3], addr_906_5, wires_3627_6,addr_3627_6);

wire[3:0] wires_3628_6;

wire[31:0] addr_3628_6;

Selector_2 s3628_6(wires_907_5[0], addr_907_5, wires_3628_6,addr_3628_6);

wire[3:0] wires_3629_6;

wire[31:0] addr_3629_6;

Selector_2 s3629_6(wires_907_5[1], addr_907_5, wires_3629_6,addr_3629_6);

wire[3:0] wires_3630_6;

wire[31:0] addr_3630_6;

Selector_2 s3630_6(wires_907_5[2], addr_907_5, wires_3630_6,addr_3630_6);

wire[3:0] wires_3631_6;

wire[31:0] addr_3631_6;

Selector_2 s3631_6(wires_907_5[3], addr_907_5, wires_3631_6,addr_3631_6);

wire[3:0] wires_3632_6;

wire[31:0] addr_3632_6;

Selector_2 s3632_6(wires_908_5[0], addr_908_5, wires_3632_6,addr_3632_6);

wire[3:0] wires_3633_6;

wire[31:0] addr_3633_6;

Selector_2 s3633_6(wires_908_5[1], addr_908_5, wires_3633_6,addr_3633_6);

wire[3:0] wires_3634_6;

wire[31:0] addr_3634_6;

Selector_2 s3634_6(wires_908_5[2], addr_908_5, wires_3634_6,addr_3634_6);

wire[3:0] wires_3635_6;

wire[31:0] addr_3635_6;

Selector_2 s3635_6(wires_908_5[3], addr_908_5, wires_3635_6,addr_3635_6);

wire[3:0] wires_3636_6;

wire[31:0] addr_3636_6;

Selector_2 s3636_6(wires_909_5[0], addr_909_5, wires_3636_6,addr_3636_6);

wire[3:0] wires_3637_6;

wire[31:0] addr_3637_6;

Selector_2 s3637_6(wires_909_5[1], addr_909_5, wires_3637_6,addr_3637_6);

wire[3:0] wires_3638_6;

wire[31:0] addr_3638_6;

Selector_2 s3638_6(wires_909_5[2], addr_909_5, wires_3638_6,addr_3638_6);

wire[3:0] wires_3639_6;

wire[31:0] addr_3639_6;

Selector_2 s3639_6(wires_909_5[3], addr_909_5, wires_3639_6,addr_3639_6);

wire[3:0] wires_3640_6;

wire[31:0] addr_3640_6;

Selector_2 s3640_6(wires_910_5[0], addr_910_5, wires_3640_6,addr_3640_6);

wire[3:0] wires_3641_6;

wire[31:0] addr_3641_6;

Selector_2 s3641_6(wires_910_5[1], addr_910_5, wires_3641_6,addr_3641_6);

wire[3:0] wires_3642_6;

wire[31:0] addr_3642_6;

Selector_2 s3642_6(wires_910_5[2], addr_910_5, wires_3642_6,addr_3642_6);

wire[3:0] wires_3643_6;

wire[31:0] addr_3643_6;

Selector_2 s3643_6(wires_910_5[3], addr_910_5, wires_3643_6,addr_3643_6);

wire[3:0] wires_3644_6;

wire[31:0] addr_3644_6;

Selector_2 s3644_6(wires_911_5[0], addr_911_5, wires_3644_6,addr_3644_6);

wire[3:0] wires_3645_6;

wire[31:0] addr_3645_6;

Selector_2 s3645_6(wires_911_5[1], addr_911_5, wires_3645_6,addr_3645_6);

wire[3:0] wires_3646_6;

wire[31:0] addr_3646_6;

Selector_2 s3646_6(wires_911_5[2], addr_911_5, wires_3646_6,addr_3646_6);

wire[3:0] wires_3647_6;

wire[31:0] addr_3647_6;

Selector_2 s3647_6(wires_911_5[3], addr_911_5, wires_3647_6,addr_3647_6);

wire[3:0] wires_3648_6;

wire[31:0] addr_3648_6;

Selector_2 s3648_6(wires_912_5[0], addr_912_5, wires_3648_6,addr_3648_6);

wire[3:0] wires_3649_6;

wire[31:0] addr_3649_6;

Selector_2 s3649_6(wires_912_5[1], addr_912_5, wires_3649_6,addr_3649_6);

wire[3:0] wires_3650_6;

wire[31:0] addr_3650_6;

Selector_2 s3650_6(wires_912_5[2], addr_912_5, wires_3650_6,addr_3650_6);

wire[3:0] wires_3651_6;

wire[31:0] addr_3651_6;

Selector_2 s3651_6(wires_912_5[3], addr_912_5, wires_3651_6,addr_3651_6);

wire[3:0] wires_3652_6;

wire[31:0] addr_3652_6;

Selector_2 s3652_6(wires_913_5[0], addr_913_5, wires_3652_6,addr_3652_6);

wire[3:0] wires_3653_6;

wire[31:0] addr_3653_6;

Selector_2 s3653_6(wires_913_5[1], addr_913_5, wires_3653_6,addr_3653_6);

wire[3:0] wires_3654_6;

wire[31:0] addr_3654_6;

Selector_2 s3654_6(wires_913_5[2], addr_913_5, wires_3654_6,addr_3654_6);

wire[3:0] wires_3655_6;

wire[31:0] addr_3655_6;

Selector_2 s3655_6(wires_913_5[3], addr_913_5, wires_3655_6,addr_3655_6);

wire[3:0] wires_3656_6;

wire[31:0] addr_3656_6;

Selector_2 s3656_6(wires_914_5[0], addr_914_5, wires_3656_6,addr_3656_6);

wire[3:0] wires_3657_6;

wire[31:0] addr_3657_6;

Selector_2 s3657_6(wires_914_5[1], addr_914_5, wires_3657_6,addr_3657_6);

wire[3:0] wires_3658_6;

wire[31:0] addr_3658_6;

Selector_2 s3658_6(wires_914_5[2], addr_914_5, wires_3658_6,addr_3658_6);

wire[3:0] wires_3659_6;

wire[31:0] addr_3659_6;

Selector_2 s3659_6(wires_914_5[3], addr_914_5, wires_3659_6,addr_3659_6);

wire[3:0] wires_3660_6;

wire[31:0] addr_3660_6;

Selector_2 s3660_6(wires_915_5[0], addr_915_5, wires_3660_6,addr_3660_6);

wire[3:0] wires_3661_6;

wire[31:0] addr_3661_6;

Selector_2 s3661_6(wires_915_5[1], addr_915_5, wires_3661_6,addr_3661_6);

wire[3:0] wires_3662_6;

wire[31:0] addr_3662_6;

Selector_2 s3662_6(wires_915_5[2], addr_915_5, wires_3662_6,addr_3662_6);

wire[3:0] wires_3663_6;

wire[31:0] addr_3663_6;

Selector_2 s3663_6(wires_915_5[3], addr_915_5, wires_3663_6,addr_3663_6);

wire[3:0] wires_3664_6;

wire[31:0] addr_3664_6;

Selector_2 s3664_6(wires_916_5[0], addr_916_5, wires_3664_6,addr_3664_6);

wire[3:0] wires_3665_6;

wire[31:0] addr_3665_6;

Selector_2 s3665_6(wires_916_5[1], addr_916_5, wires_3665_6,addr_3665_6);

wire[3:0] wires_3666_6;

wire[31:0] addr_3666_6;

Selector_2 s3666_6(wires_916_5[2], addr_916_5, wires_3666_6,addr_3666_6);

wire[3:0] wires_3667_6;

wire[31:0] addr_3667_6;

Selector_2 s3667_6(wires_916_5[3], addr_916_5, wires_3667_6,addr_3667_6);

wire[3:0] wires_3668_6;

wire[31:0] addr_3668_6;

Selector_2 s3668_6(wires_917_5[0], addr_917_5, wires_3668_6,addr_3668_6);

wire[3:0] wires_3669_6;

wire[31:0] addr_3669_6;

Selector_2 s3669_6(wires_917_5[1], addr_917_5, wires_3669_6,addr_3669_6);

wire[3:0] wires_3670_6;

wire[31:0] addr_3670_6;

Selector_2 s3670_6(wires_917_5[2], addr_917_5, wires_3670_6,addr_3670_6);

wire[3:0] wires_3671_6;

wire[31:0] addr_3671_6;

Selector_2 s3671_6(wires_917_5[3], addr_917_5, wires_3671_6,addr_3671_6);

wire[3:0] wires_3672_6;

wire[31:0] addr_3672_6;

Selector_2 s3672_6(wires_918_5[0], addr_918_5, wires_3672_6,addr_3672_6);

wire[3:0] wires_3673_6;

wire[31:0] addr_3673_6;

Selector_2 s3673_6(wires_918_5[1], addr_918_5, wires_3673_6,addr_3673_6);

wire[3:0] wires_3674_6;

wire[31:0] addr_3674_6;

Selector_2 s3674_6(wires_918_5[2], addr_918_5, wires_3674_6,addr_3674_6);

wire[3:0] wires_3675_6;

wire[31:0] addr_3675_6;

Selector_2 s3675_6(wires_918_5[3], addr_918_5, wires_3675_6,addr_3675_6);

wire[3:0] wires_3676_6;

wire[31:0] addr_3676_6;

Selector_2 s3676_6(wires_919_5[0], addr_919_5, wires_3676_6,addr_3676_6);

wire[3:0] wires_3677_6;

wire[31:0] addr_3677_6;

Selector_2 s3677_6(wires_919_5[1], addr_919_5, wires_3677_6,addr_3677_6);

wire[3:0] wires_3678_6;

wire[31:0] addr_3678_6;

Selector_2 s3678_6(wires_919_5[2], addr_919_5, wires_3678_6,addr_3678_6);

wire[3:0] wires_3679_6;

wire[31:0] addr_3679_6;

Selector_2 s3679_6(wires_919_5[3], addr_919_5, wires_3679_6,addr_3679_6);

wire[3:0] wires_3680_6;

wire[31:0] addr_3680_6;

Selector_2 s3680_6(wires_920_5[0], addr_920_5, wires_3680_6,addr_3680_6);

wire[3:0] wires_3681_6;

wire[31:0] addr_3681_6;

Selector_2 s3681_6(wires_920_5[1], addr_920_5, wires_3681_6,addr_3681_6);

wire[3:0] wires_3682_6;

wire[31:0] addr_3682_6;

Selector_2 s3682_6(wires_920_5[2], addr_920_5, wires_3682_6,addr_3682_6);

wire[3:0] wires_3683_6;

wire[31:0] addr_3683_6;

Selector_2 s3683_6(wires_920_5[3], addr_920_5, wires_3683_6,addr_3683_6);

wire[3:0] wires_3684_6;

wire[31:0] addr_3684_6;

Selector_2 s3684_6(wires_921_5[0], addr_921_5, wires_3684_6,addr_3684_6);

wire[3:0] wires_3685_6;

wire[31:0] addr_3685_6;

Selector_2 s3685_6(wires_921_5[1], addr_921_5, wires_3685_6,addr_3685_6);

wire[3:0] wires_3686_6;

wire[31:0] addr_3686_6;

Selector_2 s3686_6(wires_921_5[2], addr_921_5, wires_3686_6,addr_3686_6);

wire[3:0] wires_3687_6;

wire[31:0] addr_3687_6;

Selector_2 s3687_6(wires_921_5[3], addr_921_5, wires_3687_6,addr_3687_6);

wire[3:0] wires_3688_6;

wire[31:0] addr_3688_6;

Selector_2 s3688_6(wires_922_5[0], addr_922_5, wires_3688_6,addr_3688_6);

wire[3:0] wires_3689_6;

wire[31:0] addr_3689_6;

Selector_2 s3689_6(wires_922_5[1], addr_922_5, wires_3689_6,addr_3689_6);

wire[3:0] wires_3690_6;

wire[31:0] addr_3690_6;

Selector_2 s3690_6(wires_922_5[2], addr_922_5, wires_3690_6,addr_3690_6);

wire[3:0] wires_3691_6;

wire[31:0] addr_3691_6;

Selector_2 s3691_6(wires_922_5[3], addr_922_5, wires_3691_6,addr_3691_6);

wire[3:0] wires_3692_6;

wire[31:0] addr_3692_6;

Selector_2 s3692_6(wires_923_5[0], addr_923_5, wires_3692_6,addr_3692_6);

wire[3:0] wires_3693_6;

wire[31:0] addr_3693_6;

Selector_2 s3693_6(wires_923_5[1], addr_923_5, wires_3693_6,addr_3693_6);

wire[3:0] wires_3694_6;

wire[31:0] addr_3694_6;

Selector_2 s3694_6(wires_923_5[2], addr_923_5, wires_3694_6,addr_3694_6);

wire[3:0] wires_3695_6;

wire[31:0] addr_3695_6;

Selector_2 s3695_6(wires_923_5[3], addr_923_5, wires_3695_6,addr_3695_6);

wire[3:0] wires_3696_6;

wire[31:0] addr_3696_6;

Selector_2 s3696_6(wires_924_5[0], addr_924_5, wires_3696_6,addr_3696_6);

wire[3:0] wires_3697_6;

wire[31:0] addr_3697_6;

Selector_2 s3697_6(wires_924_5[1], addr_924_5, wires_3697_6,addr_3697_6);

wire[3:0] wires_3698_6;

wire[31:0] addr_3698_6;

Selector_2 s3698_6(wires_924_5[2], addr_924_5, wires_3698_6,addr_3698_6);

wire[3:0] wires_3699_6;

wire[31:0] addr_3699_6;

Selector_2 s3699_6(wires_924_5[3], addr_924_5, wires_3699_6,addr_3699_6);

wire[3:0] wires_3700_6;

wire[31:0] addr_3700_6;

Selector_2 s3700_6(wires_925_5[0], addr_925_5, wires_3700_6,addr_3700_6);

wire[3:0] wires_3701_6;

wire[31:0] addr_3701_6;

Selector_2 s3701_6(wires_925_5[1], addr_925_5, wires_3701_6,addr_3701_6);

wire[3:0] wires_3702_6;

wire[31:0] addr_3702_6;

Selector_2 s3702_6(wires_925_5[2], addr_925_5, wires_3702_6,addr_3702_6);

wire[3:0] wires_3703_6;

wire[31:0] addr_3703_6;

Selector_2 s3703_6(wires_925_5[3], addr_925_5, wires_3703_6,addr_3703_6);

wire[3:0] wires_3704_6;

wire[31:0] addr_3704_6;

Selector_2 s3704_6(wires_926_5[0], addr_926_5, wires_3704_6,addr_3704_6);

wire[3:0] wires_3705_6;

wire[31:0] addr_3705_6;

Selector_2 s3705_6(wires_926_5[1], addr_926_5, wires_3705_6,addr_3705_6);

wire[3:0] wires_3706_6;

wire[31:0] addr_3706_6;

Selector_2 s3706_6(wires_926_5[2], addr_926_5, wires_3706_6,addr_3706_6);

wire[3:0] wires_3707_6;

wire[31:0] addr_3707_6;

Selector_2 s3707_6(wires_926_5[3], addr_926_5, wires_3707_6,addr_3707_6);

wire[3:0] wires_3708_6;

wire[31:0] addr_3708_6;

Selector_2 s3708_6(wires_927_5[0], addr_927_5, wires_3708_6,addr_3708_6);

wire[3:0] wires_3709_6;

wire[31:0] addr_3709_6;

Selector_2 s3709_6(wires_927_5[1], addr_927_5, wires_3709_6,addr_3709_6);

wire[3:0] wires_3710_6;

wire[31:0] addr_3710_6;

Selector_2 s3710_6(wires_927_5[2], addr_927_5, wires_3710_6,addr_3710_6);

wire[3:0] wires_3711_6;

wire[31:0] addr_3711_6;

Selector_2 s3711_6(wires_927_5[3], addr_927_5, wires_3711_6,addr_3711_6);

wire[3:0] wires_3712_6;

wire[31:0] addr_3712_6;

Selector_2 s3712_6(wires_928_5[0], addr_928_5, wires_3712_6,addr_3712_6);

wire[3:0] wires_3713_6;

wire[31:0] addr_3713_6;

Selector_2 s3713_6(wires_928_5[1], addr_928_5, wires_3713_6,addr_3713_6);

wire[3:0] wires_3714_6;

wire[31:0] addr_3714_6;

Selector_2 s3714_6(wires_928_5[2], addr_928_5, wires_3714_6,addr_3714_6);

wire[3:0] wires_3715_6;

wire[31:0] addr_3715_6;

Selector_2 s3715_6(wires_928_5[3], addr_928_5, wires_3715_6,addr_3715_6);

wire[3:0] wires_3716_6;

wire[31:0] addr_3716_6;

Selector_2 s3716_6(wires_929_5[0], addr_929_5, wires_3716_6,addr_3716_6);

wire[3:0] wires_3717_6;

wire[31:0] addr_3717_6;

Selector_2 s3717_6(wires_929_5[1], addr_929_5, wires_3717_6,addr_3717_6);

wire[3:0] wires_3718_6;

wire[31:0] addr_3718_6;

Selector_2 s3718_6(wires_929_5[2], addr_929_5, wires_3718_6,addr_3718_6);

wire[3:0] wires_3719_6;

wire[31:0] addr_3719_6;

Selector_2 s3719_6(wires_929_5[3], addr_929_5, wires_3719_6,addr_3719_6);

wire[3:0] wires_3720_6;

wire[31:0] addr_3720_6;

Selector_2 s3720_6(wires_930_5[0], addr_930_5, wires_3720_6,addr_3720_6);

wire[3:0] wires_3721_6;

wire[31:0] addr_3721_6;

Selector_2 s3721_6(wires_930_5[1], addr_930_5, wires_3721_6,addr_3721_6);

wire[3:0] wires_3722_6;

wire[31:0] addr_3722_6;

Selector_2 s3722_6(wires_930_5[2], addr_930_5, wires_3722_6,addr_3722_6);

wire[3:0] wires_3723_6;

wire[31:0] addr_3723_6;

Selector_2 s3723_6(wires_930_5[3], addr_930_5, wires_3723_6,addr_3723_6);

wire[3:0] wires_3724_6;

wire[31:0] addr_3724_6;

Selector_2 s3724_6(wires_931_5[0], addr_931_5, wires_3724_6,addr_3724_6);

wire[3:0] wires_3725_6;

wire[31:0] addr_3725_6;

Selector_2 s3725_6(wires_931_5[1], addr_931_5, wires_3725_6,addr_3725_6);

wire[3:0] wires_3726_6;

wire[31:0] addr_3726_6;

Selector_2 s3726_6(wires_931_5[2], addr_931_5, wires_3726_6,addr_3726_6);

wire[3:0] wires_3727_6;

wire[31:0] addr_3727_6;

Selector_2 s3727_6(wires_931_5[3], addr_931_5, wires_3727_6,addr_3727_6);

wire[3:0] wires_3728_6;

wire[31:0] addr_3728_6;

Selector_2 s3728_6(wires_932_5[0], addr_932_5, wires_3728_6,addr_3728_6);

wire[3:0] wires_3729_6;

wire[31:0] addr_3729_6;

Selector_2 s3729_6(wires_932_5[1], addr_932_5, wires_3729_6,addr_3729_6);

wire[3:0] wires_3730_6;

wire[31:0] addr_3730_6;

Selector_2 s3730_6(wires_932_5[2], addr_932_5, wires_3730_6,addr_3730_6);

wire[3:0] wires_3731_6;

wire[31:0] addr_3731_6;

Selector_2 s3731_6(wires_932_5[3], addr_932_5, wires_3731_6,addr_3731_6);

wire[3:0] wires_3732_6;

wire[31:0] addr_3732_6;

Selector_2 s3732_6(wires_933_5[0], addr_933_5, wires_3732_6,addr_3732_6);

wire[3:0] wires_3733_6;

wire[31:0] addr_3733_6;

Selector_2 s3733_6(wires_933_5[1], addr_933_5, wires_3733_6,addr_3733_6);

wire[3:0] wires_3734_6;

wire[31:0] addr_3734_6;

Selector_2 s3734_6(wires_933_5[2], addr_933_5, wires_3734_6,addr_3734_6);

wire[3:0] wires_3735_6;

wire[31:0] addr_3735_6;

Selector_2 s3735_6(wires_933_5[3], addr_933_5, wires_3735_6,addr_3735_6);

wire[3:0] wires_3736_6;

wire[31:0] addr_3736_6;

Selector_2 s3736_6(wires_934_5[0], addr_934_5, wires_3736_6,addr_3736_6);

wire[3:0] wires_3737_6;

wire[31:0] addr_3737_6;

Selector_2 s3737_6(wires_934_5[1], addr_934_5, wires_3737_6,addr_3737_6);

wire[3:0] wires_3738_6;

wire[31:0] addr_3738_6;

Selector_2 s3738_6(wires_934_5[2], addr_934_5, wires_3738_6,addr_3738_6);

wire[3:0] wires_3739_6;

wire[31:0] addr_3739_6;

Selector_2 s3739_6(wires_934_5[3], addr_934_5, wires_3739_6,addr_3739_6);

wire[3:0] wires_3740_6;

wire[31:0] addr_3740_6;

Selector_2 s3740_6(wires_935_5[0], addr_935_5, wires_3740_6,addr_3740_6);

wire[3:0] wires_3741_6;

wire[31:0] addr_3741_6;

Selector_2 s3741_6(wires_935_5[1], addr_935_5, wires_3741_6,addr_3741_6);

wire[3:0] wires_3742_6;

wire[31:0] addr_3742_6;

Selector_2 s3742_6(wires_935_5[2], addr_935_5, wires_3742_6,addr_3742_6);

wire[3:0] wires_3743_6;

wire[31:0] addr_3743_6;

Selector_2 s3743_6(wires_935_5[3], addr_935_5, wires_3743_6,addr_3743_6);

wire[3:0] wires_3744_6;

wire[31:0] addr_3744_6;

Selector_2 s3744_6(wires_936_5[0], addr_936_5, wires_3744_6,addr_3744_6);

wire[3:0] wires_3745_6;

wire[31:0] addr_3745_6;

Selector_2 s3745_6(wires_936_5[1], addr_936_5, wires_3745_6,addr_3745_6);

wire[3:0] wires_3746_6;

wire[31:0] addr_3746_6;

Selector_2 s3746_6(wires_936_5[2], addr_936_5, wires_3746_6,addr_3746_6);

wire[3:0] wires_3747_6;

wire[31:0] addr_3747_6;

Selector_2 s3747_6(wires_936_5[3], addr_936_5, wires_3747_6,addr_3747_6);

wire[3:0] wires_3748_6;

wire[31:0] addr_3748_6;

Selector_2 s3748_6(wires_937_5[0], addr_937_5, wires_3748_6,addr_3748_6);

wire[3:0] wires_3749_6;

wire[31:0] addr_3749_6;

Selector_2 s3749_6(wires_937_5[1], addr_937_5, wires_3749_6,addr_3749_6);

wire[3:0] wires_3750_6;

wire[31:0] addr_3750_6;

Selector_2 s3750_6(wires_937_5[2], addr_937_5, wires_3750_6,addr_3750_6);

wire[3:0] wires_3751_6;

wire[31:0] addr_3751_6;

Selector_2 s3751_6(wires_937_5[3], addr_937_5, wires_3751_6,addr_3751_6);

wire[3:0] wires_3752_6;

wire[31:0] addr_3752_6;

Selector_2 s3752_6(wires_938_5[0], addr_938_5, wires_3752_6,addr_3752_6);

wire[3:0] wires_3753_6;

wire[31:0] addr_3753_6;

Selector_2 s3753_6(wires_938_5[1], addr_938_5, wires_3753_6,addr_3753_6);

wire[3:0] wires_3754_6;

wire[31:0] addr_3754_6;

Selector_2 s3754_6(wires_938_5[2], addr_938_5, wires_3754_6,addr_3754_6);

wire[3:0] wires_3755_6;

wire[31:0] addr_3755_6;

Selector_2 s3755_6(wires_938_5[3], addr_938_5, wires_3755_6,addr_3755_6);

wire[3:0] wires_3756_6;

wire[31:0] addr_3756_6;

Selector_2 s3756_6(wires_939_5[0], addr_939_5, wires_3756_6,addr_3756_6);

wire[3:0] wires_3757_6;

wire[31:0] addr_3757_6;

Selector_2 s3757_6(wires_939_5[1], addr_939_5, wires_3757_6,addr_3757_6);

wire[3:0] wires_3758_6;

wire[31:0] addr_3758_6;

Selector_2 s3758_6(wires_939_5[2], addr_939_5, wires_3758_6,addr_3758_6);

wire[3:0] wires_3759_6;

wire[31:0] addr_3759_6;

Selector_2 s3759_6(wires_939_5[3], addr_939_5, wires_3759_6,addr_3759_6);

wire[3:0] wires_3760_6;

wire[31:0] addr_3760_6;

Selector_2 s3760_6(wires_940_5[0], addr_940_5, wires_3760_6,addr_3760_6);

wire[3:0] wires_3761_6;

wire[31:0] addr_3761_6;

Selector_2 s3761_6(wires_940_5[1], addr_940_5, wires_3761_6,addr_3761_6);

wire[3:0] wires_3762_6;

wire[31:0] addr_3762_6;

Selector_2 s3762_6(wires_940_5[2], addr_940_5, wires_3762_6,addr_3762_6);

wire[3:0] wires_3763_6;

wire[31:0] addr_3763_6;

Selector_2 s3763_6(wires_940_5[3], addr_940_5, wires_3763_6,addr_3763_6);

wire[3:0] wires_3764_6;

wire[31:0] addr_3764_6;

Selector_2 s3764_6(wires_941_5[0], addr_941_5, wires_3764_6,addr_3764_6);

wire[3:0] wires_3765_6;

wire[31:0] addr_3765_6;

Selector_2 s3765_6(wires_941_5[1], addr_941_5, wires_3765_6,addr_3765_6);

wire[3:0] wires_3766_6;

wire[31:0] addr_3766_6;

Selector_2 s3766_6(wires_941_5[2], addr_941_5, wires_3766_6,addr_3766_6);

wire[3:0] wires_3767_6;

wire[31:0] addr_3767_6;

Selector_2 s3767_6(wires_941_5[3], addr_941_5, wires_3767_6,addr_3767_6);

wire[3:0] wires_3768_6;

wire[31:0] addr_3768_6;

Selector_2 s3768_6(wires_942_5[0], addr_942_5, wires_3768_6,addr_3768_6);

wire[3:0] wires_3769_6;

wire[31:0] addr_3769_6;

Selector_2 s3769_6(wires_942_5[1], addr_942_5, wires_3769_6,addr_3769_6);

wire[3:0] wires_3770_6;

wire[31:0] addr_3770_6;

Selector_2 s3770_6(wires_942_5[2], addr_942_5, wires_3770_6,addr_3770_6);

wire[3:0] wires_3771_6;

wire[31:0] addr_3771_6;

Selector_2 s3771_6(wires_942_5[3], addr_942_5, wires_3771_6,addr_3771_6);

wire[3:0] wires_3772_6;

wire[31:0] addr_3772_6;

Selector_2 s3772_6(wires_943_5[0], addr_943_5, wires_3772_6,addr_3772_6);

wire[3:0] wires_3773_6;

wire[31:0] addr_3773_6;

Selector_2 s3773_6(wires_943_5[1], addr_943_5, wires_3773_6,addr_3773_6);

wire[3:0] wires_3774_6;

wire[31:0] addr_3774_6;

Selector_2 s3774_6(wires_943_5[2], addr_943_5, wires_3774_6,addr_3774_6);

wire[3:0] wires_3775_6;

wire[31:0] addr_3775_6;

Selector_2 s3775_6(wires_943_5[3], addr_943_5, wires_3775_6,addr_3775_6);

wire[3:0] wires_3776_6;

wire[31:0] addr_3776_6;

Selector_2 s3776_6(wires_944_5[0], addr_944_5, wires_3776_6,addr_3776_6);

wire[3:0] wires_3777_6;

wire[31:0] addr_3777_6;

Selector_2 s3777_6(wires_944_5[1], addr_944_5, wires_3777_6,addr_3777_6);

wire[3:0] wires_3778_6;

wire[31:0] addr_3778_6;

Selector_2 s3778_6(wires_944_5[2], addr_944_5, wires_3778_6,addr_3778_6);

wire[3:0] wires_3779_6;

wire[31:0] addr_3779_6;

Selector_2 s3779_6(wires_944_5[3], addr_944_5, wires_3779_6,addr_3779_6);

wire[3:0] wires_3780_6;

wire[31:0] addr_3780_6;

Selector_2 s3780_6(wires_945_5[0], addr_945_5, wires_3780_6,addr_3780_6);

wire[3:0] wires_3781_6;

wire[31:0] addr_3781_6;

Selector_2 s3781_6(wires_945_5[1], addr_945_5, wires_3781_6,addr_3781_6);

wire[3:0] wires_3782_6;

wire[31:0] addr_3782_6;

Selector_2 s3782_6(wires_945_5[2], addr_945_5, wires_3782_6,addr_3782_6);

wire[3:0] wires_3783_6;

wire[31:0] addr_3783_6;

Selector_2 s3783_6(wires_945_5[3], addr_945_5, wires_3783_6,addr_3783_6);

wire[3:0] wires_3784_6;

wire[31:0] addr_3784_6;

Selector_2 s3784_6(wires_946_5[0], addr_946_5, wires_3784_6,addr_3784_6);

wire[3:0] wires_3785_6;

wire[31:0] addr_3785_6;

Selector_2 s3785_6(wires_946_5[1], addr_946_5, wires_3785_6,addr_3785_6);

wire[3:0] wires_3786_6;

wire[31:0] addr_3786_6;

Selector_2 s3786_6(wires_946_5[2], addr_946_5, wires_3786_6,addr_3786_6);

wire[3:0] wires_3787_6;

wire[31:0] addr_3787_6;

Selector_2 s3787_6(wires_946_5[3], addr_946_5, wires_3787_6,addr_3787_6);

wire[3:0] wires_3788_6;

wire[31:0] addr_3788_6;

Selector_2 s3788_6(wires_947_5[0], addr_947_5, wires_3788_6,addr_3788_6);

wire[3:0] wires_3789_6;

wire[31:0] addr_3789_6;

Selector_2 s3789_6(wires_947_5[1], addr_947_5, wires_3789_6,addr_3789_6);

wire[3:0] wires_3790_6;

wire[31:0] addr_3790_6;

Selector_2 s3790_6(wires_947_5[2], addr_947_5, wires_3790_6,addr_3790_6);

wire[3:0] wires_3791_6;

wire[31:0] addr_3791_6;

Selector_2 s3791_6(wires_947_5[3], addr_947_5, wires_3791_6,addr_3791_6);

wire[3:0] wires_3792_6;

wire[31:0] addr_3792_6;

Selector_2 s3792_6(wires_948_5[0], addr_948_5, wires_3792_6,addr_3792_6);

wire[3:0] wires_3793_6;

wire[31:0] addr_3793_6;

Selector_2 s3793_6(wires_948_5[1], addr_948_5, wires_3793_6,addr_3793_6);

wire[3:0] wires_3794_6;

wire[31:0] addr_3794_6;

Selector_2 s3794_6(wires_948_5[2], addr_948_5, wires_3794_6,addr_3794_6);

wire[3:0] wires_3795_6;

wire[31:0] addr_3795_6;

Selector_2 s3795_6(wires_948_5[3], addr_948_5, wires_3795_6,addr_3795_6);

wire[3:0] wires_3796_6;

wire[31:0] addr_3796_6;

Selector_2 s3796_6(wires_949_5[0], addr_949_5, wires_3796_6,addr_3796_6);

wire[3:0] wires_3797_6;

wire[31:0] addr_3797_6;

Selector_2 s3797_6(wires_949_5[1], addr_949_5, wires_3797_6,addr_3797_6);

wire[3:0] wires_3798_6;

wire[31:0] addr_3798_6;

Selector_2 s3798_6(wires_949_5[2], addr_949_5, wires_3798_6,addr_3798_6);

wire[3:0] wires_3799_6;

wire[31:0] addr_3799_6;

Selector_2 s3799_6(wires_949_5[3], addr_949_5, wires_3799_6,addr_3799_6);

wire[3:0] wires_3800_6;

wire[31:0] addr_3800_6;

Selector_2 s3800_6(wires_950_5[0], addr_950_5, wires_3800_6,addr_3800_6);

wire[3:0] wires_3801_6;

wire[31:0] addr_3801_6;

Selector_2 s3801_6(wires_950_5[1], addr_950_5, wires_3801_6,addr_3801_6);

wire[3:0] wires_3802_6;

wire[31:0] addr_3802_6;

Selector_2 s3802_6(wires_950_5[2], addr_950_5, wires_3802_6,addr_3802_6);

wire[3:0] wires_3803_6;

wire[31:0] addr_3803_6;

Selector_2 s3803_6(wires_950_5[3], addr_950_5, wires_3803_6,addr_3803_6);

wire[3:0] wires_3804_6;

wire[31:0] addr_3804_6;

Selector_2 s3804_6(wires_951_5[0], addr_951_5, wires_3804_6,addr_3804_6);

wire[3:0] wires_3805_6;

wire[31:0] addr_3805_6;

Selector_2 s3805_6(wires_951_5[1], addr_951_5, wires_3805_6,addr_3805_6);

wire[3:0] wires_3806_6;

wire[31:0] addr_3806_6;

Selector_2 s3806_6(wires_951_5[2], addr_951_5, wires_3806_6,addr_3806_6);

wire[3:0] wires_3807_6;

wire[31:0] addr_3807_6;

Selector_2 s3807_6(wires_951_5[3], addr_951_5, wires_3807_6,addr_3807_6);

wire[3:0] wires_3808_6;

wire[31:0] addr_3808_6;

Selector_2 s3808_6(wires_952_5[0], addr_952_5, wires_3808_6,addr_3808_6);

wire[3:0] wires_3809_6;

wire[31:0] addr_3809_6;

Selector_2 s3809_6(wires_952_5[1], addr_952_5, wires_3809_6,addr_3809_6);

wire[3:0] wires_3810_6;

wire[31:0] addr_3810_6;

Selector_2 s3810_6(wires_952_5[2], addr_952_5, wires_3810_6,addr_3810_6);

wire[3:0] wires_3811_6;

wire[31:0] addr_3811_6;

Selector_2 s3811_6(wires_952_5[3], addr_952_5, wires_3811_6,addr_3811_6);

wire[3:0] wires_3812_6;

wire[31:0] addr_3812_6;

Selector_2 s3812_6(wires_953_5[0], addr_953_5, wires_3812_6,addr_3812_6);

wire[3:0] wires_3813_6;

wire[31:0] addr_3813_6;

Selector_2 s3813_6(wires_953_5[1], addr_953_5, wires_3813_6,addr_3813_6);

wire[3:0] wires_3814_6;

wire[31:0] addr_3814_6;

Selector_2 s3814_6(wires_953_5[2], addr_953_5, wires_3814_6,addr_3814_6);

wire[3:0] wires_3815_6;

wire[31:0] addr_3815_6;

Selector_2 s3815_6(wires_953_5[3], addr_953_5, wires_3815_6,addr_3815_6);

wire[3:0] wires_3816_6;

wire[31:0] addr_3816_6;

Selector_2 s3816_6(wires_954_5[0], addr_954_5, wires_3816_6,addr_3816_6);

wire[3:0] wires_3817_6;

wire[31:0] addr_3817_6;

Selector_2 s3817_6(wires_954_5[1], addr_954_5, wires_3817_6,addr_3817_6);

wire[3:0] wires_3818_6;

wire[31:0] addr_3818_6;

Selector_2 s3818_6(wires_954_5[2], addr_954_5, wires_3818_6,addr_3818_6);

wire[3:0] wires_3819_6;

wire[31:0] addr_3819_6;

Selector_2 s3819_6(wires_954_5[3], addr_954_5, wires_3819_6,addr_3819_6);

wire[3:0] wires_3820_6;

wire[31:0] addr_3820_6;

Selector_2 s3820_6(wires_955_5[0], addr_955_5, wires_3820_6,addr_3820_6);

wire[3:0] wires_3821_6;

wire[31:0] addr_3821_6;

Selector_2 s3821_6(wires_955_5[1], addr_955_5, wires_3821_6,addr_3821_6);

wire[3:0] wires_3822_6;

wire[31:0] addr_3822_6;

Selector_2 s3822_6(wires_955_5[2], addr_955_5, wires_3822_6,addr_3822_6);

wire[3:0] wires_3823_6;

wire[31:0] addr_3823_6;

Selector_2 s3823_6(wires_955_5[3], addr_955_5, wires_3823_6,addr_3823_6);

wire[3:0] wires_3824_6;

wire[31:0] addr_3824_6;

Selector_2 s3824_6(wires_956_5[0], addr_956_5, wires_3824_6,addr_3824_6);

wire[3:0] wires_3825_6;

wire[31:0] addr_3825_6;

Selector_2 s3825_6(wires_956_5[1], addr_956_5, wires_3825_6,addr_3825_6);

wire[3:0] wires_3826_6;

wire[31:0] addr_3826_6;

Selector_2 s3826_6(wires_956_5[2], addr_956_5, wires_3826_6,addr_3826_6);

wire[3:0] wires_3827_6;

wire[31:0] addr_3827_6;

Selector_2 s3827_6(wires_956_5[3], addr_956_5, wires_3827_6,addr_3827_6);

wire[3:0] wires_3828_6;

wire[31:0] addr_3828_6;

Selector_2 s3828_6(wires_957_5[0], addr_957_5, wires_3828_6,addr_3828_6);

wire[3:0] wires_3829_6;

wire[31:0] addr_3829_6;

Selector_2 s3829_6(wires_957_5[1], addr_957_5, wires_3829_6,addr_3829_6);

wire[3:0] wires_3830_6;

wire[31:0] addr_3830_6;

Selector_2 s3830_6(wires_957_5[2], addr_957_5, wires_3830_6,addr_3830_6);

wire[3:0] wires_3831_6;

wire[31:0] addr_3831_6;

Selector_2 s3831_6(wires_957_5[3], addr_957_5, wires_3831_6,addr_3831_6);

wire[3:0] wires_3832_6;

wire[31:0] addr_3832_6;

Selector_2 s3832_6(wires_958_5[0], addr_958_5, wires_3832_6,addr_3832_6);

wire[3:0] wires_3833_6;

wire[31:0] addr_3833_6;

Selector_2 s3833_6(wires_958_5[1], addr_958_5, wires_3833_6,addr_3833_6);

wire[3:0] wires_3834_6;

wire[31:0] addr_3834_6;

Selector_2 s3834_6(wires_958_5[2], addr_958_5, wires_3834_6,addr_3834_6);

wire[3:0] wires_3835_6;

wire[31:0] addr_3835_6;

Selector_2 s3835_6(wires_958_5[3], addr_958_5, wires_3835_6,addr_3835_6);

wire[3:0] wires_3836_6;

wire[31:0] addr_3836_6;

Selector_2 s3836_6(wires_959_5[0], addr_959_5, wires_3836_6,addr_3836_6);

wire[3:0] wires_3837_6;

wire[31:0] addr_3837_6;

Selector_2 s3837_6(wires_959_5[1], addr_959_5, wires_3837_6,addr_3837_6);

wire[3:0] wires_3838_6;

wire[31:0] addr_3838_6;

Selector_2 s3838_6(wires_959_5[2], addr_959_5, wires_3838_6,addr_3838_6);

wire[3:0] wires_3839_6;

wire[31:0] addr_3839_6;

Selector_2 s3839_6(wires_959_5[3], addr_959_5, wires_3839_6,addr_3839_6);

wire[3:0] wires_3840_6;

wire[31:0] addr_3840_6;

Selector_2 s3840_6(wires_960_5[0], addr_960_5, wires_3840_6,addr_3840_6);

wire[3:0] wires_3841_6;

wire[31:0] addr_3841_6;

Selector_2 s3841_6(wires_960_5[1], addr_960_5, wires_3841_6,addr_3841_6);

wire[3:0] wires_3842_6;

wire[31:0] addr_3842_6;

Selector_2 s3842_6(wires_960_5[2], addr_960_5, wires_3842_6,addr_3842_6);

wire[3:0] wires_3843_6;

wire[31:0] addr_3843_6;

Selector_2 s3843_6(wires_960_5[3], addr_960_5, wires_3843_6,addr_3843_6);

wire[3:0] wires_3844_6;

wire[31:0] addr_3844_6;

Selector_2 s3844_6(wires_961_5[0], addr_961_5, wires_3844_6,addr_3844_6);

wire[3:0] wires_3845_6;

wire[31:0] addr_3845_6;

Selector_2 s3845_6(wires_961_5[1], addr_961_5, wires_3845_6,addr_3845_6);

wire[3:0] wires_3846_6;

wire[31:0] addr_3846_6;

Selector_2 s3846_6(wires_961_5[2], addr_961_5, wires_3846_6,addr_3846_6);

wire[3:0] wires_3847_6;

wire[31:0] addr_3847_6;

Selector_2 s3847_6(wires_961_5[3], addr_961_5, wires_3847_6,addr_3847_6);

wire[3:0] wires_3848_6;

wire[31:0] addr_3848_6;

Selector_2 s3848_6(wires_962_5[0], addr_962_5, wires_3848_6,addr_3848_6);

wire[3:0] wires_3849_6;

wire[31:0] addr_3849_6;

Selector_2 s3849_6(wires_962_5[1], addr_962_5, wires_3849_6,addr_3849_6);

wire[3:0] wires_3850_6;

wire[31:0] addr_3850_6;

Selector_2 s3850_6(wires_962_5[2], addr_962_5, wires_3850_6,addr_3850_6);

wire[3:0] wires_3851_6;

wire[31:0] addr_3851_6;

Selector_2 s3851_6(wires_962_5[3], addr_962_5, wires_3851_6,addr_3851_6);

wire[3:0] wires_3852_6;

wire[31:0] addr_3852_6;

Selector_2 s3852_6(wires_963_5[0], addr_963_5, wires_3852_6,addr_3852_6);

wire[3:0] wires_3853_6;

wire[31:0] addr_3853_6;

Selector_2 s3853_6(wires_963_5[1], addr_963_5, wires_3853_6,addr_3853_6);

wire[3:0] wires_3854_6;

wire[31:0] addr_3854_6;

Selector_2 s3854_6(wires_963_5[2], addr_963_5, wires_3854_6,addr_3854_6);

wire[3:0] wires_3855_6;

wire[31:0] addr_3855_6;

Selector_2 s3855_6(wires_963_5[3], addr_963_5, wires_3855_6,addr_3855_6);

wire[3:0] wires_3856_6;

wire[31:0] addr_3856_6;

Selector_2 s3856_6(wires_964_5[0], addr_964_5, wires_3856_6,addr_3856_6);

wire[3:0] wires_3857_6;

wire[31:0] addr_3857_6;

Selector_2 s3857_6(wires_964_5[1], addr_964_5, wires_3857_6,addr_3857_6);

wire[3:0] wires_3858_6;

wire[31:0] addr_3858_6;

Selector_2 s3858_6(wires_964_5[2], addr_964_5, wires_3858_6,addr_3858_6);

wire[3:0] wires_3859_6;

wire[31:0] addr_3859_6;

Selector_2 s3859_6(wires_964_5[3], addr_964_5, wires_3859_6,addr_3859_6);

wire[3:0] wires_3860_6;

wire[31:0] addr_3860_6;

Selector_2 s3860_6(wires_965_5[0], addr_965_5, wires_3860_6,addr_3860_6);

wire[3:0] wires_3861_6;

wire[31:0] addr_3861_6;

Selector_2 s3861_6(wires_965_5[1], addr_965_5, wires_3861_6,addr_3861_6);

wire[3:0] wires_3862_6;

wire[31:0] addr_3862_6;

Selector_2 s3862_6(wires_965_5[2], addr_965_5, wires_3862_6,addr_3862_6);

wire[3:0] wires_3863_6;

wire[31:0] addr_3863_6;

Selector_2 s3863_6(wires_965_5[3], addr_965_5, wires_3863_6,addr_3863_6);

wire[3:0] wires_3864_6;

wire[31:0] addr_3864_6;

Selector_2 s3864_6(wires_966_5[0], addr_966_5, wires_3864_6,addr_3864_6);

wire[3:0] wires_3865_6;

wire[31:0] addr_3865_6;

Selector_2 s3865_6(wires_966_5[1], addr_966_5, wires_3865_6,addr_3865_6);

wire[3:0] wires_3866_6;

wire[31:0] addr_3866_6;

Selector_2 s3866_6(wires_966_5[2], addr_966_5, wires_3866_6,addr_3866_6);

wire[3:0] wires_3867_6;

wire[31:0] addr_3867_6;

Selector_2 s3867_6(wires_966_5[3], addr_966_5, wires_3867_6,addr_3867_6);

wire[3:0] wires_3868_6;

wire[31:0] addr_3868_6;

Selector_2 s3868_6(wires_967_5[0], addr_967_5, wires_3868_6,addr_3868_6);

wire[3:0] wires_3869_6;

wire[31:0] addr_3869_6;

Selector_2 s3869_6(wires_967_5[1], addr_967_5, wires_3869_6,addr_3869_6);

wire[3:0] wires_3870_6;

wire[31:0] addr_3870_6;

Selector_2 s3870_6(wires_967_5[2], addr_967_5, wires_3870_6,addr_3870_6);

wire[3:0] wires_3871_6;

wire[31:0] addr_3871_6;

Selector_2 s3871_6(wires_967_5[3], addr_967_5, wires_3871_6,addr_3871_6);

wire[3:0] wires_3872_6;

wire[31:0] addr_3872_6;

Selector_2 s3872_6(wires_968_5[0], addr_968_5, wires_3872_6,addr_3872_6);

wire[3:0] wires_3873_6;

wire[31:0] addr_3873_6;

Selector_2 s3873_6(wires_968_5[1], addr_968_5, wires_3873_6,addr_3873_6);

wire[3:0] wires_3874_6;

wire[31:0] addr_3874_6;

Selector_2 s3874_6(wires_968_5[2], addr_968_5, wires_3874_6,addr_3874_6);

wire[3:0] wires_3875_6;

wire[31:0] addr_3875_6;

Selector_2 s3875_6(wires_968_5[3], addr_968_5, wires_3875_6,addr_3875_6);

wire[3:0] wires_3876_6;

wire[31:0] addr_3876_6;

Selector_2 s3876_6(wires_969_5[0], addr_969_5, wires_3876_6,addr_3876_6);

wire[3:0] wires_3877_6;

wire[31:0] addr_3877_6;

Selector_2 s3877_6(wires_969_5[1], addr_969_5, wires_3877_6,addr_3877_6);

wire[3:0] wires_3878_6;

wire[31:0] addr_3878_6;

Selector_2 s3878_6(wires_969_5[2], addr_969_5, wires_3878_6,addr_3878_6);

wire[3:0] wires_3879_6;

wire[31:0] addr_3879_6;

Selector_2 s3879_6(wires_969_5[3], addr_969_5, wires_3879_6,addr_3879_6);

wire[3:0] wires_3880_6;

wire[31:0] addr_3880_6;

Selector_2 s3880_6(wires_970_5[0], addr_970_5, wires_3880_6,addr_3880_6);

wire[3:0] wires_3881_6;

wire[31:0] addr_3881_6;

Selector_2 s3881_6(wires_970_5[1], addr_970_5, wires_3881_6,addr_3881_6);

wire[3:0] wires_3882_6;

wire[31:0] addr_3882_6;

Selector_2 s3882_6(wires_970_5[2], addr_970_5, wires_3882_6,addr_3882_6);

wire[3:0] wires_3883_6;

wire[31:0] addr_3883_6;

Selector_2 s3883_6(wires_970_5[3], addr_970_5, wires_3883_6,addr_3883_6);

wire[3:0] wires_3884_6;

wire[31:0] addr_3884_6;

Selector_2 s3884_6(wires_971_5[0], addr_971_5, wires_3884_6,addr_3884_6);

wire[3:0] wires_3885_6;

wire[31:0] addr_3885_6;

Selector_2 s3885_6(wires_971_5[1], addr_971_5, wires_3885_6,addr_3885_6);

wire[3:0] wires_3886_6;

wire[31:0] addr_3886_6;

Selector_2 s3886_6(wires_971_5[2], addr_971_5, wires_3886_6,addr_3886_6);

wire[3:0] wires_3887_6;

wire[31:0] addr_3887_6;

Selector_2 s3887_6(wires_971_5[3], addr_971_5, wires_3887_6,addr_3887_6);

wire[3:0] wires_3888_6;

wire[31:0] addr_3888_6;

Selector_2 s3888_6(wires_972_5[0], addr_972_5, wires_3888_6,addr_3888_6);

wire[3:0] wires_3889_6;

wire[31:0] addr_3889_6;

Selector_2 s3889_6(wires_972_5[1], addr_972_5, wires_3889_6,addr_3889_6);

wire[3:0] wires_3890_6;

wire[31:0] addr_3890_6;

Selector_2 s3890_6(wires_972_5[2], addr_972_5, wires_3890_6,addr_3890_6);

wire[3:0] wires_3891_6;

wire[31:0] addr_3891_6;

Selector_2 s3891_6(wires_972_5[3], addr_972_5, wires_3891_6,addr_3891_6);

wire[3:0] wires_3892_6;

wire[31:0] addr_3892_6;

Selector_2 s3892_6(wires_973_5[0], addr_973_5, wires_3892_6,addr_3892_6);

wire[3:0] wires_3893_6;

wire[31:0] addr_3893_6;

Selector_2 s3893_6(wires_973_5[1], addr_973_5, wires_3893_6,addr_3893_6);

wire[3:0] wires_3894_6;

wire[31:0] addr_3894_6;

Selector_2 s3894_6(wires_973_5[2], addr_973_5, wires_3894_6,addr_3894_6);

wire[3:0] wires_3895_6;

wire[31:0] addr_3895_6;

Selector_2 s3895_6(wires_973_5[3], addr_973_5, wires_3895_6,addr_3895_6);

wire[3:0] wires_3896_6;

wire[31:0] addr_3896_6;

Selector_2 s3896_6(wires_974_5[0], addr_974_5, wires_3896_6,addr_3896_6);

wire[3:0] wires_3897_6;

wire[31:0] addr_3897_6;

Selector_2 s3897_6(wires_974_5[1], addr_974_5, wires_3897_6,addr_3897_6);

wire[3:0] wires_3898_6;

wire[31:0] addr_3898_6;

Selector_2 s3898_6(wires_974_5[2], addr_974_5, wires_3898_6,addr_3898_6);

wire[3:0] wires_3899_6;

wire[31:0] addr_3899_6;

Selector_2 s3899_6(wires_974_5[3], addr_974_5, wires_3899_6,addr_3899_6);

wire[3:0] wires_3900_6;

wire[31:0] addr_3900_6;

Selector_2 s3900_6(wires_975_5[0], addr_975_5, wires_3900_6,addr_3900_6);

wire[3:0] wires_3901_6;

wire[31:0] addr_3901_6;

Selector_2 s3901_6(wires_975_5[1], addr_975_5, wires_3901_6,addr_3901_6);

wire[3:0] wires_3902_6;

wire[31:0] addr_3902_6;

Selector_2 s3902_6(wires_975_5[2], addr_975_5, wires_3902_6,addr_3902_6);

wire[3:0] wires_3903_6;

wire[31:0] addr_3903_6;

Selector_2 s3903_6(wires_975_5[3], addr_975_5, wires_3903_6,addr_3903_6);

wire[3:0] wires_3904_6;

wire[31:0] addr_3904_6;

Selector_2 s3904_6(wires_976_5[0], addr_976_5, wires_3904_6,addr_3904_6);

wire[3:0] wires_3905_6;

wire[31:0] addr_3905_6;

Selector_2 s3905_6(wires_976_5[1], addr_976_5, wires_3905_6,addr_3905_6);

wire[3:0] wires_3906_6;

wire[31:0] addr_3906_6;

Selector_2 s3906_6(wires_976_5[2], addr_976_5, wires_3906_6,addr_3906_6);

wire[3:0] wires_3907_6;

wire[31:0] addr_3907_6;

Selector_2 s3907_6(wires_976_5[3], addr_976_5, wires_3907_6,addr_3907_6);

wire[3:0] wires_3908_6;

wire[31:0] addr_3908_6;

Selector_2 s3908_6(wires_977_5[0], addr_977_5, wires_3908_6,addr_3908_6);

wire[3:0] wires_3909_6;

wire[31:0] addr_3909_6;

Selector_2 s3909_6(wires_977_5[1], addr_977_5, wires_3909_6,addr_3909_6);

wire[3:0] wires_3910_6;

wire[31:0] addr_3910_6;

Selector_2 s3910_6(wires_977_5[2], addr_977_5, wires_3910_6,addr_3910_6);

wire[3:0] wires_3911_6;

wire[31:0] addr_3911_6;

Selector_2 s3911_6(wires_977_5[3], addr_977_5, wires_3911_6,addr_3911_6);

wire[3:0] wires_3912_6;

wire[31:0] addr_3912_6;

Selector_2 s3912_6(wires_978_5[0], addr_978_5, wires_3912_6,addr_3912_6);

wire[3:0] wires_3913_6;

wire[31:0] addr_3913_6;

Selector_2 s3913_6(wires_978_5[1], addr_978_5, wires_3913_6,addr_3913_6);

wire[3:0] wires_3914_6;

wire[31:0] addr_3914_6;

Selector_2 s3914_6(wires_978_5[2], addr_978_5, wires_3914_6,addr_3914_6);

wire[3:0] wires_3915_6;

wire[31:0] addr_3915_6;

Selector_2 s3915_6(wires_978_5[3], addr_978_5, wires_3915_6,addr_3915_6);

wire[3:0] wires_3916_6;

wire[31:0] addr_3916_6;

Selector_2 s3916_6(wires_979_5[0], addr_979_5, wires_3916_6,addr_3916_6);

wire[3:0] wires_3917_6;

wire[31:0] addr_3917_6;

Selector_2 s3917_6(wires_979_5[1], addr_979_5, wires_3917_6,addr_3917_6);

wire[3:0] wires_3918_6;

wire[31:0] addr_3918_6;

Selector_2 s3918_6(wires_979_5[2], addr_979_5, wires_3918_6,addr_3918_6);

wire[3:0] wires_3919_6;

wire[31:0] addr_3919_6;

Selector_2 s3919_6(wires_979_5[3], addr_979_5, wires_3919_6,addr_3919_6);

wire[3:0] wires_3920_6;

wire[31:0] addr_3920_6;

Selector_2 s3920_6(wires_980_5[0], addr_980_5, wires_3920_6,addr_3920_6);

wire[3:0] wires_3921_6;

wire[31:0] addr_3921_6;

Selector_2 s3921_6(wires_980_5[1], addr_980_5, wires_3921_6,addr_3921_6);

wire[3:0] wires_3922_6;

wire[31:0] addr_3922_6;

Selector_2 s3922_6(wires_980_5[2], addr_980_5, wires_3922_6,addr_3922_6);

wire[3:0] wires_3923_6;

wire[31:0] addr_3923_6;

Selector_2 s3923_6(wires_980_5[3], addr_980_5, wires_3923_6,addr_3923_6);

wire[3:0] wires_3924_6;

wire[31:0] addr_3924_6;

Selector_2 s3924_6(wires_981_5[0], addr_981_5, wires_3924_6,addr_3924_6);

wire[3:0] wires_3925_6;

wire[31:0] addr_3925_6;

Selector_2 s3925_6(wires_981_5[1], addr_981_5, wires_3925_6,addr_3925_6);

wire[3:0] wires_3926_6;

wire[31:0] addr_3926_6;

Selector_2 s3926_6(wires_981_5[2], addr_981_5, wires_3926_6,addr_3926_6);

wire[3:0] wires_3927_6;

wire[31:0] addr_3927_6;

Selector_2 s3927_6(wires_981_5[3], addr_981_5, wires_3927_6,addr_3927_6);

wire[3:0] wires_3928_6;

wire[31:0] addr_3928_6;

Selector_2 s3928_6(wires_982_5[0], addr_982_5, wires_3928_6,addr_3928_6);

wire[3:0] wires_3929_6;

wire[31:0] addr_3929_6;

Selector_2 s3929_6(wires_982_5[1], addr_982_5, wires_3929_6,addr_3929_6);

wire[3:0] wires_3930_6;

wire[31:0] addr_3930_6;

Selector_2 s3930_6(wires_982_5[2], addr_982_5, wires_3930_6,addr_3930_6);

wire[3:0] wires_3931_6;

wire[31:0] addr_3931_6;

Selector_2 s3931_6(wires_982_5[3], addr_982_5, wires_3931_6,addr_3931_6);

wire[3:0] wires_3932_6;

wire[31:0] addr_3932_6;

Selector_2 s3932_6(wires_983_5[0], addr_983_5, wires_3932_6,addr_3932_6);

wire[3:0] wires_3933_6;

wire[31:0] addr_3933_6;

Selector_2 s3933_6(wires_983_5[1], addr_983_5, wires_3933_6,addr_3933_6);

wire[3:0] wires_3934_6;

wire[31:0] addr_3934_6;

Selector_2 s3934_6(wires_983_5[2], addr_983_5, wires_3934_6,addr_3934_6);

wire[3:0] wires_3935_6;

wire[31:0] addr_3935_6;

Selector_2 s3935_6(wires_983_5[3], addr_983_5, wires_3935_6,addr_3935_6);

wire[3:0] wires_3936_6;

wire[31:0] addr_3936_6;

Selector_2 s3936_6(wires_984_5[0], addr_984_5, wires_3936_6,addr_3936_6);

wire[3:0] wires_3937_6;

wire[31:0] addr_3937_6;

Selector_2 s3937_6(wires_984_5[1], addr_984_5, wires_3937_6,addr_3937_6);

wire[3:0] wires_3938_6;

wire[31:0] addr_3938_6;

Selector_2 s3938_6(wires_984_5[2], addr_984_5, wires_3938_6,addr_3938_6);

wire[3:0] wires_3939_6;

wire[31:0] addr_3939_6;

Selector_2 s3939_6(wires_984_5[3], addr_984_5, wires_3939_6,addr_3939_6);

wire[3:0] wires_3940_6;

wire[31:0] addr_3940_6;

Selector_2 s3940_6(wires_985_5[0], addr_985_5, wires_3940_6,addr_3940_6);

wire[3:0] wires_3941_6;

wire[31:0] addr_3941_6;

Selector_2 s3941_6(wires_985_5[1], addr_985_5, wires_3941_6,addr_3941_6);

wire[3:0] wires_3942_6;

wire[31:0] addr_3942_6;

Selector_2 s3942_6(wires_985_5[2], addr_985_5, wires_3942_6,addr_3942_6);

wire[3:0] wires_3943_6;

wire[31:0] addr_3943_6;

Selector_2 s3943_6(wires_985_5[3], addr_985_5, wires_3943_6,addr_3943_6);

wire[3:0] wires_3944_6;

wire[31:0] addr_3944_6;

Selector_2 s3944_6(wires_986_5[0], addr_986_5, wires_3944_6,addr_3944_6);

wire[3:0] wires_3945_6;

wire[31:0] addr_3945_6;

Selector_2 s3945_6(wires_986_5[1], addr_986_5, wires_3945_6,addr_3945_6);

wire[3:0] wires_3946_6;

wire[31:0] addr_3946_6;

Selector_2 s3946_6(wires_986_5[2], addr_986_5, wires_3946_6,addr_3946_6);

wire[3:0] wires_3947_6;

wire[31:0] addr_3947_6;

Selector_2 s3947_6(wires_986_5[3], addr_986_5, wires_3947_6,addr_3947_6);

wire[3:0] wires_3948_6;

wire[31:0] addr_3948_6;

Selector_2 s3948_6(wires_987_5[0], addr_987_5, wires_3948_6,addr_3948_6);

wire[3:0] wires_3949_6;

wire[31:0] addr_3949_6;

Selector_2 s3949_6(wires_987_5[1], addr_987_5, wires_3949_6,addr_3949_6);

wire[3:0] wires_3950_6;

wire[31:0] addr_3950_6;

Selector_2 s3950_6(wires_987_5[2], addr_987_5, wires_3950_6,addr_3950_6);

wire[3:0] wires_3951_6;

wire[31:0] addr_3951_6;

Selector_2 s3951_6(wires_987_5[3], addr_987_5, wires_3951_6,addr_3951_6);

wire[3:0] wires_3952_6;

wire[31:0] addr_3952_6;

Selector_2 s3952_6(wires_988_5[0], addr_988_5, wires_3952_6,addr_3952_6);

wire[3:0] wires_3953_6;

wire[31:0] addr_3953_6;

Selector_2 s3953_6(wires_988_5[1], addr_988_5, wires_3953_6,addr_3953_6);

wire[3:0] wires_3954_6;

wire[31:0] addr_3954_6;

Selector_2 s3954_6(wires_988_5[2], addr_988_5, wires_3954_6,addr_3954_6);

wire[3:0] wires_3955_6;

wire[31:0] addr_3955_6;

Selector_2 s3955_6(wires_988_5[3], addr_988_5, wires_3955_6,addr_3955_6);

wire[3:0] wires_3956_6;

wire[31:0] addr_3956_6;

Selector_2 s3956_6(wires_989_5[0], addr_989_5, wires_3956_6,addr_3956_6);

wire[3:0] wires_3957_6;

wire[31:0] addr_3957_6;

Selector_2 s3957_6(wires_989_5[1], addr_989_5, wires_3957_6,addr_3957_6);

wire[3:0] wires_3958_6;

wire[31:0] addr_3958_6;

Selector_2 s3958_6(wires_989_5[2], addr_989_5, wires_3958_6,addr_3958_6);

wire[3:0] wires_3959_6;

wire[31:0] addr_3959_6;

Selector_2 s3959_6(wires_989_5[3], addr_989_5, wires_3959_6,addr_3959_6);

wire[3:0] wires_3960_6;

wire[31:0] addr_3960_6;

Selector_2 s3960_6(wires_990_5[0], addr_990_5, wires_3960_6,addr_3960_6);

wire[3:0] wires_3961_6;

wire[31:0] addr_3961_6;

Selector_2 s3961_6(wires_990_5[1], addr_990_5, wires_3961_6,addr_3961_6);

wire[3:0] wires_3962_6;

wire[31:0] addr_3962_6;

Selector_2 s3962_6(wires_990_5[2], addr_990_5, wires_3962_6,addr_3962_6);

wire[3:0] wires_3963_6;

wire[31:0] addr_3963_6;

Selector_2 s3963_6(wires_990_5[3], addr_990_5, wires_3963_6,addr_3963_6);

wire[3:0] wires_3964_6;

wire[31:0] addr_3964_6;

Selector_2 s3964_6(wires_991_5[0], addr_991_5, wires_3964_6,addr_3964_6);

wire[3:0] wires_3965_6;

wire[31:0] addr_3965_6;

Selector_2 s3965_6(wires_991_5[1], addr_991_5, wires_3965_6,addr_3965_6);

wire[3:0] wires_3966_6;

wire[31:0] addr_3966_6;

Selector_2 s3966_6(wires_991_5[2], addr_991_5, wires_3966_6,addr_3966_6);

wire[3:0] wires_3967_6;

wire[31:0] addr_3967_6;

Selector_2 s3967_6(wires_991_5[3], addr_991_5, wires_3967_6,addr_3967_6);

wire[3:0] wires_3968_6;

wire[31:0] addr_3968_6;

Selector_2 s3968_6(wires_992_5[0], addr_992_5, wires_3968_6,addr_3968_6);

wire[3:0] wires_3969_6;

wire[31:0] addr_3969_6;

Selector_2 s3969_6(wires_992_5[1], addr_992_5, wires_3969_6,addr_3969_6);

wire[3:0] wires_3970_6;

wire[31:0] addr_3970_6;

Selector_2 s3970_6(wires_992_5[2], addr_992_5, wires_3970_6,addr_3970_6);

wire[3:0] wires_3971_6;

wire[31:0] addr_3971_6;

Selector_2 s3971_6(wires_992_5[3], addr_992_5, wires_3971_6,addr_3971_6);

wire[3:0] wires_3972_6;

wire[31:0] addr_3972_6;

Selector_2 s3972_6(wires_993_5[0], addr_993_5, wires_3972_6,addr_3972_6);

wire[3:0] wires_3973_6;

wire[31:0] addr_3973_6;

Selector_2 s3973_6(wires_993_5[1], addr_993_5, wires_3973_6,addr_3973_6);

wire[3:0] wires_3974_6;

wire[31:0] addr_3974_6;

Selector_2 s3974_6(wires_993_5[2], addr_993_5, wires_3974_6,addr_3974_6);

wire[3:0] wires_3975_6;

wire[31:0] addr_3975_6;

Selector_2 s3975_6(wires_993_5[3], addr_993_5, wires_3975_6,addr_3975_6);

wire[3:0] wires_3976_6;

wire[31:0] addr_3976_6;

Selector_2 s3976_6(wires_994_5[0], addr_994_5, wires_3976_6,addr_3976_6);

wire[3:0] wires_3977_6;

wire[31:0] addr_3977_6;

Selector_2 s3977_6(wires_994_5[1], addr_994_5, wires_3977_6,addr_3977_6);

wire[3:0] wires_3978_6;

wire[31:0] addr_3978_6;

Selector_2 s3978_6(wires_994_5[2], addr_994_5, wires_3978_6,addr_3978_6);

wire[3:0] wires_3979_6;

wire[31:0] addr_3979_6;

Selector_2 s3979_6(wires_994_5[3], addr_994_5, wires_3979_6,addr_3979_6);

wire[3:0] wires_3980_6;

wire[31:0] addr_3980_6;

Selector_2 s3980_6(wires_995_5[0], addr_995_5, wires_3980_6,addr_3980_6);

wire[3:0] wires_3981_6;

wire[31:0] addr_3981_6;

Selector_2 s3981_6(wires_995_5[1], addr_995_5, wires_3981_6,addr_3981_6);

wire[3:0] wires_3982_6;

wire[31:0] addr_3982_6;

Selector_2 s3982_6(wires_995_5[2], addr_995_5, wires_3982_6,addr_3982_6);

wire[3:0] wires_3983_6;

wire[31:0] addr_3983_6;

Selector_2 s3983_6(wires_995_5[3], addr_995_5, wires_3983_6,addr_3983_6);

wire[3:0] wires_3984_6;

wire[31:0] addr_3984_6;

Selector_2 s3984_6(wires_996_5[0], addr_996_5, wires_3984_6,addr_3984_6);

wire[3:0] wires_3985_6;

wire[31:0] addr_3985_6;

Selector_2 s3985_6(wires_996_5[1], addr_996_5, wires_3985_6,addr_3985_6);

wire[3:0] wires_3986_6;

wire[31:0] addr_3986_6;

Selector_2 s3986_6(wires_996_5[2], addr_996_5, wires_3986_6,addr_3986_6);

wire[3:0] wires_3987_6;

wire[31:0] addr_3987_6;

Selector_2 s3987_6(wires_996_5[3], addr_996_5, wires_3987_6,addr_3987_6);

wire[3:0] wires_3988_6;

wire[31:0] addr_3988_6;

Selector_2 s3988_6(wires_997_5[0], addr_997_5, wires_3988_6,addr_3988_6);

wire[3:0] wires_3989_6;

wire[31:0] addr_3989_6;

Selector_2 s3989_6(wires_997_5[1], addr_997_5, wires_3989_6,addr_3989_6);

wire[3:0] wires_3990_6;

wire[31:0] addr_3990_6;

Selector_2 s3990_6(wires_997_5[2], addr_997_5, wires_3990_6,addr_3990_6);

wire[3:0] wires_3991_6;

wire[31:0] addr_3991_6;

Selector_2 s3991_6(wires_997_5[3], addr_997_5, wires_3991_6,addr_3991_6);

wire[3:0] wires_3992_6;

wire[31:0] addr_3992_6;

Selector_2 s3992_6(wires_998_5[0], addr_998_5, wires_3992_6,addr_3992_6);

wire[3:0] wires_3993_6;

wire[31:0] addr_3993_6;

Selector_2 s3993_6(wires_998_5[1], addr_998_5, wires_3993_6,addr_3993_6);

wire[3:0] wires_3994_6;

wire[31:0] addr_3994_6;

Selector_2 s3994_6(wires_998_5[2], addr_998_5, wires_3994_6,addr_3994_6);

wire[3:0] wires_3995_6;

wire[31:0] addr_3995_6;

Selector_2 s3995_6(wires_998_5[3], addr_998_5, wires_3995_6,addr_3995_6);

wire[3:0] wires_3996_6;

wire[31:0] addr_3996_6;

Selector_2 s3996_6(wires_999_5[0], addr_999_5, wires_3996_6,addr_3996_6);

wire[3:0] wires_3997_6;

wire[31:0] addr_3997_6;

Selector_2 s3997_6(wires_999_5[1], addr_999_5, wires_3997_6,addr_3997_6);

wire[3:0] wires_3998_6;

wire[31:0] addr_3998_6;

Selector_2 s3998_6(wires_999_5[2], addr_999_5, wires_3998_6,addr_3998_6);

wire[3:0] wires_3999_6;

wire[31:0] addr_3999_6;

Selector_2 s3999_6(wires_999_5[3], addr_999_5, wires_3999_6,addr_3999_6);

wire[3:0] wires_4000_6;

wire[31:0] addr_4000_6;

Selector_2 s4000_6(wires_1000_5[0], addr_1000_5, wires_4000_6,addr_4000_6);

wire[3:0] wires_4001_6;

wire[31:0] addr_4001_6;

Selector_2 s4001_6(wires_1000_5[1], addr_1000_5, wires_4001_6,addr_4001_6);

wire[3:0] wires_4002_6;

wire[31:0] addr_4002_6;

Selector_2 s4002_6(wires_1000_5[2], addr_1000_5, wires_4002_6,addr_4002_6);

wire[3:0] wires_4003_6;

wire[31:0] addr_4003_6;

Selector_2 s4003_6(wires_1000_5[3], addr_1000_5, wires_4003_6,addr_4003_6);

wire[3:0] wires_4004_6;

wire[31:0] addr_4004_6;

Selector_2 s4004_6(wires_1001_5[0], addr_1001_5, wires_4004_6,addr_4004_6);

wire[3:0] wires_4005_6;

wire[31:0] addr_4005_6;

Selector_2 s4005_6(wires_1001_5[1], addr_1001_5, wires_4005_6,addr_4005_6);

wire[3:0] wires_4006_6;

wire[31:0] addr_4006_6;

Selector_2 s4006_6(wires_1001_5[2], addr_1001_5, wires_4006_6,addr_4006_6);

wire[3:0] wires_4007_6;

wire[31:0] addr_4007_6;

Selector_2 s4007_6(wires_1001_5[3], addr_1001_5, wires_4007_6,addr_4007_6);

wire[3:0] wires_4008_6;

wire[31:0] addr_4008_6;

Selector_2 s4008_6(wires_1002_5[0], addr_1002_5, wires_4008_6,addr_4008_6);

wire[3:0] wires_4009_6;

wire[31:0] addr_4009_6;

Selector_2 s4009_6(wires_1002_5[1], addr_1002_5, wires_4009_6,addr_4009_6);

wire[3:0] wires_4010_6;

wire[31:0] addr_4010_6;

Selector_2 s4010_6(wires_1002_5[2], addr_1002_5, wires_4010_6,addr_4010_6);

wire[3:0] wires_4011_6;

wire[31:0] addr_4011_6;

Selector_2 s4011_6(wires_1002_5[3], addr_1002_5, wires_4011_6,addr_4011_6);

wire[3:0] wires_4012_6;

wire[31:0] addr_4012_6;

Selector_2 s4012_6(wires_1003_5[0], addr_1003_5, wires_4012_6,addr_4012_6);

wire[3:0] wires_4013_6;

wire[31:0] addr_4013_6;

Selector_2 s4013_6(wires_1003_5[1], addr_1003_5, wires_4013_6,addr_4013_6);

wire[3:0] wires_4014_6;

wire[31:0] addr_4014_6;

Selector_2 s4014_6(wires_1003_5[2], addr_1003_5, wires_4014_6,addr_4014_6);

wire[3:0] wires_4015_6;

wire[31:0] addr_4015_6;

Selector_2 s4015_6(wires_1003_5[3], addr_1003_5, wires_4015_6,addr_4015_6);

wire[3:0] wires_4016_6;

wire[31:0] addr_4016_6;

Selector_2 s4016_6(wires_1004_5[0], addr_1004_5, wires_4016_6,addr_4016_6);

wire[3:0] wires_4017_6;

wire[31:0] addr_4017_6;

Selector_2 s4017_6(wires_1004_5[1], addr_1004_5, wires_4017_6,addr_4017_6);

wire[3:0] wires_4018_6;

wire[31:0] addr_4018_6;

Selector_2 s4018_6(wires_1004_5[2], addr_1004_5, wires_4018_6,addr_4018_6);

wire[3:0] wires_4019_6;

wire[31:0] addr_4019_6;

Selector_2 s4019_6(wires_1004_5[3], addr_1004_5, wires_4019_6,addr_4019_6);

wire[3:0] wires_4020_6;

wire[31:0] addr_4020_6;

Selector_2 s4020_6(wires_1005_5[0], addr_1005_5, wires_4020_6,addr_4020_6);

wire[3:0] wires_4021_6;

wire[31:0] addr_4021_6;

Selector_2 s4021_6(wires_1005_5[1], addr_1005_5, wires_4021_6,addr_4021_6);

wire[3:0] wires_4022_6;

wire[31:0] addr_4022_6;

Selector_2 s4022_6(wires_1005_5[2], addr_1005_5, wires_4022_6,addr_4022_6);

wire[3:0] wires_4023_6;

wire[31:0] addr_4023_6;

Selector_2 s4023_6(wires_1005_5[3], addr_1005_5, wires_4023_6,addr_4023_6);

wire[3:0] wires_4024_6;

wire[31:0] addr_4024_6;

Selector_2 s4024_6(wires_1006_5[0], addr_1006_5, wires_4024_6,addr_4024_6);

wire[3:0] wires_4025_6;

wire[31:0] addr_4025_6;

Selector_2 s4025_6(wires_1006_5[1], addr_1006_5, wires_4025_6,addr_4025_6);

wire[3:0] wires_4026_6;

wire[31:0] addr_4026_6;

Selector_2 s4026_6(wires_1006_5[2], addr_1006_5, wires_4026_6,addr_4026_6);

wire[3:0] wires_4027_6;

wire[31:0] addr_4027_6;

Selector_2 s4027_6(wires_1006_5[3], addr_1006_5, wires_4027_6,addr_4027_6);

wire[3:0] wires_4028_6;

wire[31:0] addr_4028_6;

Selector_2 s4028_6(wires_1007_5[0], addr_1007_5, wires_4028_6,addr_4028_6);

wire[3:0] wires_4029_6;

wire[31:0] addr_4029_6;

Selector_2 s4029_6(wires_1007_5[1], addr_1007_5, wires_4029_6,addr_4029_6);

wire[3:0] wires_4030_6;

wire[31:0] addr_4030_6;

Selector_2 s4030_6(wires_1007_5[2], addr_1007_5, wires_4030_6,addr_4030_6);

wire[3:0] wires_4031_6;

wire[31:0] addr_4031_6;

Selector_2 s4031_6(wires_1007_5[3], addr_1007_5, wires_4031_6,addr_4031_6);

wire[3:0] wires_4032_6;

wire[31:0] addr_4032_6;

Selector_2 s4032_6(wires_1008_5[0], addr_1008_5, wires_4032_6,addr_4032_6);

wire[3:0] wires_4033_6;

wire[31:0] addr_4033_6;

Selector_2 s4033_6(wires_1008_5[1], addr_1008_5, wires_4033_6,addr_4033_6);

wire[3:0] wires_4034_6;

wire[31:0] addr_4034_6;

Selector_2 s4034_6(wires_1008_5[2], addr_1008_5, wires_4034_6,addr_4034_6);

wire[3:0] wires_4035_6;

wire[31:0] addr_4035_6;

Selector_2 s4035_6(wires_1008_5[3], addr_1008_5, wires_4035_6,addr_4035_6);

wire[3:0] wires_4036_6;

wire[31:0] addr_4036_6;

Selector_2 s4036_6(wires_1009_5[0], addr_1009_5, wires_4036_6,addr_4036_6);

wire[3:0] wires_4037_6;

wire[31:0] addr_4037_6;

Selector_2 s4037_6(wires_1009_5[1], addr_1009_5, wires_4037_6,addr_4037_6);

wire[3:0] wires_4038_6;

wire[31:0] addr_4038_6;

Selector_2 s4038_6(wires_1009_5[2], addr_1009_5, wires_4038_6,addr_4038_6);

wire[3:0] wires_4039_6;

wire[31:0] addr_4039_6;

Selector_2 s4039_6(wires_1009_5[3], addr_1009_5, wires_4039_6,addr_4039_6);

wire[3:0] wires_4040_6;

wire[31:0] addr_4040_6;

Selector_2 s4040_6(wires_1010_5[0], addr_1010_5, wires_4040_6,addr_4040_6);

wire[3:0] wires_4041_6;

wire[31:0] addr_4041_6;

Selector_2 s4041_6(wires_1010_5[1], addr_1010_5, wires_4041_6,addr_4041_6);

wire[3:0] wires_4042_6;

wire[31:0] addr_4042_6;

Selector_2 s4042_6(wires_1010_5[2], addr_1010_5, wires_4042_6,addr_4042_6);

wire[3:0] wires_4043_6;

wire[31:0] addr_4043_6;

Selector_2 s4043_6(wires_1010_5[3], addr_1010_5, wires_4043_6,addr_4043_6);

wire[3:0] wires_4044_6;

wire[31:0] addr_4044_6;

Selector_2 s4044_6(wires_1011_5[0], addr_1011_5, wires_4044_6,addr_4044_6);

wire[3:0] wires_4045_6;

wire[31:0] addr_4045_6;

Selector_2 s4045_6(wires_1011_5[1], addr_1011_5, wires_4045_6,addr_4045_6);

wire[3:0] wires_4046_6;

wire[31:0] addr_4046_6;

Selector_2 s4046_6(wires_1011_5[2], addr_1011_5, wires_4046_6,addr_4046_6);

wire[3:0] wires_4047_6;

wire[31:0] addr_4047_6;

Selector_2 s4047_6(wires_1011_5[3], addr_1011_5, wires_4047_6,addr_4047_6);

wire[3:0] wires_4048_6;

wire[31:0] addr_4048_6;

Selector_2 s4048_6(wires_1012_5[0], addr_1012_5, wires_4048_6,addr_4048_6);

wire[3:0] wires_4049_6;

wire[31:0] addr_4049_6;

Selector_2 s4049_6(wires_1012_5[1], addr_1012_5, wires_4049_6,addr_4049_6);

wire[3:0] wires_4050_6;

wire[31:0] addr_4050_6;

Selector_2 s4050_6(wires_1012_5[2], addr_1012_5, wires_4050_6,addr_4050_6);

wire[3:0] wires_4051_6;

wire[31:0] addr_4051_6;

Selector_2 s4051_6(wires_1012_5[3], addr_1012_5, wires_4051_6,addr_4051_6);

wire[3:0] wires_4052_6;

wire[31:0] addr_4052_6;

Selector_2 s4052_6(wires_1013_5[0], addr_1013_5, wires_4052_6,addr_4052_6);

wire[3:0] wires_4053_6;

wire[31:0] addr_4053_6;

Selector_2 s4053_6(wires_1013_5[1], addr_1013_5, wires_4053_6,addr_4053_6);

wire[3:0] wires_4054_6;

wire[31:0] addr_4054_6;

Selector_2 s4054_6(wires_1013_5[2], addr_1013_5, wires_4054_6,addr_4054_6);

wire[3:0] wires_4055_6;

wire[31:0] addr_4055_6;

Selector_2 s4055_6(wires_1013_5[3], addr_1013_5, wires_4055_6,addr_4055_6);

wire[3:0] wires_4056_6;

wire[31:0] addr_4056_6;

Selector_2 s4056_6(wires_1014_5[0], addr_1014_5, wires_4056_6,addr_4056_6);

wire[3:0] wires_4057_6;

wire[31:0] addr_4057_6;

Selector_2 s4057_6(wires_1014_5[1], addr_1014_5, wires_4057_6,addr_4057_6);

wire[3:0] wires_4058_6;

wire[31:0] addr_4058_6;

Selector_2 s4058_6(wires_1014_5[2], addr_1014_5, wires_4058_6,addr_4058_6);

wire[3:0] wires_4059_6;

wire[31:0] addr_4059_6;

Selector_2 s4059_6(wires_1014_5[3], addr_1014_5, wires_4059_6,addr_4059_6);

wire[3:0] wires_4060_6;

wire[31:0] addr_4060_6;

Selector_2 s4060_6(wires_1015_5[0], addr_1015_5, wires_4060_6,addr_4060_6);

wire[3:0] wires_4061_6;

wire[31:0] addr_4061_6;

Selector_2 s4061_6(wires_1015_5[1], addr_1015_5, wires_4061_6,addr_4061_6);

wire[3:0] wires_4062_6;

wire[31:0] addr_4062_6;

Selector_2 s4062_6(wires_1015_5[2], addr_1015_5, wires_4062_6,addr_4062_6);

wire[3:0] wires_4063_6;

wire[31:0] addr_4063_6;

Selector_2 s4063_6(wires_1015_5[3], addr_1015_5, wires_4063_6,addr_4063_6);

wire[3:0] wires_4064_6;

wire[31:0] addr_4064_6;

Selector_2 s4064_6(wires_1016_5[0], addr_1016_5, wires_4064_6,addr_4064_6);

wire[3:0] wires_4065_6;

wire[31:0] addr_4065_6;

Selector_2 s4065_6(wires_1016_5[1], addr_1016_5, wires_4065_6,addr_4065_6);

wire[3:0] wires_4066_6;

wire[31:0] addr_4066_6;

Selector_2 s4066_6(wires_1016_5[2], addr_1016_5, wires_4066_6,addr_4066_6);

wire[3:0] wires_4067_6;

wire[31:0] addr_4067_6;

Selector_2 s4067_6(wires_1016_5[3], addr_1016_5, wires_4067_6,addr_4067_6);

wire[3:0] wires_4068_6;

wire[31:0] addr_4068_6;

Selector_2 s4068_6(wires_1017_5[0], addr_1017_5, wires_4068_6,addr_4068_6);

wire[3:0] wires_4069_6;

wire[31:0] addr_4069_6;

Selector_2 s4069_6(wires_1017_5[1], addr_1017_5, wires_4069_6,addr_4069_6);

wire[3:0] wires_4070_6;

wire[31:0] addr_4070_6;

Selector_2 s4070_6(wires_1017_5[2], addr_1017_5, wires_4070_6,addr_4070_6);

wire[3:0] wires_4071_6;

wire[31:0] addr_4071_6;

Selector_2 s4071_6(wires_1017_5[3], addr_1017_5, wires_4071_6,addr_4071_6);

wire[3:0] wires_4072_6;

wire[31:0] addr_4072_6;

Selector_2 s4072_6(wires_1018_5[0], addr_1018_5, wires_4072_6,addr_4072_6);

wire[3:0] wires_4073_6;

wire[31:0] addr_4073_6;

Selector_2 s4073_6(wires_1018_5[1], addr_1018_5, wires_4073_6,addr_4073_6);

wire[3:0] wires_4074_6;

wire[31:0] addr_4074_6;

Selector_2 s4074_6(wires_1018_5[2], addr_1018_5, wires_4074_6,addr_4074_6);

wire[3:0] wires_4075_6;

wire[31:0] addr_4075_6;

Selector_2 s4075_6(wires_1018_5[3], addr_1018_5, wires_4075_6,addr_4075_6);

wire[3:0] wires_4076_6;

wire[31:0] addr_4076_6;

Selector_2 s4076_6(wires_1019_5[0], addr_1019_5, wires_4076_6,addr_4076_6);

wire[3:0] wires_4077_6;

wire[31:0] addr_4077_6;

Selector_2 s4077_6(wires_1019_5[1], addr_1019_5, wires_4077_6,addr_4077_6);

wire[3:0] wires_4078_6;

wire[31:0] addr_4078_6;

Selector_2 s4078_6(wires_1019_5[2], addr_1019_5, wires_4078_6,addr_4078_6);

wire[3:0] wires_4079_6;

wire[31:0] addr_4079_6;

Selector_2 s4079_6(wires_1019_5[3], addr_1019_5, wires_4079_6,addr_4079_6);

wire[3:0] wires_4080_6;

wire[31:0] addr_4080_6;

Selector_2 s4080_6(wires_1020_5[0], addr_1020_5, wires_4080_6,addr_4080_6);

wire[3:0] wires_4081_6;

wire[31:0] addr_4081_6;

Selector_2 s4081_6(wires_1020_5[1], addr_1020_5, wires_4081_6,addr_4081_6);

wire[3:0] wires_4082_6;

wire[31:0] addr_4082_6;

Selector_2 s4082_6(wires_1020_5[2], addr_1020_5, wires_4082_6,addr_4082_6);

wire[3:0] wires_4083_6;

wire[31:0] addr_4083_6;

Selector_2 s4083_6(wires_1020_5[3], addr_1020_5, wires_4083_6,addr_4083_6);

wire[3:0] wires_4084_6;

wire[31:0] addr_4084_6;

Selector_2 s4084_6(wires_1021_5[0], addr_1021_5, wires_4084_6,addr_4084_6);

wire[3:0] wires_4085_6;

wire[31:0] addr_4085_6;

Selector_2 s4085_6(wires_1021_5[1], addr_1021_5, wires_4085_6,addr_4085_6);

wire[3:0] wires_4086_6;

wire[31:0] addr_4086_6;

Selector_2 s4086_6(wires_1021_5[2], addr_1021_5, wires_4086_6,addr_4086_6);

wire[3:0] wires_4087_6;

wire[31:0] addr_4087_6;

Selector_2 s4087_6(wires_1021_5[3], addr_1021_5, wires_4087_6,addr_4087_6);

wire[3:0] wires_4088_6;

wire[31:0] addr_4088_6;

Selector_2 s4088_6(wires_1022_5[0], addr_1022_5, wires_4088_6,addr_4088_6);

wire[3:0] wires_4089_6;

wire[31:0] addr_4089_6;

Selector_2 s4089_6(wires_1022_5[1], addr_1022_5, wires_4089_6,addr_4089_6);

wire[3:0] wires_4090_6;

wire[31:0] addr_4090_6;

Selector_2 s4090_6(wires_1022_5[2], addr_1022_5, wires_4090_6,addr_4090_6);

wire[3:0] wires_4091_6;

wire[31:0] addr_4091_6;

Selector_2 s4091_6(wires_1022_5[3], addr_1022_5, wires_4091_6,addr_4091_6);

wire[3:0] wires_4092_6;

wire[31:0] addr_4092_6;

Selector_2 s4092_6(wires_1023_5[0], addr_1023_5, wires_4092_6,addr_4092_6);

wire[3:0] wires_4093_6;

wire[31:0] addr_4093_6;

Selector_2 s4093_6(wires_1023_5[1], addr_1023_5, wires_4093_6,addr_4093_6);

wire[3:0] wires_4094_6;

wire[31:0] addr_4094_6;

Selector_2 s4094_6(wires_1023_5[2], addr_1023_5, wires_4094_6,addr_4094_6);

wire[3:0] wires_4095_6;

wire[31:0] addr_4095_6;

Selector_2 s4095_6(wires_1023_5[3], addr_1023_5, wires_4095_6,addr_4095_6);

wire[31:0] addr_0_7;

Selector_2 s0_7(wires_0_6[0], addr_0_6, addr_positional[3:0], addr_0_7);

wire[31:0] addr_1_7;

Selector_2 s1_7(wires_0_6[1], addr_0_6, addr_positional[7:4], addr_1_7);

wire[31:0] addr_2_7;

Selector_2 s2_7(wires_0_6[2], addr_0_6, addr_positional[11:8], addr_2_7);

wire[31:0] addr_3_7;

Selector_2 s3_7(wires_0_6[3], addr_0_6, addr_positional[15:12], addr_3_7);

wire[31:0] addr_4_7;

Selector_2 s4_7(wires_1_6[0], addr_1_6, addr_positional[19:16], addr_4_7);

wire[31:0] addr_5_7;

Selector_2 s5_7(wires_1_6[1], addr_1_6, addr_positional[23:20], addr_5_7);

wire[31:0] addr_6_7;

Selector_2 s6_7(wires_1_6[2], addr_1_6, addr_positional[27:24], addr_6_7);

wire[31:0] addr_7_7;

Selector_2 s7_7(wires_1_6[3], addr_1_6, addr_positional[31:28], addr_7_7);

wire[31:0] addr_8_7;

Selector_2 s8_7(wires_2_6[0], addr_2_6, addr_positional[35:32], addr_8_7);

wire[31:0] addr_9_7;

Selector_2 s9_7(wires_2_6[1], addr_2_6, addr_positional[39:36], addr_9_7);

wire[31:0] addr_10_7;

Selector_2 s10_7(wires_2_6[2], addr_2_6, addr_positional[43:40], addr_10_7);

wire[31:0] addr_11_7;

Selector_2 s11_7(wires_2_6[3], addr_2_6, addr_positional[47:44], addr_11_7);

wire[31:0] addr_12_7;

Selector_2 s12_7(wires_3_6[0], addr_3_6, addr_positional[51:48], addr_12_7);

wire[31:0] addr_13_7;

Selector_2 s13_7(wires_3_6[1], addr_3_6, addr_positional[55:52], addr_13_7);

wire[31:0] addr_14_7;

Selector_2 s14_7(wires_3_6[2], addr_3_6, addr_positional[59:56], addr_14_7);

wire[31:0] addr_15_7;

Selector_2 s15_7(wires_3_6[3], addr_3_6, addr_positional[63:60], addr_15_7);

wire[31:0] addr_16_7;

Selector_2 s16_7(wires_4_6[0], addr_4_6, addr_positional[67:64], addr_16_7);

wire[31:0] addr_17_7;

Selector_2 s17_7(wires_4_6[1], addr_4_6, addr_positional[71:68], addr_17_7);

wire[31:0] addr_18_7;

Selector_2 s18_7(wires_4_6[2], addr_4_6, addr_positional[75:72], addr_18_7);

wire[31:0] addr_19_7;

Selector_2 s19_7(wires_4_6[3], addr_4_6, addr_positional[79:76], addr_19_7);

wire[31:0] addr_20_7;

Selector_2 s20_7(wires_5_6[0], addr_5_6, addr_positional[83:80], addr_20_7);

wire[31:0] addr_21_7;

Selector_2 s21_7(wires_5_6[1], addr_5_6, addr_positional[87:84], addr_21_7);

wire[31:0] addr_22_7;

Selector_2 s22_7(wires_5_6[2], addr_5_6, addr_positional[91:88], addr_22_7);

wire[31:0] addr_23_7;

Selector_2 s23_7(wires_5_6[3], addr_5_6, addr_positional[95:92], addr_23_7);

wire[31:0] addr_24_7;

Selector_2 s24_7(wires_6_6[0], addr_6_6, addr_positional[99:96], addr_24_7);

wire[31:0] addr_25_7;

Selector_2 s25_7(wires_6_6[1], addr_6_6, addr_positional[103:100], addr_25_7);

wire[31:0] addr_26_7;

Selector_2 s26_7(wires_6_6[2], addr_6_6, addr_positional[107:104], addr_26_7);

wire[31:0] addr_27_7;

Selector_2 s27_7(wires_6_6[3], addr_6_6, addr_positional[111:108], addr_27_7);

wire[31:0] addr_28_7;

Selector_2 s28_7(wires_7_6[0], addr_7_6, addr_positional[115:112], addr_28_7);

wire[31:0] addr_29_7;

Selector_2 s29_7(wires_7_6[1], addr_7_6, addr_positional[119:116], addr_29_7);

wire[31:0] addr_30_7;

Selector_2 s30_7(wires_7_6[2], addr_7_6, addr_positional[123:120], addr_30_7);

wire[31:0] addr_31_7;

Selector_2 s31_7(wires_7_6[3], addr_7_6, addr_positional[127:124], addr_31_7);

wire[31:0] addr_32_7;

Selector_2 s32_7(wires_8_6[0], addr_8_6, addr_positional[131:128], addr_32_7);

wire[31:0] addr_33_7;

Selector_2 s33_7(wires_8_6[1], addr_8_6, addr_positional[135:132], addr_33_7);

wire[31:0] addr_34_7;

Selector_2 s34_7(wires_8_6[2], addr_8_6, addr_positional[139:136], addr_34_7);

wire[31:0] addr_35_7;

Selector_2 s35_7(wires_8_6[3], addr_8_6, addr_positional[143:140], addr_35_7);

wire[31:0] addr_36_7;

Selector_2 s36_7(wires_9_6[0], addr_9_6, addr_positional[147:144], addr_36_7);

wire[31:0] addr_37_7;

Selector_2 s37_7(wires_9_6[1], addr_9_6, addr_positional[151:148], addr_37_7);

wire[31:0] addr_38_7;

Selector_2 s38_7(wires_9_6[2], addr_9_6, addr_positional[155:152], addr_38_7);

wire[31:0] addr_39_7;

Selector_2 s39_7(wires_9_6[3], addr_9_6, addr_positional[159:156], addr_39_7);

wire[31:0] addr_40_7;

Selector_2 s40_7(wires_10_6[0], addr_10_6, addr_positional[163:160], addr_40_7);

wire[31:0] addr_41_7;

Selector_2 s41_7(wires_10_6[1], addr_10_6, addr_positional[167:164], addr_41_7);

wire[31:0] addr_42_7;

Selector_2 s42_7(wires_10_6[2], addr_10_6, addr_positional[171:168], addr_42_7);

wire[31:0] addr_43_7;

Selector_2 s43_7(wires_10_6[3], addr_10_6, addr_positional[175:172], addr_43_7);

wire[31:0] addr_44_7;

Selector_2 s44_7(wires_11_6[0], addr_11_6, addr_positional[179:176], addr_44_7);

wire[31:0] addr_45_7;

Selector_2 s45_7(wires_11_6[1], addr_11_6, addr_positional[183:180], addr_45_7);

wire[31:0] addr_46_7;

Selector_2 s46_7(wires_11_6[2], addr_11_6, addr_positional[187:184], addr_46_7);

wire[31:0] addr_47_7;

Selector_2 s47_7(wires_11_6[3], addr_11_6, addr_positional[191:188], addr_47_7);

wire[31:0] addr_48_7;

Selector_2 s48_7(wires_12_6[0], addr_12_6, addr_positional[195:192], addr_48_7);

wire[31:0] addr_49_7;

Selector_2 s49_7(wires_12_6[1], addr_12_6, addr_positional[199:196], addr_49_7);

wire[31:0] addr_50_7;

Selector_2 s50_7(wires_12_6[2], addr_12_6, addr_positional[203:200], addr_50_7);

wire[31:0] addr_51_7;

Selector_2 s51_7(wires_12_6[3], addr_12_6, addr_positional[207:204], addr_51_7);

wire[31:0] addr_52_7;

Selector_2 s52_7(wires_13_6[0], addr_13_6, addr_positional[211:208], addr_52_7);

wire[31:0] addr_53_7;

Selector_2 s53_7(wires_13_6[1], addr_13_6, addr_positional[215:212], addr_53_7);

wire[31:0] addr_54_7;

Selector_2 s54_7(wires_13_6[2], addr_13_6, addr_positional[219:216], addr_54_7);

wire[31:0] addr_55_7;

Selector_2 s55_7(wires_13_6[3], addr_13_6, addr_positional[223:220], addr_55_7);

wire[31:0] addr_56_7;

Selector_2 s56_7(wires_14_6[0], addr_14_6, addr_positional[227:224], addr_56_7);

wire[31:0] addr_57_7;

Selector_2 s57_7(wires_14_6[1], addr_14_6, addr_positional[231:228], addr_57_7);

wire[31:0] addr_58_7;

Selector_2 s58_7(wires_14_6[2], addr_14_6, addr_positional[235:232], addr_58_7);

wire[31:0] addr_59_7;

Selector_2 s59_7(wires_14_6[3], addr_14_6, addr_positional[239:236], addr_59_7);

wire[31:0] addr_60_7;

Selector_2 s60_7(wires_15_6[0], addr_15_6, addr_positional[243:240], addr_60_7);

wire[31:0] addr_61_7;

Selector_2 s61_7(wires_15_6[1], addr_15_6, addr_positional[247:244], addr_61_7);

wire[31:0] addr_62_7;

Selector_2 s62_7(wires_15_6[2], addr_15_6, addr_positional[251:248], addr_62_7);

wire[31:0] addr_63_7;

Selector_2 s63_7(wires_15_6[3], addr_15_6, addr_positional[255:252], addr_63_7);

wire[31:0] addr_64_7;

Selector_2 s64_7(wires_16_6[0], addr_16_6, addr_positional[259:256], addr_64_7);

wire[31:0] addr_65_7;

Selector_2 s65_7(wires_16_6[1], addr_16_6, addr_positional[263:260], addr_65_7);

wire[31:0] addr_66_7;

Selector_2 s66_7(wires_16_6[2], addr_16_6, addr_positional[267:264], addr_66_7);

wire[31:0] addr_67_7;

Selector_2 s67_7(wires_16_6[3], addr_16_6, addr_positional[271:268], addr_67_7);

wire[31:0] addr_68_7;

Selector_2 s68_7(wires_17_6[0], addr_17_6, addr_positional[275:272], addr_68_7);

wire[31:0] addr_69_7;

Selector_2 s69_7(wires_17_6[1], addr_17_6, addr_positional[279:276], addr_69_7);

wire[31:0] addr_70_7;

Selector_2 s70_7(wires_17_6[2], addr_17_6, addr_positional[283:280], addr_70_7);

wire[31:0] addr_71_7;

Selector_2 s71_7(wires_17_6[3], addr_17_6, addr_positional[287:284], addr_71_7);

wire[31:0] addr_72_7;

Selector_2 s72_7(wires_18_6[0], addr_18_6, addr_positional[291:288], addr_72_7);

wire[31:0] addr_73_7;

Selector_2 s73_7(wires_18_6[1], addr_18_6, addr_positional[295:292], addr_73_7);

wire[31:0] addr_74_7;

Selector_2 s74_7(wires_18_6[2], addr_18_6, addr_positional[299:296], addr_74_7);

wire[31:0] addr_75_7;

Selector_2 s75_7(wires_18_6[3], addr_18_6, addr_positional[303:300], addr_75_7);

wire[31:0] addr_76_7;

Selector_2 s76_7(wires_19_6[0], addr_19_6, addr_positional[307:304], addr_76_7);

wire[31:0] addr_77_7;

Selector_2 s77_7(wires_19_6[1], addr_19_6, addr_positional[311:308], addr_77_7);

wire[31:0] addr_78_7;

Selector_2 s78_7(wires_19_6[2], addr_19_6, addr_positional[315:312], addr_78_7);

wire[31:0] addr_79_7;

Selector_2 s79_7(wires_19_6[3], addr_19_6, addr_positional[319:316], addr_79_7);

wire[31:0] addr_80_7;

Selector_2 s80_7(wires_20_6[0], addr_20_6, addr_positional[323:320], addr_80_7);

wire[31:0] addr_81_7;

Selector_2 s81_7(wires_20_6[1], addr_20_6, addr_positional[327:324], addr_81_7);

wire[31:0] addr_82_7;

Selector_2 s82_7(wires_20_6[2], addr_20_6, addr_positional[331:328], addr_82_7);

wire[31:0] addr_83_7;

Selector_2 s83_7(wires_20_6[3], addr_20_6, addr_positional[335:332], addr_83_7);

wire[31:0] addr_84_7;

Selector_2 s84_7(wires_21_6[0], addr_21_6, addr_positional[339:336], addr_84_7);

wire[31:0] addr_85_7;

Selector_2 s85_7(wires_21_6[1], addr_21_6, addr_positional[343:340], addr_85_7);

wire[31:0] addr_86_7;

Selector_2 s86_7(wires_21_6[2], addr_21_6, addr_positional[347:344], addr_86_7);

wire[31:0] addr_87_7;

Selector_2 s87_7(wires_21_6[3], addr_21_6, addr_positional[351:348], addr_87_7);

wire[31:0] addr_88_7;

Selector_2 s88_7(wires_22_6[0], addr_22_6, addr_positional[355:352], addr_88_7);

wire[31:0] addr_89_7;

Selector_2 s89_7(wires_22_6[1], addr_22_6, addr_positional[359:356], addr_89_7);

wire[31:0] addr_90_7;

Selector_2 s90_7(wires_22_6[2], addr_22_6, addr_positional[363:360], addr_90_7);

wire[31:0] addr_91_7;

Selector_2 s91_7(wires_22_6[3], addr_22_6, addr_positional[367:364], addr_91_7);

wire[31:0] addr_92_7;

Selector_2 s92_7(wires_23_6[0], addr_23_6, addr_positional[371:368], addr_92_7);

wire[31:0] addr_93_7;

Selector_2 s93_7(wires_23_6[1], addr_23_6, addr_positional[375:372], addr_93_7);

wire[31:0] addr_94_7;

Selector_2 s94_7(wires_23_6[2], addr_23_6, addr_positional[379:376], addr_94_7);

wire[31:0] addr_95_7;

Selector_2 s95_7(wires_23_6[3], addr_23_6, addr_positional[383:380], addr_95_7);

wire[31:0] addr_96_7;

Selector_2 s96_7(wires_24_6[0], addr_24_6, addr_positional[387:384], addr_96_7);

wire[31:0] addr_97_7;

Selector_2 s97_7(wires_24_6[1], addr_24_6, addr_positional[391:388], addr_97_7);

wire[31:0] addr_98_7;

Selector_2 s98_7(wires_24_6[2], addr_24_6, addr_positional[395:392], addr_98_7);

wire[31:0] addr_99_7;

Selector_2 s99_7(wires_24_6[3], addr_24_6, addr_positional[399:396], addr_99_7);

wire[31:0] addr_100_7;

Selector_2 s100_7(wires_25_6[0], addr_25_6, addr_positional[403:400], addr_100_7);

wire[31:0] addr_101_7;

Selector_2 s101_7(wires_25_6[1], addr_25_6, addr_positional[407:404], addr_101_7);

wire[31:0] addr_102_7;

Selector_2 s102_7(wires_25_6[2], addr_25_6, addr_positional[411:408], addr_102_7);

wire[31:0] addr_103_7;

Selector_2 s103_7(wires_25_6[3], addr_25_6, addr_positional[415:412], addr_103_7);

wire[31:0] addr_104_7;

Selector_2 s104_7(wires_26_6[0], addr_26_6, addr_positional[419:416], addr_104_7);

wire[31:0] addr_105_7;

Selector_2 s105_7(wires_26_6[1], addr_26_6, addr_positional[423:420], addr_105_7);

wire[31:0] addr_106_7;

Selector_2 s106_7(wires_26_6[2], addr_26_6, addr_positional[427:424], addr_106_7);

wire[31:0] addr_107_7;

Selector_2 s107_7(wires_26_6[3], addr_26_6, addr_positional[431:428], addr_107_7);

wire[31:0] addr_108_7;

Selector_2 s108_7(wires_27_6[0], addr_27_6, addr_positional[435:432], addr_108_7);

wire[31:0] addr_109_7;

Selector_2 s109_7(wires_27_6[1], addr_27_6, addr_positional[439:436], addr_109_7);

wire[31:0] addr_110_7;

Selector_2 s110_7(wires_27_6[2], addr_27_6, addr_positional[443:440], addr_110_7);

wire[31:0] addr_111_7;

Selector_2 s111_7(wires_27_6[3], addr_27_6, addr_positional[447:444], addr_111_7);

wire[31:0] addr_112_7;

Selector_2 s112_7(wires_28_6[0], addr_28_6, addr_positional[451:448], addr_112_7);

wire[31:0] addr_113_7;

Selector_2 s113_7(wires_28_6[1], addr_28_6, addr_positional[455:452], addr_113_7);

wire[31:0] addr_114_7;

Selector_2 s114_7(wires_28_6[2], addr_28_6, addr_positional[459:456], addr_114_7);

wire[31:0] addr_115_7;

Selector_2 s115_7(wires_28_6[3], addr_28_6, addr_positional[463:460], addr_115_7);

wire[31:0] addr_116_7;

Selector_2 s116_7(wires_29_6[0], addr_29_6, addr_positional[467:464], addr_116_7);

wire[31:0] addr_117_7;

Selector_2 s117_7(wires_29_6[1], addr_29_6, addr_positional[471:468], addr_117_7);

wire[31:0] addr_118_7;

Selector_2 s118_7(wires_29_6[2], addr_29_6, addr_positional[475:472], addr_118_7);

wire[31:0] addr_119_7;

Selector_2 s119_7(wires_29_6[3], addr_29_6, addr_positional[479:476], addr_119_7);

wire[31:0] addr_120_7;

Selector_2 s120_7(wires_30_6[0], addr_30_6, addr_positional[483:480], addr_120_7);

wire[31:0] addr_121_7;

Selector_2 s121_7(wires_30_6[1], addr_30_6, addr_positional[487:484], addr_121_7);

wire[31:0] addr_122_7;

Selector_2 s122_7(wires_30_6[2], addr_30_6, addr_positional[491:488], addr_122_7);

wire[31:0] addr_123_7;

Selector_2 s123_7(wires_30_6[3], addr_30_6, addr_positional[495:492], addr_123_7);

wire[31:0] addr_124_7;

Selector_2 s124_7(wires_31_6[0], addr_31_6, addr_positional[499:496], addr_124_7);

wire[31:0] addr_125_7;

Selector_2 s125_7(wires_31_6[1], addr_31_6, addr_positional[503:500], addr_125_7);

wire[31:0] addr_126_7;

Selector_2 s126_7(wires_31_6[2], addr_31_6, addr_positional[507:504], addr_126_7);

wire[31:0] addr_127_7;

Selector_2 s127_7(wires_31_6[3], addr_31_6, addr_positional[511:508], addr_127_7);

wire[31:0] addr_128_7;

Selector_2 s128_7(wires_32_6[0], addr_32_6, addr_positional[515:512], addr_128_7);

wire[31:0] addr_129_7;

Selector_2 s129_7(wires_32_6[1], addr_32_6, addr_positional[519:516], addr_129_7);

wire[31:0] addr_130_7;

Selector_2 s130_7(wires_32_6[2], addr_32_6, addr_positional[523:520], addr_130_7);

wire[31:0] addr_131_7;

Selector_2 s131_7(wires_32_6[3], addr_32_6, addr_positional[527:524], addr_131_7);

wire[31:0] addr_132_7;

Selector_2 s132_7(wires_33_6[0], addr_33_6, addr_positional[531:528], addr_132_7);

wire[31:0] addr_133_7;

Selector_2 s133_7(wires_33_6[1], addr_33_6, addr_positional[535:532], addr_133_7);

wire[31:0] addr_134_7;

Selector_2 s134_7(wires_33_6[2], addr_33_6, addr_positional[539:536], addr_134_7);

wire[31:0] addr_135_7;

Selector_2 s135_7(wires_33_6[3], addr_33_6, addr_positional[543:540], addr_135_7);

wire[31:0] addr_136_7;

Selector_2 s136_7(wires_34_6[0], addr_34_6, addr_positional[547:544], addr_136_7);

wire[31:0] addr_137_7;

Selector_2 s137_7(wires_34_6[1], addr_34_6, addr_positional[551:548], addr_137_7);

wire[31:0] addr_138_7;

Selector_2 s138_7(wires_34_6[2], addr_34_6, addr_positional[555:552], addr_138_7);

wire[31:0] addr_139_7;

Selector_2 s139_7(wires_34_6[3], addr_34_6, addr_positional[559:556], addr_139_7);

wire[31:0] addr_140_7;

Selector_2 s140_7(wires_35_6[0], addr_35_6, addr_positional[563:560], addr_140_7);

wire[31:0] addr_141_7;

Selector_2 s141_7(wires_35_6[1], addr_35_6, addr_positional[567:564], addr_141_7);

wire[31:0] addr_142_7;

Selector_2 s142_7(wires_35_6[2], addr_35_6, addr_positional[571:568], addr_142_7);

wire[31:0] addr_143_7;

Selector_2 s143_7(wires_35_6[3], addr_35_6, addr_positional[575:572], addr_143_7);

wire[31:0] addr_144_7;

Selector_2 s144_7(wires_36_6[0], addr_36_6, addr_positional[579:576], addr_144_7);

wire[31:0] addr_145_7;

Selector_2 s145_7(wires_36_6[1], addr_36_6, addr_positional[583:580], addr_145_7);

wire[31:0] addr_146_7;

Selector_2 s146_7(wires_36_6[2], addr_36_6, addr_positional[587:584], addr_146_7);

wire[31:0] addr_147_7;

Selector_2 s147_7(wires_36_6[3], addr_36_6, addr_positional[591:588], addr_147_7);

wire[31:0] addr_148_7;

Selector_2 s148_7(wires_37_6[0], addr_37_6, addr_positional[595:592], addr_148_7);

wire[31:0] addr_149_7;

Selector_2 s149_7(wires_37_6[1], addr_37_6, addr_positional[599:596], addr_149_7);

wire[31:0] addr_150_7;

Selector_2 s150_7(wires_37_6[2], addr_37_6, addr_positional[603:600], addr_150_7);

wire[31:0] addr_151_7;

Selector_2 s151_7(wires_37_6[3], addr_37_6, addr_positional[607:604], addr_151_7);

wire[31:0] addr_152_7;

Selector_2 s152_7(wires_38_6[0], addr_38_6, addr_positional[611:608], addr_152_7);

wire[31:0] addr_153_7;

Selector_2 s153_7(wires_38_6[1], addr_38_6, addr_positional[615:612], addr_153_7);

wire[31:0] addr_154_7;

Selector_2 s154_7(wires_38_6[2], addr_38_6, addr_positional[619:616], addr_154_7);

wire[31:0] addr_155_7;

Selector_2 s155_7(wires_38_6[3], addr_38_6, addr_positional[623:620], addr_155_7);

wire[31:0] addr_156_7;

Selector_2 s156_7(wires_39_6[0], addr_39_6, addr_positional[627:624], addr_156_7);

wire[31:0] addr_157_7;

Selector_2 s157_7(wires_39_6[1], addr_39_6, addr_positional[631:628], addr_157_7);

wire[31:0] addr_158_7;

Selector_2 s158_7(wires_39_6[2], addr_39_6, addr_positional[635:632], addr_158_7);

wire[31:0] addr_159_7;

Selector_2 s159_7(wires_39_6[3], addr_39_6, addr_positional[639:636], addr_159_7);

wire[31:0] addr_160_7;

Selector_2 s160_7(wires_40_6[0], addr_40_6, addr_positional[643:640], addr_160_7);

wire[31:0] addr_161_7;

Selector_2 s161_7(wires_40_6[1], addr_40_6, addr_positional[647:644], addr_161_7);

wire[31:0] addr_162_7;

Selector_2 s162_7(wires_40_6[2], addr_40_6, addr_positional[651:648], addr_162_7);

wire[31:0] addr_163_7;

Selector_2 s163_7(wires_40_6[3], addr_40_6, addr_positional[655:652], addr_163_7);

wire[31:0] addr_164_7;

Selector_2 s164_7(wires_41_6[0], addr_41_6, addr_positional[659:656], addr_164_7);

wire[31:0] addr_165_7;

Selector_2 s165_7(wires_41_6[1], addr_41_6, addr_positional[663:660], addr_165_7);

wire[31:0] addr_166_7;

Selector_2 s166_7(wires_41_6[2], addr_41_6, addr_positional[667:664], addr_166_7);

wire[31:0] addr_167_7;

Selector_2 s167_7(wires_41_6[3], addr_41_6, addr_positional[671:668], addr_167_7);

wire[31:0] addr_168_7;

Selector_2 s168_7(wires_42_6[0], addr_42_6, addr_positional[675:672], addr_168_7);

wire[31:0] addr_169_7;

Selector_2 s169_7(wires_42_6[1], addr_42_6, addr_positional[679:676], addr_169_7);

wire[31:0] addr_170_7;

Selector_2 s170_7(wires_42_6[2], addr_42_6, addr_positional[683:680], addr_170_7);

wire[31:0] addr_171_7;

Selector_2 s171_7(wires_42_6[3], addr_42_6, addr_positional[687:684], addr_171_7);

wire[31:0] addr_172_7;

Selector_2 s172_7(wires_43_6[0], addr_43_6, addr_positional[691:688], addr_172_7);

wire[31:0] addr_173_7;

Selector_2 s173_7(wires_43_6[1], addr_43_6, addr_positional[695:692], addr_173_7);

wire[31:0] addr_174_7;

Selector_2 s174_7(wires_43_6[2], addr_43_6, addr_positional[699:696], addr_174_7);

wire[31:0] addr_175_7;

Selector_2 s175_7(wires_43_6[3], addr_43_6, addr_positional[703:700], addr_175_7);

wire[31:0] addr_176_7;

Selector_2 s176_7(wires_44_6[0], addr_44_6, addr_positional[707:704], addr_176_7);

wire[31:0] addr_177_7;

Selector_2 s177_7(wires_44_6[1], addr_44_6, addr_positional[711:708], addr_177_7);

wire[31:0] addr_178_7;

Selector_2 s178_7(wires_44_6[2], addr_44_6, addr_positional[715:712], addr_178_7);

wire[31:0] addr_179_7;

Selector_2 s179_7(wires_44_6[3], addr_44_6, addr_positional[719:716], addr_179_7);

wire[31:0] addr_180_7;

Selector_2 s180_7(wires_45_6[0], addr_45_6, addr_positional[723:720], addr_180_7);

wire[31:0] addr_181_7;

Selector_2 s181_7(wires_45_6[1], addr_45_6, addr_positional[727:724], addr_181_7);

wire[31:0] addr_182_7;

Selector_2 s182_7(wires_45_6[2], addr_45_6, addr_positional[731:728], addr_182_7);

wire[31:0] addr_183_7;

Selector_2 s183_7(wires_45_6[3], addr_45_6, addr_positional[735:732], addr_183_7);

wire[31:0] addr_184_7;

Selector_2 s184_7(wires_46_6[0], addr_46_6, addr_positional[739:736], addr_184_7);

wire[31:0] addr_185_7;

Selector_2 s185_7(wires_46_6[1], addr_46_6, addr_positional[743:740], addr_185_7);

wire[31:0] addr_186_7;

Selector_2 s186_7(wires_46_6[2], addr_46_6, addr_positional[747:744], addr_186_7);

wire[31:0] addr_187_7;

Selector_2 s187_7(wires_46_6[3], addr_46_6, addr_positional[751:748], addr_187_7);

wire[31:0] addr_188_7;

Selector_2 s188_7(wires_47_6[0], addr_47_6, addr_positional[755:752], addr_188_7);

wire[31:0] addr_189_7;

Selector_2 s189_7(wires_47_6[1], addr_47_6, addr_positional[759:756], addr_189_7);

wire[31:0] addr_190_7;

Selector_2 s190_7(wires_47_6[2], addr_47_6, addr_positional[763:760], addr_190_7);

wire[31:0] addr_191_7;

Selector_2 s191_7(wires_47_6[3], addr_47_6, addr_positional[767:764], addr_191_7);

wire[31:0] addr_192_7;

Selector_2 s192_7(wires_48_6[0], addr_48_6, addr_positional[771:768], addr_192_7);

wire[31:0] addr_193_7;

Selector_2 s193_7(wires_48_6[1], addr_48_6, addr_positional[775:772], addr_193_7);

wire[31:0] addr_194_7;

Selector_2 s194_7(wires_48_6[2], addr_48_6, addr_positional[779:776], addr_194_7);

wire[31:0] addr_195_7;

Selector_2 s195_7(wires_48_6[3], addr_48_6, addr_positional[783:780], addr_195_7);

wire[31:0] addr_196_7;

Selector_2 s196_7(wires_49_6[0], addr_49_6, addr_positional[787:784], addr_196_7);

wire[31:0] addr_197_7;

Selector_2 s197_7(wires_49_6[1], addr_49_6, addr_positional[791:788], addr_197_7);

wire[31:0] addr_198_7;

Selector_2 s198_7(wires_49_6[2], addr_49_6, addr_positional[795:792], addr_198_7);

wire[31:0] addr_199_7;

Selector_2 s199_7(wires_49_6[3], addr_49_6, addr_positional[799:796], addr_199_7);

wire[31:0] addr_200_7;

Selector_2 s200_7(wires_50_6[0], addr_50_6, addr_positional[803:800], addr_200_7);

wire[31:0] addr_201_7;

Selector_2 s201_7(wires_50_6[1], addr_50_6, addr_positional[807:804], addr_201_7);

wire[31:0] addr_202_7;

Selector_2 s202_7(wires_50_6[2], addr_50_6, addr_positional[811:808], addr_202_7);

wire[31:0] addr_203_7;

Selector_2 s203_7(wires_50_6[3], addr_50_6, addr_positional[815:812], addr_203_7);

wire[31:0] addr_204_7;

Selector_2 s204_7(wires_51_6[0], addr_51_6, addr_positional[819:816], addr_204_7);

wire[31:0] addr_205_7;

Selector_2 s205_7(wires_51_6[1], addr_51_6, addr_positional[823:820], addr_205_7);

wire[31:0] addr_206_7;

Selector_2 s206_7(wires_51_6[2], addr_51_6, addr_positional[827:824], addr_206_7);

wire[31:0] addr_207_7;

Selector_2 s207_7(wires_51_6[3], addr_51_6, addr_positional[831:828], addr_207_7);

wire[31:0] addr_208_7;

Selector_2 s208_7(wires_52_6[0], addr_52_6, addr_positional[835:832], addr_208_7);

wire[31:0] addr_209_7;

Selector_2 s209_7(wires_52_6[1], addr_52_6, addr_positional[839:836], addr_209_7);

wire[31:0] addr_210_7;

Selector_2 s210_7(wires_52_6[2], addr_52_6, addr_positional[843:840], addr_210_7);

wire[31:0] addr_211_7;

Selector_2 s211_7(wires_52_6[3], addr_52_6, addr_positional[847:844], addr_211_7);

wire[31:0] addr_212_7;

Selector_2 s212_7(wires_53_6[0], addr_53_6, addr_positional[851:848], addr_212_7);

wire[31:0] addr_213_7;

Selector_2 s213_7(wires_53_6[1], addr_53_6, addr_positional[855:852], addr_213_7);

wire[31:0] addr_214_7;

Selector_2 s214_7(wires_53_6[2], addr_53_6, addr_positional[859:856], addr_214_7);

wire[31:0] addr_215_7;

Selector_2 s215_7(wires_53_6[3], addr_53_6, addr_positional[863:860], addr_215_7);

wire[31:0] addr_216_7;

Selector_2 s216_7(wires_54_6[0], addr_54_6, addr_positional[867:864], addr_216_7);

wire[31:0] addr_217_7;

Selector_2 s217_7(wires_54_6[1], addr_54_6, addr_positional[871:868], addr_217_7);

wire[31:0] addr_218_7;

Selector_2 s218_7(wires_54_6[2], addr_54_6, addr_positional[875:872], addr_218_7);

wire[31:0] addr_219_7;

Selector_2 s219_7(wires_54_6[3], addr_54_6, addr_positional[879:876], addr_219_7);

wire[31:0] addr_220_7;

Selector_2 s220_7(wires_55_6[0], addr_55_6, addr_positional[883:880], addr_220_7);

wire[31:0] addr_221_7;

Selector_2 s221_7(wires_55_6[1], addr_55_6, addr_positional[887:884], addr_221_7);

wire[31:0] addr_222_7;

Selector_2 s222_7(wires_55_6[2], addr_55_6, addr_positional[891:888], addr_222_7);

wire[31:0] addr_223_7;

Selector_2 s223_7(wires_55_6[3], addr_55_6, addr_positional[895:892], addr_223_7);

wire[31:0] addr_224_7;

Selector_2 s224_7(wires_56_6[0], addr_56_6, addr_positional[899:896], addr_224_7);

wire[31:0] addr_225_7;

Selector_2 s225_7(wires_56_6[1], addr_56_6, addr_positional[903:900], addr_225_7);

wire[31:0] addr_226_7;

Selector_2 s226_7(wires_56_6[2], addr_56_6, addr_positional[907:904], addr_226_7);

wire[31:0] addr_227_7;

Selector_2 s227_7(wires_56_6[3], addr_56_6, addr_positional[911:908], addr_227_7);

wire[31:0] addr_228_7;

Selector_2 s228_7(wires_57_6[0], addr_57_6, addr_positional[915:912], addr_228_7);

wire[31:0] addr_229_7;

Selector_2 s229_7(wires_57_6[1], addr_57_6, addr_positional[919:916], addr_229_7);

wire[31:0] addr_230_7;

Selector_2 s230_7(wires_57_6[2], addr_57_6, addr_positional[923:920], addr_230_7);

wire[31:0] addr_231_7;

Selector_2 s231_7(wires_57_6[3], addr_57_6, addr_positional[927:924], addr_231_7);

wire[31:0] addr_232_7;

Selector_2 s232_7(wires_58_6[0], addr_58_6, addr_positional[931:928], addr_232_7);

wire[31:0] addr_233_7;

Selector_2 s233_7(wires_58_6[1], addr_58_6, addr_positional[935:932], addr_233_7);

wire[31:0] addr_234_7;

Selector_2 s234_7(wires_58_6[2], addr_58_6, addr_positional[939:936], addr_234_7);

wire[31:0] addr_235_7;

Selector_2 s235_7(wires_58_6[3], addr_58_6, addr_positional[943:940], addr_235_7);

wire[31:0] addr_236_7;

Selector_2 s236_7(wires_59_6[0], addr_59_6, addr_positional[947:944], addr_236_7);

wire[31:0] addr_237_7;

Selector_2 s237_7(wires_59_6[1], addr_59_6, addr_positional[951:948], addr_237_7);

wire[31:0] addr_238_7;

Selector_2 s238_7(wires_59_6[2], addr_59_6, addr_positional[955:952], addr_238_7);

wire[31:0] addr_239_7;

Selector_2 s239_7(wires_59_6[3], addr_59_6, addr_positional[959:956], addr_239_7);

wire[31:0] addr_240_7;

Selector_2 s240_7(wires_60_6[0], addr_60_6, addr_positional[963:960], addr_240_7);

wire[31:0] addr_241_7;

Selector_2 s241_7(wires_60_6[1], addr_60_6, addr_positional[967:964], addr_241_7);

wire[31:0] addr_242_7;

Selector_2 s242_7(wires_60_6[2], addr_60_6, addr_positional[971:968], addr_242_7);

wire[31:0] addr_243_7;

Selector_2 s243_7(wires_60_6[3], addr_60_6, addr_positional[975:972], addr_243_7);

wire[31:0] addr_244_7;

Selector_2 s244_7(wires_61_6[0], addr_61_6, addr_positional[979:976], addr_244_7);

wire[31:0] addr_245_7;

Selector_2 s245_7(wires_61_6[1], addr_61_6, addr_positional[983:980], addr_245_7);

wire[31:0] addr_246_7;

Selector_2 s246_7(wires_61_6[2], addr_61_6, addr_positional[987:984], addr_246_7);

wire[31:0] addr_247_7;

Selector_2 s247_7(wires_61_6[3], addr_61_6, addr_positional[991:988], addr_247_7);

wire[31:0] addr_248_7;

Selector_2 s248_7(wires_62_6[0], addr_62_6, addr_positional[995:992], addr_248_7);

wire[31:0] addr_249_7;

Selector_2 s249_7(wires_62_6[1], addr_62_6, addr_positional[999:996], addr_249_7);

wire[31:0] addr_250_7;

Selector_2 s250_7(wires_62_6[2], addr_62_6, addr_positional[1003:1000], addr_250_7);

wire[31:0] addr_251_7;

Selector_2 s251_7(wires_62_6[3], addr_62_6, addr_positional[1007:1004], addr_251_7);

wire[31:0] addr_252_7;

Selector_2 s252_7(wires_63_6[0], addr_63_6, addr_positional[1011:1008], addr_252_7);

wire[31:0] addr_253_7;

Selector_2 s253_7(wires_63_6[1], addr_63_6, addr_positional[1015:1012], addr_253_7);

wire[31:0] addr_254_7;

Selector_2 s254_7(wires_63_6[2], addr_63_6, addr_positional[1019:1016], addr_254_7);

wire[31:0] addr_255_7;

Selector_2 s255_7(wires_63_6[3], addr_63_6, addr_positional[1023:1020], addr_255_7);

wire[31:0] addr_256_7;

Selector_2 s256_7(wires_64_6[0], addr_64_6, addr_positional[1027:1024], addr_256_7);

wire[31:0] addr_257_7;

Selector_2 s257_7(wires_64_6[1], addr_64_6, addr_positional[1031:1028], addr_257_7);

wire[31:0] addr_258_7;

Selector_2 s258_7(wires_64_6[2], addr_64_6, addr_positional[1035:1032], addr_258_7);

wire[31:0] addr_259_7;

Selector_2 s259_7(wires_64_6[3], addr_64_6, addr_positional[1039:1036], addr_259_7);

wire[31:0] addr_260_7;

Selector_2 s260_7(wires_65_6[0], addr_65_6, addr_positional[1043:1040], addr_260_7);

wire[31:0] addr_261_7;

Selector_2 s261_7(wires_65_6[1], addr_65_6, addr_positional[1047:1044], addr_261_7);

wire[31:0] addr_262_7;

Selector_2 s262_7(wires_65_6[2], addr_65_6, addr_positional[1051:1048], addr_262_7);

wire[31:0] addr_263_7;

Selector_2 s263_7(wires_65_6[3], addr_65_6, addr_positional[1055:1052], addr_263_7);

wire[31:0] addr_264_7;

Selector_2 s264_7(wires_66_6[0], addr_66_6, addr_positional[1059:1056], addr_264_7);

wire[31:0] addr_265_7;

Selector_2 s265_7(wires_66_6[1], addr_66_6, addr_positional[1063:1060], addr_265_7);

wire[31:0] addr_266_7;

Selector_2 s266_7(wires_66_6[2], addr_66_6, addr_positional[1067:1064], addr_266_7);

wire[31:0] addr_267_7;

Selector_2 s267_7(wires_66_6[3], addr_66_6, addr_positional[1071:1068], addr_267_7);

wire[31:0] addr_268_7;

Selector_2 s268_7(wires_67_6[0], addr_67_6, addr_positional[1075:1072], addr_268_7);

wire[31:0] addr_269_7;

Selector_2 s269_7(wires_67_6[1], addr_67_6, addr_positional[1079:1076], addr_269_7);

wire[31:0] addr_270_7;

Selector_2 s270_7(wires_67_6[2], addr_67_6, addr_positional[1083:1080], addr_270_7);

wire[31:0] addr_271_7;

Selector_2 s271_7(wires_67_6[3], addr_67_6, addr_positional[1087:1084], addr_271_7);

wire[31:0] addr_272_7;

Selector_2 s272_7(wires_68_6[0], addr_68_6, addr_positional[1091:1088], addr_272_7);

wire[31:0] addr_273_7;

Selector_2 s273_7(wires_68_6[1], addr_68_6, addr_positional[1095:1092], addr_273_7);

wire[31:0] addr_274_7;

Selector_2 s274_7(wires_68_6[2], addr_68_6, addr_positional[1099:1096], addr_274_7);

wire[31:0] addr_275_7;

Selector_2 s275_7(wires_68_6[3], addr_68_6, addr_positional[1103:1100], addr_275_7);

wire[31:0] addr_276_7;

Selector_2 s276_7(wires_69_6[0], addr_69_6, addr_positional[1107:1104], addr_276_7);

wire[31:0] addr_277_7;

Selector_2 s277_7(wires_69_6[1], addr_69_6, addr_positional[1111:1108], addr_277_7);

wire[31:0] addr_278_7;

Selector_2 s278_7(wires_69_6[2], addr_69_6, addr_positional[1115:1112], addr_278_7);

wire[31:0] addr_279_7;

Selector_2 s279_7(wires_69_6[3], addr_69_6, addr_positional[1119:1116], addr_279_7);

wire[31:0] addr_280_7;

Selector_2 s280_7(wires_70_6[0], addr_70_6, addr_positional[1123:1120], addr_280_7);

wire[31:0] addr_281_7;

Selector_2 s281_7(wires_70_6[1], addr_70_6, addr_positional[1127:1124], addr_281_7);

wire[31:0] addr_282_7;

Selector_2 s282_7(wires_70_6[2], addr_70_6, addr_positional[1131:1128], addr_282_7);

wire[31:0] addr_283_7;

Selector_2 s283_7(wires_70_6[3], addr_70_6, addr_positional[1135:1132], addr_283_7);

wire[31:0] addr_284_7;

Selector_2 s284_7(wires_71_6[0], addr_71_6, addr_positional[1139:1136], addr_284_7);

wire[31:0] addr_285_7;

Selector_2 s285_7(wires_71_6[1], addr_71_6, addr_positional[1143:1140], addr_285_7);

wire[31:0] addr_286_7;

Selector_2 s286_7(wires_71_6[2], addr_71_6, addr_positional[1147:1144], addr_286_7);

wire[31:0] addr_287_7;

Selector_2 s287_7(wires_71_6[3], addr_71_6, addr_positional[1151:1148], addr_287_7);

wire[31:0] addr_288_7;

Selector_2 s288_7(wires_72_6[0], addr_72_6, addr_positional[1155:1152], addr_288_7);

wire[31:0] addr_289_7;

Selector_2 s289_7(wires_72_6[1], addr_72_6, addr_positional[1159:1156], addr_289_7);

wire[31:0] addr_290_7;

Selector_2 s290_7(wires_72_6[2], addr_72_6, addr_positional[1163:1160], addr_290_7);

wire[31:0] addr_291_7;

Selector_2 s291_7(wires_72_6[3], addr_72_6, addr_positional[1167:1164], addr_291_7);

wire[31:0] addr_292_7;

Selector_2 s292_7(wires_73_6[0], addr_73_6, addr_positional[1171:1168], addr_292_7);

wire[31:0] addr_293_7;

Selector_2 s293_7(wires_73_6[1], addr_73_6, addr_positional[1175:1172], addr_293_7);

wire[31:0] addr_294_7;

Selector_2 s294_7(wires_73_6[2], addr_73_6, addr_positional[1179:1176], addr_294_7);

wire[31:0] addr_295_7;

Selector_2 s295_7(wires_73_6[3], addr_73_6, addr_positional[1183:1180], addr_295_7);

wire[31:0] addr_296_7;

Selector_2 s296_7(wires_74_6[0], addr_74_6, addr_positional[1187:1184], addr_296_7);

wire[31:0] addr_297_7;

Selector_2 s297_7(wires_74_6[1], addr_74_6, addr_positional[1191:1188], addr_297_7);

wire[31:0] addr_298_7;

Selector_2 s298_7(wires_74_6[2], addr_74_6, addr_positional[1195:1192], addr_298_7);

wire[31:0] addr_299_7;

Selector_2 s299_7(wires_74_6[3], addr_74_6, addr_positional[1199:1196], addr_299_7);

wire[31:0] addr_300_7;

Selector_2 s300_7(wires_75_6[0], addr_75_6, addr_positional[1203:1200], addr_300_7);

wire[31:0] addr_301_7;

Selector_2 s301_7(wires_75_6[1], addr_75_6, addr_positional[1207:1204], addr_301_7);

wire[31:0] addr_302_7;

Selector_2 s302_7(wires_75_6[2], addr_75_6, addr_positional[1211:1208], addr_302_7);

wire[31:0] addr_303_7;

Selector_2 s303_7(wires_75_6[3], addr_75_6, addr_positional[1215:1212], addr_303_7);

wire[31:0] addr_304_7;

Selector_2 s304_7(wires_76_6[0], addr_76_6, addr_positional[1219:1216], addr_304_7);

wire[31:0] addr_305_7;

Selector_2 s305_7(wires_76_6[1], addr_76_6, addr_positional[1223:1220], addr_305_7);

wire[31:0] addr_306_7;

Selector_2 s306_7(wires_76_6[2], addr_76_6, addr_positional[1227:1224], addr_306_7);

wire[31:0] addr_307_7;

Selector_2 s307_7(wires_76_6[3], addr_76_6, addr_positional[1231:1228], addr_307_7);

wire[31:0] addr_308_7;

Selector_2 s308_7(wires_77_6[0], addr_77_6, addr_positional[1235:1232], addr_308_7);

wire[31:0] addr_309_7;

Selector_2 s309_7(wires_77_6[1], addr_77_6, addr_positional[1239:1236], addr_309_7);

wire[31:0] addr_310_7;

Selector_2 s310_7(wires_77_6[2], addr_77_6, addr_positional[1243:1240], addr_310_7);

wire[31:0] addr_311_7;

Selector_2 s311_7(wires_77_6[3], addr_77_6, addr_positional[1247:1244], addr_311_7);

wire[31:0] addr_312_7;

Selector_2 s312_7(wires_78_6[0], addr_78_6, addr_positional[1251:1248], addr_312_7);

wire[31:0] addr_313_7;

Selector_2 s313_7(wires_78_6[1], addr_78_6, addr_positional[1255:1252], addr_313_7);

wire[31:0] addr_314_7;

Selector_2 s314_7(wires_78_6[2], addr_78_6, addr_positional[1259:1256], addr_314_7);

wire[31:0] addr_315_7;

Selector_2 s315_7(wires_78_6[3], addr_78_6, addr_positional[1263:1260], addr_315_7);

wire[31:0] addr_316_7;

Selector_2 s316_7(wires_79_6[0], addr_79_6, addr_positional[1267:1264], addr_316_7);

wire[31:0] addr_317_7;

Selector_2 s317_7(wires_79_6[1], addr_79_6, addr_positional[1271:1268], addr_317_7);

wire[31:0] addr_318_7;

Selector_2 s318_7(wires_79_6[2], addr_79_6, addr_positional[1275:1272], addr_318_7);

wire[31:0] addr_319_7;

Selector_2 s319_7(wires_79_6[3], addr_79_6, addr_positional[1279:1276], addr_319_7);

wire[31:0] addr_320_7;

Selector_2 s320_7(wires_80_6[0], addr_80_6, addr_positional[1283:1280], addr_320_7);

wire[31:0] addr_321_7;

Selector_2 s321_7(wires_80_6[1], addr_80_6, addr_positional[1287:1284], addr_321_7);

wire[31:0] addr_322_7;

Selector_2 s322_7(wires_80_6[2], addr_80_6, addr_positional[1291:1288], addr_322_7);

wire[31:0] addr_323_7;

Selector_2 s323_7(wires_80_6[3], addr_80_6, addr_positional[1295:1292], addr_323_7);

wire[31:0] addr_324_7;

Selector_2 s324_7(wires_81_6[0], addr_81_6, addr_positional[1299:1296], addr_324_7);

wire[31:0] addr_325_7;

Selector_2 s325_7(wires_81_6[1], addr_81_6, addr_positional[1303:1300], addr_325_7);

wire[31:0] addr_326_7;

Selector_2 s326_7(wires_81_6[2], addr_81_6, addr_positional[1307:1304], addr_326_7);

wire[31:0] addr_327_7;

Selector_2 s327_7(wires_81_6[3], addr_81_6, addr_positional[1311:1308], addr_327_7);

wire[31:0] addr_328_7;

Selector_2 s328_7(wires_82_6[0], addr_82_6, addr_positional[1315:1312], addr_328_7);

wire[31:0] addr_329_7;

Selector_2 s329_7(wires_82_6[1], addr_82_6, addr_positional[1319:1316], addr_329_7);

wire[31:0] addr_330_7;

Selector_2 s330_7(wires_82_6[2], addr_82_6, addr_positional[1323:1320], addr_330_7);

wire[31:0] addr_331_7;

Selector_2 s331_7(wires_82_6[3], addr_82_6, addr_positional[1327:1324], addr_331_7);

wire[31:0] addr_332_7;

Selector_2 s332_7(wires_83_6[0], addr_83_6, addr_positional[1331:1328], addr_332_7);

wire[31:0] addr_333_7;

Selector_2 s333_7(wires_83_6[1], addr_83_6, addr_positional[1335:1332], addr_333_7);

wire[31:0] addr_334_7;

Selector_2 s334_7(wires_83_6[2], addr_83_6, addr_positional[1339:1336], addr_334_7);

wire[31:0] addr_335_7;

Selector_2 s335_7(wires_83_6[3], addr_83_6, addr_positional[1343:1340], addr_335_7);

wire[31:0] addr_336_7;

Selector_2 s336_7(wires_84_6[0], addr_84_6, addr_positional[1347:1344], addr_336_7);

wire[31:0] addr_337_7;

Selector_2 s337_7(wires_84_6[1], addr_84_6, addr_positional[1351:1348], addr_337_7);

wire[31:0] addr_338_7;

Selector_2 s338_7(wires_84_6[2], addr_84_6, addr_positional[1355:1352], addr_338_7);

wire[31:0] addr_339_7;

Selector_2 s339_7(wires_84_6[3], addr_84_6, addr_positional[1359:1356], addr_339_7);

wire[31:0] addr_340_7;

Selector_2 s340_7(wires_85_6[0], addr_85_6, addr_positional[1363:1360], addr_340_7);

wire[31:0] addr_341_7;

Selector_2 s341_7(wires_85_6[1], addr_85_6, addr_positional[1367:1364], addr_341_7);

wire[31:0] addr_342_7;

Selector_2 s342_7(wires_85_6[2], addr_85_6, addr_positional[1371:1368], addr_342_7);

wire[31:0] addr_343_7;

Selector_2 s343_7(wires_85_6[3], addr_85_6, addr_positional[1375:1372], addr_343_7);

wire[31:0] addr_344_7;

Selector_2 s344_7(wires_86_6[0], addr_86_6, addr_positional[1379:1376], addr_344_7);

wire[31:0] addr_345_7;

Selector_2 s345_7(wires_86_6[1], addr_86_6, addr_positional[1383:1380], addr_345_7);

wire[31:0] addr_346_7;

Selector_2 s346_7(wires_86_6[2], addr_86_6, addr_positional[1387:1384], addr_346_7);

wire[31:0] addr_347_7;

Selector_2 s347_7(wires_86_6[3], addr_86_6, addr_positional[1391:1388], addr_347_7);

wire[31:0] addr_348_7;

Selector_2 s348_7(wires_87_6[0], addr_87_6, addr_positional[1395:1392], addr_348_7);

wire[31:0] addr_349_7;

Selector_2 s349_7(wires_87_6[1], addr_87_6, addr_positional[1399:1396], addr_349_7);

wire[31:0] addr_350_7;

Selector_2 s350_7(wires_87_6[2], addr_87_6, addr_positional[1403:1400], addr_350_7);

wire[31:0] addr_351_7;

Selector_2 s351_7(wires_87_6[3], addr_87_6, addr_positional[1407:1404], addr_351_7);

wire[31:0] addr_352_7;

Selector_2 s352_7(wires_88_6[0], addr_88_6, addr_positional[1411:1408], addr_352_7);

wire[31:0] addr_353_7;

Selector_2 s353_7(wires_88_6[1], addr_88_6, addr_positional[1415:1412], addr_353_7);

wire[31:0] addr_354_7;

Selector_2 s354_7(wires_88_6[2], addr_88_6, addr_positional[1419:1416], addr_354_7);

wire[31:0] addr_355_7;

Selector_2 s355_7(wires_88_6[3], addr_88_6, addr_positional[1423:1420], addr_355_7);

wire[31:0] addr_356_7;

Selector_2 s356_7(wires_89_6[0], addr_89_6, addr_positional[1427:1424], addr_356_7);

wire[31:0] addr_357_7;

Selector_2 s357_7(wires_89_6[1], addr_89_6, addr_positional[1431:1428], addr_357_7);

wire[31:0] addr_358_7;

Selector_2 s358_7(wires_89_6[2], addr_89_6, addr_positional[1435:1432], addr_358_7);

wire[31:0] addr_359_7;

Selector_2 s359_7(wires_89_6[3], addr_89_6, addr_positional[1439:1436], addr_359_7);

wire[31:0] addr_360_7;

Selector_2 s360_7(wires_90_6[0], addr_90_6, addr_positional[1443:1440], addr_360_7);

wire[31:0] addr_361_7;

Selector_2 s361_7(wires_90_6[1], addr_90_6, addr_positional[1447:1444], addr_361_7);

wire[31:0] addr_362_7;

Selector_2 s362_7(wires_90_6[2], addr_90_6, addr_positional[1451:1448], addr_362_7);

wire[31:0] addr_363_7;

Selector_2 s363_7(wires_90_6[3], addr_90_6, addr_positional[1455:1452], addr_363_7);

wire[31:0] addr_364_7;

Selector_2 s364_7(wires_91_6[0], addr_91_6, addr_positional[1459:1456], addr_364_7);

wire[31:0] addr_365_7;

Selector_2 s365_7(wires_91_6[1], addr_91_6, addr_positional[1463:1460], addr_365_7);

wire[31:0] addr_366_7;

Selector_2 s366_7(wires_91_6[2], addr_91_6, addr_positional[1467:1464], addr_366_7);

wire[31:0] addr_367_7;

Selector_2 s367_7(wires_91_6[3], addr_91_6, addr_positional[1471:1468], addr_367_7);

wire[31:0] addr_368_7;

Selector_2 s368_7(wires_92_6[0], addr_92_6, addr_positional[1475:1472], addr_368_7);

wire[31:0] addr_369_7;

Selector_2 s369_7(wires_92_6[1], addr_92_6, addr_positional[1479:1476], addr_369_7);

wire[31:0] addr_370_7;

Selector_2 s370_7(wires_92_6[2], addr_92_6, addr_positional[1483:1480], addr_370_7);

wire[31:0] addr_371_7;

Selector_2 s371_7(wires_92_6[3], addr_92_6, addr_positional[1487:1484], addr_371_7);

wire[31:0] addr_372_7;

Selector_2 s372_7(wires_93_6[0], addr_93_6, addr_positional[1491:1488], addr_372_7);

wire[31:0] addr_373_7;

Selector_2 s373_7(wires_93_6[1], addr_93_6, addr_positional[1495:1492], addr_373_7);

wire[31:0] addr_374_7;

Selector_2 s374_7(wires_93_6[2], addr_93_6, addr_positional[1499:1496], addr_374_7);

wire[31:0] addr_375_7;

Selector_2 s375_7(wires_93_6[3], addr_93_6, addr_positional[1503:1500], addr_375_7);

wire[31:0] addr_376_7;

Selector_2 s376_7(wires_94_6[0], addr_94_6, addr_positional[1507:1504], addr_376_7);

wire[31:0] addr_377_7;

Selector_2 s377_7(wires_94_6[1], addr_94_6, addr_positional[1511:1508], addr_377_7);

wire[31:0] addr_378_7;

Selector_2 s378_7(wires_94_6[2], addr_94_6, addr_positional[1515:1512], addr_378_7);

wire[31:0] addr_379_7;

Selector_2 s379_7(wires_94_6[3], addr_94_6, addr_positional[1519:1516], addr_379_7);

wire[31:0] addr_380_7;

Selector_2 s380_7(wires_95_6[0], addr_95_6, addr_positional[1523:1520], addr_380_7);

wire[31:0] addr_381_7;

Selector_2 s381_7(wires_95_6[1], addr_95_6, addr_positional[1527:1524], addr_381_7);

wire[31:0] addr_382_7;

Selector_2 s382_7(wires_95_6[2], addr_95_6, addr_positional[1531:1528], addr_382_7);

wire[31:0] addr_383_7;

Selector_2 s383_7(wires_95_6[3], addr_95_6, addr_positional[1535:1532], addr_383_7);

wire[31:0] addr_384_7;

Selector_2 s384_7(wires_96_6[0], addr_96_6, addr_positional[1539:1536], addr_384_7);

wire[31:0] addr_385_7;

Selector_2 s385_7(wires_96_6[1], addr_96_6, addr_positional[1543:1540], addr_385_7);

wire[31:0] addr_386_7;

Selector_2 s386_7(wires_96_6[2], addr_96_6, addr_positional[1547:1544], addr_386_7);

wire[31:0] addr_387_7;

Selector_2 s387_7(wires_96_6[3], addr_96_6, addr_positional[1551:1548], addr_387_7);

wire[31:0] addr_388_7;

Selector_2 s388_7(wires_97_6[0], addr_97_6, addr_positional[1555:1552], addr_388_7);

wire[31:0] addr_389_7;

Selector_2 s389_7(wires_97_6[1], addr_97_6, addr_positional[1559:1556], addr_389_7);

wire[31:0] addr_390_7;

Selector_2 s390_7(wires_97_6[2], addr_97_6, addr_positional[1563:1560], addr_390_7);

wire[31:0] addr_391_7;

Selector_2 s391_7(wires_97_6[3], addr_97_6, addr_positional[1567:1564], addr_391_7);

wire[31:0] addr_392_7;

Selector_2 s392_7(wires_98_6[0], addr_98_6, addr_positional[1571:1568], addr_392_7);

wire[31:0] addr_393_7;

Selector_2 s393_7(wires_98_6[1], addr_98_6, addr_positional[1575:1572], addr_393_7);

wire[31:0] addr_394_7;

Selector_2 s394_7(wires_98_6[2], addr_98_6, addr_positional[1579:1576], addr_394_7);

wire[31:0] addr_395_7;

Selector_2 s395_7(wires_98_6[3], addr_98_6, addr_positional[1583:1580], addr_395_7);

wire[31:0] addr_396_7;

Selector_2 s396_7(wires_99_6[0], addr_99_6, addr_positional[1587:1584], addr_396_7);

wire[31:0] addr_397_7;

Selector_2 s397_7(wires_99_6[1], addr_99_6, addr_positional[1591:1588], addr_397_7);

wire[31:0] addr_398_7;

Selector_2 s398_7(wires_99_6[2], addr_99_6, addr_positional[1595:1592], addr_398_7);

wire[31:0] addr_399_7;

Selector_2 s399_7(wires_99_6[3], addr_99_6, addr_positional[1599:1596], addr_399_7);

wire[31:0] addr_400_7;

Selector_2 s400_7(wires_100_6[0], addr_100_6, addr_positional[1603:1600], addr_400_7);

wire[31:0] addr_401_7;

Selector_2 s401_7(wires_100_6[1], addr_100_6, addr_positional[1607:1604], addr_401_7);

wire[31:0] addr_402_7;

Selector_2 s402_7(wires_100_6[2], addr_100_6, addr_positional[1611:1608], addr_402_7);

wire[31:0] addr_403_7;

Selector_2 s403_7(wires_100_6[3], addr_100_6, addr_positional[1615:1612], addr_403_7);

wire[31:0] addr_404_7;

Selector_2 s404_7(wires_101_6[0], addr_101_6, addr_positional[1619:1616], addr_404_7);

wire[31:0] addr_405_7;

Selector_2 s405_7(wires_101_6[1], addr_101_6, addr_positional[1623:1620], addr_405_7);

wire[31:0] addr_406_7;

Selector_2 s406_7(wires_101_6[2], addr_101_6, addr_positional[1627:1624], addr_406_7);

wire[31:0] addr_407_7;

Selector_2 s407_7(wires_101_6[3], addr_101_6, addr_positional[1631:1628], addr_407_7);

wire[31:0] addr_408_7;

Selector_2 s408_7(wires_102_6[0], addr_102_6, addr_positional[1635:1632], addr_408_7);

wire[31:0] addr_409_7;

Selector_2 s409_7(wires_102_6[1], addr_102_6, addr_positional[1639:1636], addr_409_7);

wire[31:0] addr_410_7;

Selector_2 s410_7(wires_102_6[2], addr_102_6, addr_positional[1643:1640], addr_410_7);

wire[31:0] addr_411_7;

Selector_2 s411_7(wires_102_6[3], addr_102_6, addr_positional[1647:1644], addr_411_7);

wire[31:0] addr_412_7;

Selector_2 s412_7(wires_103_6[0], addr_103_6, addr_positional[1651:1648], addr_412_7);

wire[31:0] addr_413_7;

Selector_2 s413_7(wires_103_6[1], addr_103_6, addr_positional[1655:1652], addr_413_7);

wire[31:0] addr_414_7;

Selector_2 s414_7(wires_103_6[2], addr_103_6, addr_positional[1659:1656], addr_414_7);

wire[31:0] addr_415_7;

Selector_2 s415_7(wires_103_6[3], addr_103_6, addr_positional[1663:1660], addr_415_7);

wire[31:0] addr_416_7;

Selector_2 s416_7(wires_104_6[0], addr_104_6, addr_positional[1667:1664], addr_416_7);

wire[31:0] addr_417_7;

Selector_2 s417_7(wires_104_6[1], addr_104_6, addr_positional[1671:1668], addr_417_7);

wire[31:0] addr_418_7;

Selector_2 s418_7(wires_104_6[2], addr_104_6, addr_positional[1675:1672], addr_418_7);

wire[31:0] addr_419_7;

Selector_2 s419_7(wires_104_6[3], addr_104_6, addr_positional[1679:1676], addr_419_7);

wire[31:0] addr_420_7;

Selector_2 s420_7(wires_105_6[0], addr_105_6, addr_positional[1683:1680], addr_420_7);

wire[31:0] addr_421_7;

Selector_2 s421_7(wires_105_6[1], addr_105_6, addr_positional[1687:1684], addr_421_7);

wire[31:0] addr_422_7;

Selector_2 s422_7(wires_105_6[2], addr_105_6, addr_positional[1691:1688], addr_422_7);

wire[31:0] addr_423_7;

Selector_2 s423_7(wires_105_6[3], addr_105_6, addr_positional[1695:1692], addr_423_7);

wire[31:0] addr_424_7;

Selector_2 s424_7(wires_106_6[0], addr_106_6, addr_positional[1699:1696], addr_424_7);

wire[31:0] addr_425_7;

Selector_2 s425_7(wires_106_6[1], addr_106_6, addr_positional[1703:1700], addr_425_7);

wire[31:0] addr_426_7;

Selector_2 s426_7(wires_106_6[2], addr_106_6, addr_positional[1707:1704], addr_426_7);

wire[31:0] addr_427_7;

Selector_2 s427_7(wires_106_6[3], addr_106_6, addr_positional[1711:1708], addr_427_7);

wire[31:0] addr_428_7;

Selector_2 s428_7(wires_107_6[0], addr_107_6, addr_positional[1715:1712], addr_428_7);

wire[31:0] addr_429_7;

Selector_2 s429_7(wires_107_6[1], addr_107_6, addr_positional[1719:1716], addr_429_7);

wire[31:0] addr_430_7;

Selector_2 s430_7(wires_107_6[2], addr_107_6, addr_positional[1723:1720], addr_430_7);

wire[31:0] addr_431_7;

Selector_2 s431_7(wires_107_6[3], addr_107_6, addr_positional[1727:1724], addr_431_7);

wire[31:0] addr_432_7;

Selector_2 s432_7(wires_108_6[0], addr_108_6, addr_positional[1731:1728], addr_432_7);

wire[31:0] addr_433_7;

Selector_2 s433_7(wires_108_6[1], addr_108_6, addr_positional[1735:1732], addr_433_7);

wire[31:0] addr_434_7;

Selector_2 s434_7(wires_108_6[2], addr_108_6, addr_positional[1739:1736], addr_434_7);

wire[31:0] addr_435_7;

Selector_2 s435_7(wires_108_6[3], addr_108_6, addr_positional[1743:1740], addr_435_7);

wire[31:0] addr_436_7;

Selector_2 s436_7(wires_109_6[0], addr_109_6, addr_positional[1747:1744], addr_436_7);

wire[31:0] addr_437_7;

Selector_2 s437_7(wires_109_6[1], addr_109_6, addr_positional[1751:1748], addr_437_7);

wire[31:0] addr_438_7;

Selector_2 s438_7(wires_109_6[2], addr_109_6, addr_positional[1755:1752], addr_438_7);

wire[31:0] addr_439_7;

Selector_2 s439_7(wires_109_6[3], addr_109_6, addr_positional[1759:1756], addr_439_7);

wire[31:0] addr_440_7;

Selector_2 s440_7(wires_110_6[0], addr_110_6, addr_positional[1763:1760], addr_440_7);

wire[31:0] addr_441_7;

Selector_2 s441_7(wires_110_6[1], addr_110_6, addr_positional[1767:1764], addr_441_7);

wire[31:0] addr_442_7;

Selector_2 s442_7(wires_110_6[2], addr_110_6, addr_positional[1771:1768], addr_442_7);

wire[31:0] addr_443_7;

Selector_2 s443_7(wires_110_6[3], addr_110_6, addr_positional[1775:1772], addr_443_7);

wire[31:0] addr_444_7;

Selector_2 s444_7(wires_111_6[0], addr_111_6, addr_positional[1779:1776], addr_444_7);

wire[31:0] addr_445_7;

Selector_2 s445_7(wires_111_6[1], addr_111_6, addr_positional[1783:1780], addr_445_7);

wire[31:0] addr_446_7;

Selector_2 s446_7(wires_111_6[2], addr_111_6, addr_positional[1787:1784], addr_446_7);

wire[31:0] addr_447_7;

Selector_2 s447_7(wires_111_6[3], addr_111_6, addr_positional[1791:1788], addr_447_7);

wire[31:0] addr_448_7;

Selector_2 s448_7(wires_112_6[0], addr_112_6, addr_positional[1795:1792], addr_448_7);

wire[31:0] addr_449_7;

Selector_2 s449_7(wires_112_6[1], addr_112_6, addr_positional[1799:1796], addr_449_7);

wire[31:0] addr_450_7;

Selector_2 s450_7(wires_112_6[2], addr_112_6, addr_positional[1803:1800], addr_450_7);

wire[31:0] addr_451_7;

Selector_2 s451_7(wires_112_6[3], addr_112_6, addr_positional[1807:1804], addr_451_7);

wire[31:0] addr_452_7;

Selector_2 s452_7(wires_113_6[0], addr_113_6, addr_positional[1811:1808], addr_452_7);

wire[31:0] addr_453_7;

Selector_2 s453_7(wires_113_6[1], addr_113_6, addr_positional[1815:1812], addr_453_7);

wire[31:0] addr_454_7;

Selector_2 s454_7(wires_113_6[2], addr_113_6, addr_positional[1819:1816], addr_454_7);

wire[31:0] addr_455_7;

Selector_2 s455_7(wires_113_6[3], addr_113_6, addr_positional[1823:1820], addr_455_7);

wire[31:0] addr_456_7;

Selector_2 s456_7(wires_114_6[0], addr_114_6, addr_positional[1827:1824], addr_456_7);

wire[31:0] addr_457_7;

Selector_2 s457_7(wires_114_6[1], addr_114_6, addr_positional[1831:1828], addr_457_7);

wire[31:0] addr_458_7;

Selector_2 s458_7(wires_114_6[2], addr_114_6, addr_positional[1835:1832], addr_458_7);

wire[31:0] addr_459_7;

Selector_2 s459_7(wires_114_6[3], addr_114_6, addr_positional[1839:1836], addr_459_7);

wire[31:0] addr_460_7;

Selector_2 s460_7(wires_115_6[0], addr_115_6, addr_positional[1843:1840], addr_460_7);

wire[31:0] addr_461_7;

Selector_2 s461_7(wires_115_6[1], addr_115_6, addr_positional[1847:1844], addr_461_7);

wire[31:0] addr_462_7;

Selector_2 s462_7(wires_115_6[2], addr_115_6, addr_positional[1851:1848], addr_462_7);

wire[31:0] addr_463_7;

Selector_2 s463_7(wires_115_6[3], addr_115_6, addr_positional[1855:1852], addr_463_7);

wire[31:0] addr_464_7;

Selector_2 s464_7(wires_116_6[0], addr_116_6, addr_positional[1859:1856], addr_464_7);

wire[31:0] addr_465_7;

Selector_2 s465_7(wires_116_6[1], addr_116_6, addr_positional[1863:1860], addr_465_7);

wire[31:0] addr_466_7;

Selector_2 s466_7(wires_116_6[2], addr_116_6, addr_positional[1867:1864], addr_466_7);

wire[31:0] addr_467_7;

Selector_2 s467_7(wires_116_6[3], addr_116_6, addr_positional[1871:1868], addr_467_7);

wire[31:0] addr_468_7;

Selector_2 s468_7(wires_117_6[0], addr_117_6, addr_positional[1875:1872], addr_468_7);

wire[31:0] addr_469_7;

Selector_2 s469_7(wires_117_6[1], addr_117_6, addr_positional[1879:1876], addr_469_7);

wire[31:0] addr_470_7;

Selector_2 s470_7(wires_117_6[2], addr_117_6, addr_positional[1883:1880], addr_470_7);

wire[31:0] addr_471_7;

Selector_2 s471_7(wires_117_6[3], addr_117_6, addr_positional[1887:1884], addr_471_7);

wire[31:0] addr_472_7;

Selector_2 s472_7(wires_118_6[0], addr_118_6, addr_positional[1891:1888], addr_472_7);

wire[31:0] addr_473_7;

Selector_2 s473_7(wires_118_6[1], addr_118_6, addr_positional[1895:1892], addr_473_7);

wire[31:0] addr_474_7;

Selector_2 s474_7(wires_118_6[2], addr_118_6, addr_positional[1899:1896], addr_474_7);

wire[31:0] addr_475_7;

Selector_2 s475_7(wires_118_6[3], addr_118_6, addr_positional[1903:1900], addr_475_7);

wire[31:0] addr_476_7;

Selector_2 s476_7(wires_119_6[0], addr_119_6, addr_positional[1907:1904], addr_476_7);

wire[31:0] addr_477_7;

Selector_2 s477_7(wires_119_6[1], addr_119_6, addr_positional[1911:1908], addr_477_7);

wire[31:0] addr_478_7;

Selector_2 s478_7(wires_119_6[2], addr_119_6, addr_positional[1915:1912], addr_478_7);

wire[31:0] addr_479_7;

Selector_2 s479_7(wires_119_6[3], addr_119_6, addr_positional[1919:1916], addr_479_7);

wire[31:0] addr_480_7;

Selector_2 s480_7(wires_120_6[0], addr_120_6, addr_positional[1923:1920], addr_480_7);

wire[31:0] addr_481_7;

Selector_2 s481_7(wires_120_6[1], addr_120_6, addr_positional[1927:1924], addr_481_7);

wire[31:0] addr_482_7;

Selector_2 s482_7(wires_120_6[2], addr_120_6, addr_positional[1931:1928], addr_482_7);

wire[31:0] addr_483_7;

Selector_2 s483_7(wires_120_6[3], addr_120_6, addr_positional[1935:1932], addr_483_7);

wire[31:0] addr_484_7;

Selector_2 s484_7(wires_121_6[0], addr_121_6, addr_positional[1939:1936], addr_484_7);

wire[31:0] addr_485_7;

Selector_2 s485_7(wires_121_6[1], addr_121_6, addr_positional[1943:1940], addr_485_7);

wire[31:0] addr_486_7;

Selector_2 s486_7(wires_121_6[2], addr_121_6, addr_positional[1947:1944], addr_486_7);

wire[31:0] addr_487_7;

Selector_2 s487_7(wires_121_6[3], addr_121_6, addr_positional[1951:1948], addr_487_7);

wire[31:0] addr_488_7;

Selector_2 s488_7(wires_122_6[0], addr_122_6, addr_positional[1955:1952], addr_488_7);

wire[31:0] addr_489_7;

Selector_2 s489_7(wires_122_6[1], addr_122_6, addr_positional[1959:1956], addr_489_7);

wire[31:0] addr_490_7;

Selector_2 s490_7(wires_122_6[2], addr_122_6, addr_positional[1963:1960], addr_490_7);

wire[31:0] addr_491_7;

Selector_2 s491_7(wires_122_6[3], addr_122_6, addr_positional[1967:1964], addr_491_7);

wire[31:0] addr_492_7;

Selector_2 s492_7(wires_123_6[0], addr_123_6, addr_positional[1971:1968], addr_492_7);

wire[31:0] addr_493_7;

Selector_2 s493_7(wires_123_6[1], addr_123_6, addr_positional[1975:1972], addr_493_7);

wire[31:0] addr_494_7;

Selector_2 s494_7(wires_123_6[2], addr_123_6, addr_positional[1979:1976], addr_494_7);

wire[31:0] addr_495_7;

Selector_2 s495_7(wires_123_6[3], addr_123_6, addr_positional[1983:1980], addr_495_7);

wire[31:0] addr_496_7;

Selector_2 s496_7(wires_124_6[0], addr_124_6, addr_positional[1987:1984], addr_496_7);

wire[31:0] addr_497_7;

Selector_2 s497_7(wires_124_6[1], addr_124_6, addr_positional[1991:1988], addr_497_7);

wire[31:0] addr_498_7;

Selector_2 s498_7(wires_124_6[2], addr_124_6, addr_positional[1995:1992], addr_498_7);

wire[31:0] addr_499_7;

Selector_2 s499_7(wires_124_6[3], addr_124_6, addr_positional[1999:1996], addr_499_7);

wire[31:0] addr_500_7;

Selector_2 s500_7(wires_125_6[0], addr_125_6, addr_positional[2003:2000], addr_500_7);

wire[31:0] addr_501_7;

Selector_2 s501_7(wires_125_6[1], addr_125_6, addr_positional[2007:2004], addr_501_7);

wire[31:0] addr_502_7;

Selector_2 s502_7(wires_125_6[2], addr_125_6, addr_positional[2011:2008], addr_502_7);

wire[31:0] addr_503_7;

Selector_2 s503_7(wires_125_6[3], addr_125_6, addr_positional[2015:2012], addr_503_7);

wire[31:0] addr_504_7;

Selector_2 s504_7(wires_126_6[0], addr_126_6, addr_positional[2019:2016], addr_504_7);

wire[31:0] addr_505_7;

Selector_2 s505_7(wires_126_6[1], addr_126_6, addr_positional[2023:2020], addr_505_7);

wire[31:0] addr_506_7;

Selector_2 s506_7(wires_126_6[2], addr_126_6, addr_positional[2027:2024], addr_506_7);

wire[31:0] addr_507_7;

Selector_2 s507_7(wires_126_6[3], addr_126_6, addr_positional[2031:2028], addr_507_7);

wire[31:0] addr_508_7;

Selector_2 s508_7(wires_127_6[0], addr_127_6, addr_positional[2035:2032], addr_508_7);

wire[31:0] addr_509_7;

Selector_2 s509_7(wires_127_6[1], addr_127_6, addr_positional[2039:2036], addr_509_7);

wire[31:0] addr_510_7;

Selector_2 s510_7(wires_127_6[2], addr_127_6, addr_positional[2043:2040], addr_510_7);

wire[31:0] addr_511_7;

Selector_2 s511_7(wires_127_6[3], addr_127_6, addr_positional[2047:2044], addr_511_7);

wire[31:0] addr_512_7;

Selector_2 s512_7(wires_128_6[0], addr_128_6, addr_positional[2051:2048], addr_512_7);

wire[31:0] addr_513_7;

Selector_2 s513_7(wires_128_6[1], addr_128_6, addr_positional[2055:2052], addr_513_7);

wire[31:0] addr_514_7;

Selector_2 s514_7(wires_128_6[2], addr_128_6, addr_positional[2059:2056], addr_514_7);

wire[31:0] addr_515_7;

Selector_2 s515_7(wires_128_6[3], addr_128_6, addr_positional[2063:2060], addr_515_7);

wire[31:0] addr_516_7;

Selector_2 s516_7(wires_129_6[0], addr_129_6, addr_positional[2067:2064], addr_516_7);

wire[31:0] addr_517_7;

Selector_2 s517_7(wires_129_6[1], addr_129_6, addr_positional[2071:2068], addr_517_7);

wire[31:0] addr_518_7;

Selector_2 s518_7(wires_129_6[2], addr_129_6, addr_positional[2075:2072], addr_518_7);

wire[31:0] addr_519_7;

Selector_2 s519_7(wires_129_6[3], addr_129_6, addr_positional[2079:2076], addr_519_7);

wire[31:0] addr_520_7;

Selector_2 s520_7(wires_130_6[0], addr_130_6, addr_positional[2083:2080], addr_520_7);

wire[31:0] addr_521_7;

Selector_2 s521_7(wires_130_6[1], addr_130_6, addr_positional[2087:2084], addr_521_7);

wire[31:0] addr_522_7;

Selector_2 s522_7(wires_130_6[2], addr_130_6, addr_positional[2091:2088], addr_522_7);

wire[31:0] addr_523_7;

Selector_2 s523_7(wires_130_6[3], addr_130_6, addr_positional[2095:2092], addr_523_7);

wire[31:0] addr_524_7;

Selector_2 s524_7(wires_131_6[0], addr_131_6, addr_positional[2099:2096], addr_524_7);

wire[31:0] addr_525_7;

Selector_2 s525_7(wires_131_6[1], addr_131_6, addr_positional[2103:2100], addr_525_7);

wire[31:0] addr_526_7;

Selector_2 s526_7(wires_131_6[2], addr_131_6, addr_positional[2107:2104], addr_526_7);

wire[31:0] addr_527_7;

Selector_2 s527_7(wires_131_6[3], addr_131_6, addr_positional[2111:2108], addr_527_7);

wire[31:0] addr_528_7;

Selector_2 s528_7(wires_132_6[0], addr_132_6, addr_positional[2115:2112], addr_528_7);

wire[31:0] addr_529_7;

Selector_2 s529_7(wires_132_6[1], addr_132_6, addr_positional[2119:2116], addr_529_7);

wire[31:0] addr_530_7;

Selector_2 s530_7(wires_132_6[2], addr_132_6, addr_positional[2123:2120], addr_530_7);

wire[31:0] addr_531_7;

Selector_2 s531_7(wires_132_6[3], addr_132_6, addr_positional[2127:2124], addr_531_7);

wire[31:0] addr_532_7;

Selector_2 s532_7(wires_133_6[0], addr_133_6, addr_positional[2131:2128], addr_532_7);

wire[31:0] addr_533_7;

Selector_2 s533_7(wires_133_6[1], addr_133_6, addr_positional[2135:2132], addr_533_7);

wire[31:0] addr_534_7;

Selector_2 s534_7(wires_133_6[2], addr_133_6, addr_positional[2139:2136], addr_534_7);

wire[31:0] addr_535_7;

Selector_2 s535_7(wires_133_6[3], addr_133_6, addr_positional[2143:2140], addr_535_7);

wire[31:0] addr_536_7;

Selector_2 s536_7(wires_134_6[0], addr_134_6, addr_positional[2147:2144], addr_536_7);

wire[31:0] addr_537_7;

Selector_2 s537_7(wires_134_6[1], addr_134_6, addr_positional[2151:2148], addr_537_7);

wire[31:0] addr_538_7;

Selector_2 s538_7(wires_134_6[2], addr_134_6, addr_positional[2155:2152], addr_538_7);

wire[31:0] addr_539_7;

Selector_2 s539_7(wires_134_6[3], addr_134_6, addr_positional[2159:2156], addr_539_7);

wire[31:0] addr_540_7;

Selector_2 s540_7(wires_135_6[0], addr_135_6, addr_positional[2163:2160], addr_540_7);

wire[31:0] addr_541_7;

Selector_2 s541_7(wires_135_6[1], addr_135_6, addr_positional[2167:2164], addr_541_7);

wire[31:0] addr_542_7;

Selector_2 s542_7(wires_135_6[2], addr_135_6, addr_positional[2171:2168], addr_542_7);

wire[31:0] addr_543_7;

Selector_2 s543_7(wires_135_6[3], addr_135_6, addr_positional[2175:2172], addr_543_7);

wire[31:0] addr_544_7;

Selector_2 s544_7(wires_136_6[0], addr_136_6, addr_positional[2179:2176], addr_544_7);

wire[31:0] addr_545_7;

Selector_2 s545_7(wires_136_6[1], addr_136_6, addr_positional[2183:2180], addr_545_7);

wire[31:0] addr_546_7;

Selector_2 s546_7(wires_136_6[2], addr_136_6, addr_positional[2187:2184], addr_546_7);

wire[31:0] addr_547_7;

Selector_2 s547_7(wires_136_6[3], addr_136_6, addr_positional[2191:2188], addr_547_7);

wire[31:0] addr_548_7;

Selector_2 s548_7(wires_137_6[0], addr_137_6, addr_positional[2195:2192], addr_548_7);

wire[31:0] addr_549_7;

Selector_2 s549_7(wires_137_6[1], addr_137_6, addr_positional[2199:2196], addr_549_7);

wire[31:0] addr_550_7;

Selector_2 s550_7(wires_137_6[2], addr_137_6, addr_positional[2203:2200], addr_550_7);

wire[31:0] addr_551_7;

Selector_2 s551_7(wires_137_6[3], addr_137_6, addr_positional[2207:2204], addr_551_7);

wire[31:0] addr_552_7;

Selector_2 s552_7(wires_138_6[0], addr_138_6, addr_positional[2211:2208], addr_552_7);

wire[31:0] addr_553_7;

Selector_2 s553_7(wires_138_6[1], addr_138_6, addr_positional[2215:2212], addr_553_7);

wire[31:0] addr_554_7;

Selector_2 s554_7(wires_138_6[2], addr_138_6, addr_positional[2219:2216], addr_554_7);

wire[31:0] addr_555_7;

Selector_2 s555_7(wires_138_6[3], addr_138_6, addr_positional[2223:2220], addr_555_7);

wire[31:0] addr_556_7;

Selector_2 s556_7(wires_139_6[0], addr_139_6, addr_positional[2227:2224], addr_556_7);

wire[31:0] addr_557_7;

Selector_2 s557_7(wires_139_6[1], addr_139_6, addr_positional[2231:2228], addr_557_7);

wire[31:0] addr_558_7;

Selector_2 s558_7(wires_139_6[2], addr_139_6, addr_positional[2235:2232], addr_558_7);

wire[31:0] addr_559_7;

Selector_2 s559_7(wires_139_6[3], addr_139_6, addr_positional[2239:2236], addr_559_7);

wire[31:0] addr_560_7;

Selector_2 s560_7(wires_140_6[0], addr_140_6, addr_positional[2243:2240], addr_560_7);

wire[31:0] addr_561_7;

Selector_2 s561_7(wires_140_6[1], addr_140_6, addr_positional[2247:2244], addr_561_7);

wire[31:0] addr_562_7;

Selector_2 s562_7(wires_140_6[2], addr_140_6, addr_positional[2251:2248], addr_562_7);

wire[31:0] addr_563_7;

Selector_2 s563_7(wires_140_6[3], addr_140_6, addr_positional[2255:2252], addr_563_7);

wire[31:0] addr_564_7;

Selector_2 s564_7(wires_141_6[0], addr_141_6, addr_positional[2259:2256], addr_564_7);

wire[31:0] addr_565_7;

Selector_2 s565_7(wires_141_6[1], addr_141_6, addr_positional[2263:2260], addr_565_7);

wire[31:0] addr_566_7;

Selector_2 s566_7(wires_141_6[2], addr_141_6, addr_positional[2267:2264], addr_566_7);

wire[31:0] addr_567_7;

Selector_2 s567_7(wires_141_6[3], addr_141_6, addr_positional[2271:2268], addr_567_7);

wire[31:0] addr_568_7;

Selector_2 s568_7(wires_142_6[0], addr_142_6, addr_positional[2275:2272], addr_568_7);

wire[31:0] addr_569_7;

Selector_2 s569_7(wires_142_6[1], addr_142_6, addr_positional[2279:2276], addr_569_7);

wire[31:0] addr_570_7;

Selector_2 s570_7(wires_142_6[2], addr_142_6, addr_positional[2283:2280], addr_570_7);

wire[31:0] addr_571_7;

Selector_2 s571_7(wires_142_6[3], addr_142_6, addr_positional[2287:2284], addr_571_7);

wire[31:0] addr_572_7;

Selector_2 s572_7(wires_143_6[0], addr_143_6, addr_positional[2291:2288], addr_572_7);

wire[31:0] addr_573_7;

Selector_2 s573_7(wires_143_6[1], addr_143_6, addr_positional[2295:2292], addr_573_7);

wire[31:0] addr_574_7;

Selector_2 s574_7(wires_143_6[2], addr_143_6, addr_positional[2299:2296], addr_574_7);

wire[31:0] addr_575_7;

Selector_2 s575_7(wires_143_6[3], addr_143_6, addr_positional[2303:2300], addr_575_7);

wire[31:0] addr_576_7;

Selector_2 s576_7(wires_144_6[0], addr_144_6, addr_positional[2307:2304], addr_576_7);

wire[31:0] addr_577_7;

Selector_2 s577_7(wires_144_6[1], addr_144_6, addr_positional[2311:2308], addr_577_7);

wire[31:0] addr_578_7;

Selector_2 s578_7(wires_144_6[2], addr_144_6, addr_positional[2315:2312], addr_578_7);

wire[31:0] addr_579_7;

Selector_2 s579_7(wires_144_6[3], addr_144_6, addr_positional[2319:2316], addr_579_7);

wire[31:0] addr_580_7;

Selector_2 s580_7(wires_145_6[0], addr_145_6, addr_positional[2323:2320], addr_580_7);

wire[31:0] addr_581_7;

Selector_2 s581_7(wires_145_6[1], addr_145_6, addr_positional[2327:2324], addr_581_7);

wire[31:0] addr_582_7;

Selector_2 s582_7(wires_145_6[2], addr_145_6, addr_positional[2331:2328], addr_582_7);

wire[31:0] addr_583_7;

Selector_2 s583_7(wires_145_6[3], addr_145_6, addr_positional[2335:2332], addr_583_7);

wire[31:0] addr_584_7;

Selector_2 s584_7(wires_146_6[0], addr_146_6, addr_positional[2339:2336], addr_584_7);

wire[31:0] addr_585_7;

Selector_2 s585_7(wires_146_6[1], addr_146_6, addr_positional[2343:2340], addr_585_7);

wire[31:0] addr_586_7;

Selector_2 s586_7(wires_146_6[2], addr_146_6, addr_positional[2347:2344], addr_586_7);

wire[31:0] addr_587_7;

Selector_2 s587_7(wires_146_6[3], addr_146_6, addr_positional[2351:2348], addr_587_7);

wire[31:0] addr_588_7;

Selector_2 s588_7(wires_147_6[0], addr_147_6, addr_positional[2355:2352], addr_588_7);

wire[31:0] addr_589_7;

Selector_2 s589_7(wires_147_6[1], addr_147_6, addr_positional[2359:2356], addr_589_7);

wire[31:0] addr_590_7;

Selector_2 s590_7(wires_147_6[2], addr_147_6, addr_positional[2363:2360], addr_590_7);

wire[31:0] addr_591_7;

Selector_2 s591_7(wires_147_6[3], addr_147_6, addr_positional[2367:2364], addr_591_7);

wire[31:0] addr_592_7;

Selector_2 s592_7(wires_148_6[0], addr_148_6, addr_positional[2371:2368], addr_592_7);

wire[31:0] addr_593_7;

Selector_2 s593_7(wires_148_6[1], addr_148_6, addr_positional[2375:2372], addr_593_7);

wire[31:0] addr_594_7;

Selector_2 s594_7(wires_148_6[2], addr_148_6, addr_positional[2379:2376], addr_594_7);

wire[31:0] addr_595_7;

Selector_2 s595_7(wires_148_6[3], addr_148_6, addr_positional[2383:2380], addr_595_7);

wire[31:0] addr_596_7;

Selector_2 s596_7(wires_149_6[0], addr_149_6, addr_positional[2387:2384], addr_596_7);

wire[31:0] addr_597_7;

Selector_2 s597_7(wires_149_6[1], addr_149_6, addr_positional[2391:2388], addr_597_7);

wire[31:0] addr_598_7;

Selector_2 s598_7(wires_149_6[2], addr_149_6, addr_positional[2395:2392], addr_598_7);

wire[31:0] addr_599_7;

Selector_2 s599_7(wires_149_6[3], addr_149_6, addr_positional[2399:2396], addr_599_7);

wire[31:0] addr_600_7;

Selector_2 s600_7(wires_150_6[0], addr_150_6, addr_positional[2403:2400], addr_600_7);

wire[31:0] addr_601_7;

Selector_2 s601_7(wires_150_6[1], addr_150_6, addr_positional[2407:2404], addr_601_7);

wire[31:0] addr_602_7;

Selector_2 s602_7(wires_150_6[2], addr_150_6, addr_positional[2411:2408], addr_602_7);

wire[31:0] addr_603_7;

Selector_2 s603_7(wires_150_6[3], addr_150_6, addr_positional[2415:2412], addr_603_7);

wire[31:0] addr_604_7;

Selector_2 s604_7(wires_151_6[0], addr_151_6, addr_positional[2419:2416], addr_604_7);

wire[31:0] addr_605_7;

Selector_2 s605_7(wires_151_6[1], addr_151_6, addr_positional[2423:2420], addr_605_7);

wire[31:0] addr_606_7;

Selector_2 s606_7(wires_151_6[2], addr_151_6, addr_positional[2427:2424], addr_606_7);

wire[31:0] addr_607_7;

Selector_2 s607_7(wires_151_6[3], addr_151_6, addr_positional[2431:2428], addr_607_7);

wire[31:0] addr_608_7;

Selector_2 s608_7(wires_152_6[0], addr_152_6, addr_positional[2435:2432], addr_608_7);

wire[31:0] addr_609_7;

Selector_2 s609_7(wires_152_6[1], addr_152_6, addr_positional[2439:2436], addr_609_7);

wire[31:0] addr_610_7;

Selector_2 s610_7(wires_152_6[2], addr_152_6, addr_positional[2443:2440], addr_610_7);

wire[31:0] addr_611_7;

Selector_2 s611_7(wires_152_6[3], addr_152_6, addr_positional[2447:2444], addr_611_7);

wire[31:0] addr_612_7;

Selector_2 s612_7(wires_153_6[0], addr_153_6, addr_positional[2451:2448], addr_612_7);

wire[31:0] addr_613_7;

Selector_2 s613_7(wires_153_6[1], addr_153_6, addr_positional[2455:2452], addr_613_7);

wire[31:0] addr_614_7;

Selector_2 s614_7(wires_153_6[2], addr_153_6, addr_positional[2459:2456], addr_614_7);

wire[31:0] addr_615_7;

Selector_2 s615_7(wires_153_6[3], addr_153_6, addr_positional[2463:2460], addr_615_7);

wire[31:0] addr_616_7;

Selector_2 s616_7(wires_154_6[0], addr_154_6, addr_positional[2467:2464], addr_616_7);

wire[31:0] addr_617_7;

Selector_2 s617_7(wires_154_6[1], addr_154_6, addr_positional[2471:2468], addr_617_7);

wire[31:0] addr_618_7;

Selector_2 s618_7(wires_154_6[2], addr_154_6, addr_positional[2475:2472], addr_618_7);

wire[31:0] addr_619_7;

Selector_2 s619_7(wires_154_6[3], addr_154_6, addr_positional[2479:2476], addr_619_7);

wire[31:0] addr_620_7;

Selector_2 s620_7(wires_155_6[0], addr_155_6, addr_positional[2483:2480], addr_620_7);

wire[31:0] addr_621_7;

Selector_2 s621_7(wires_155_6[1], addr_155_6, addr_positional[2487:2484], addr_621_7);

wire[31:0] addr_622_7;

Selector_2 s622_7(wires_155_6[2], addr_155_6, addr_positional[2491:2488], addr_622_7);

wire[31:0] addr_623_7;

Selector_2 s623_7(wires_155_6[3], addr_155_6, addr_positional[2495:2492], addr_623_7);

wire[31:0] addr_624_7;

Selector_2 s624_7(wires_156_6[0], addr_156_6, addr_positional[2499:2496], addr_624_7);

wire[31:0] addr_625_7;

Selector_2 s625_7(wires_156_6[1], addr_156_6, addr_positional[2503:2500], addr_625_7);

wire[31:0] addr_626_7;

Selector_2 s626_7(wires_156_6[2], addr_156_6, addr_positional[2507:2504], addr_626_7);

wire[31:0] addr_627_7;

Selector_2 s627_7(wires_156_6[3], addr_156_6, addr_positional[2511:2508], addr_627_7);

wire[31:0] addr_628_7;

Selector_2 s628_7(wires_157_6[0], addr_157_6, addr_positional[2515:2512], addr_628_7);

wire[31:0] addr_629_7;

Selector_2 s629_7(wires_157_6[1], addr_157_6, addr_positional[2519:2516], addr_629_7);

wire[31:0] addr_630_7;

Selector_2 s630_7(wires_157_6[2], addr_157_6, addr_positional[2523:2520], addr_630_7);

wire[31:0] addr_631_7;

Selector_2 s631_7(wires_157_6[3], addr_157_6, addr_positional[2527:2524], addr_631_7);

wire[31:0] addr_632_7;

Selector_2 s632_7(wires_158_6[0], addr_158_6, addr_positional[2531:2528], addr_632_7);

wire[31:0] addr_633_7;

Selector_2 s633_7(wires_158_6[1], addr_158_6, addr_positional[2535:2532], addr_633_7);

wire[31:0] addr_634_7;

Selector_2 s634_7(wires_158_6[2], addr_158_6, addr_positional[2539:2536], addr_634_7);

wire[31:0] addr_635_7;

Selector_2 s635_7(wires_158_6[3], addr_158_6, addr_positional[2543:2540], addr_635_7);

wire[31:0] addr_636_7;

Selector_2 s636_7(wires_159_6[0], addr_159_6, addr_positional[2547:2544], addr_636_7);

wire[31:0] addr_637_7;

Selector_2 s637_7(wires_159_6[1], addr_159_6, addr_positional[2551:2548], addr_637_7);

wire[31:0] addr_638_7;

Selector_2 s638_7(wires_159_6[2], addr_159_6, addr_positional[2555:2552], addr_638_7);

wire[31:0] addr_639_7;

Selector_2 s639_7(wires_159_6[3], addr_159_6, addr_positional[2559:2556], addr_639_7);

wire[31:0] addr_640_7;

Selector_2 s640_7(wires_160_6[0], addr_160_6, addr_positional[2563:2560], addr_640_7);

wire[31:0] addr_641_7;

Selector_2 s641_7(wires_160_6[1], addr_160_6, addr_positional[2567:2564], addr_641_7);

wire[31:0] addr_642_7;

Selector_2 s642_7(wires_160_6[2], addr_160_6, addr_positional[2571:2568], addr_642_7);

wire[31:0] addr_643_7;

Selector_2 s643_7(wires_160_6[3], addr_160_6, addr_positional[2575:2572], addr_643_7);

wire[31:0] addr_644_7;

Selector_2 s644_7(wires_161_6[0], addr_161_6, addr_positional[2579:2576], addr_644_7);

wire[31:0] addr_645_7;

Selector_2 s645_7(wires_161_6[1], addr_161_6, addr_positional[2583:2580], addr_645_7);

wire[31:0] addr_646_7;

Selector_2 s646_7(wires_161_6[2], addr_161_6, addr_positional[2587:2584], addr_646_7);

wire[31:0] addr_647_7;

Selector_2 s647_7(wires_161_6[3], addr_161_6, addr_positional[2591:2588], addr_647_7);

wire[31:0] addr_648_7;

Selector_2 s648_7(wires_162_6[0], addr_162_6, addr_positional[2595:2592], addr_648_7);

wire[31:0] addr_649_7;

Selector_2 s649_7(wires_162_6[1], addr_162_6, addr_positional[2599:2596], addr_649_7);

wire[31:0] addr_650_7;

Selector_2 s650_7(wires_162_6[2], addr_162_6, addr_positional[2603:2600], addr_650_7);

wire[31:0] addr_651_7;

Selector_2 s651_7(wires_162_6[3], addr_162_6, addr_positional[2607:2604], addr_651_7);

wire[31:0] addr_652_7;

Selector_2 s652_7(wires_163_6[0], addr_163_6, addr_positional[2611:2608], addr_652_7);

wire[31:0] addr_653_7;

Selector_2 s653_7(wires_163_6[1], addr_163_6, addr_positional[2615:2612], addr_653_7);

wire[31:0] addr_654_7;

Selector_2 s654_7(wires_163_6[2], addr_163_6, addr_positional[2619:2616], addr_654_7);

wire[31:0] addr_655_7;

Selector_2 s655_7(wires_163_6[3], addr_163_6, addr_positional[2623:2620], addr_655_7);

wire[31:0] addr_656_7;

Selector_2 s656_7(wires_164_6[0], addr_164_6, addr_positional[2627:2624], addr_656_7);

wire[31:0] addr_657_7;

Selector_2 s657_7(wires_164_6[1], addr_164_6, addr_positional[2631:2628], addr_657_7);

wire[31:0] addr_658_7;

Selector_2 s658_7(wires_164_6[2], addr_164_6, addr_positional[2635:2632], addr_658_7);

wire[31:0] addr_659_7;

Selector_2 s659_7(wires_164_6[3], addr_164_6, addr_positional[2639:2636], addr_659_7);

wire[31:0] addr_660_7;

Selector_2 s660_7(wires_165_6[0], addr_165_6, addr_positional[2643:2640], addr_660_7);

wire[31:0] addr_661_7;

Selector_2 s661_7(wires_165_6[1], addr_165_6, addr_positional[2647:2644], addr_661_7);

wire[31:0] addr_662_7;

Selector_2 s662_7(wires_165_6[2], addr_165_6, addr_positional[2651:2648], addr_662_7);

wire[31:0] addr_663_7;

Selector_2 s663_7(wires_165_6[3], addr_165_6, addr_positional[2655:2652], addr_663_7);

wire[31:0] addr_664_7;

Selector_2 s664_7(wires_166_6[0], addr_166_6, addr_positional[2659:2656], addr_664_7);

wire[31:0] addr_665_7;

Selector_2 s665_7(wires_166_6[1], addr_166_6, addr_positional[2663:2660], addr_665_7);

wire[31:0] addr_666_7;

Selector_2 s666_7(wires_166_6[2], addr_166_6, addr_positional[2667:2664], addr_666_7);

wire[31:0] addr_667_7;

Selector_2 s667_7(wires_166_6[3], addr_166_6, addr_positional[2671:2668], addr_667_7);

wire[31:0] addr_668_7;

Selector_2 s668_7(wires_167_6[0], addr_167_6, addr_positional[2675:2672], addr_668_7);

wire[31:0] addr_669_7;

Selector_2 s669_7(wires_167_6[1], addr_167_6, addr_positional[2679:2676], addr_669_7);

wire[31:0] addr_670_7;

Selector_2 s670_7(wires_167_6[2], addr_167_6, addr_positional[2683:2680], addr_670_7);

wire[31:0] addr_671_7;

Selector_2 s671_7(wires_167_6[3], addr_167_6, addr_positional[2687:2684], addr_671_7);

wire[31:0] addr_672_7;

Selector_2 s672_7(wires_168_6[0], addr_168_6, addr_positional[2691:2688], addr_672_7);

wire[31:0] addr_673_7;

Selector_2 s673_7(wires_168_6[1], addr_168_6, addr_positional[2695:2692], addr_673_7);

wire[31:0] addr_674_7;

Selector_2 s674_7(wires_168_6[2], addr_168_6, addr_positional[2699:2696], addr_674_7);

wire[31:0] addr_675_7;

Selector_2 s675_7(wires_168_6[3], addr_168_6, addr_positional[2703:2700], addr_675_7);

wire[31:0] addr_676_7;

Selector_2 s676_7(wires_169_6[0], addr_169_6, addr_positional[2707:2704], addr_676_7);

wire[31:0] addr_677_7;

Selector_2 s677_7(wires_169_6[1], addr_169_6, addr_positional[2711:2708], addr_677_7);

wire[31:0] addr_678_7;

Selector_2 s678_7(wires_169_6[2], addr_169_6, addr_positional[2715:2712], addr_678_7);

wire[31:0] addr_679_7;

Selector_2 s679_7(wires_169_6[3], addr_169_6, addr_positional[2719:2716], addr_679_7);

wire[31:0] addr_680_7;

Selector_2 s680_7(wires_170_6[0], addr_170_6, addr_positional[2723:2720], addr_680_7);

wire[31:0] addr_681_7;

Selector_2 s681_7(wires_170_6[1], addr_170_6, addr_positional[2727:2724], addr_681_7);

wire[31:0] addr_682_7;

Selector_2 s682_7(wires_170_6[2], addr_170_6, addr_positional[2731:2728], addr_682_7);

wire[31:0] addr_683_7;

Selector_2 s683_7(wires_170_6[3], addr_170_6, addr_positional[2735:2732], addr_683_7);

wire[31:0] addr_684_7;

Selector_2 s684_7(wires_171_6[0], addr_171_6, addr_positional[2739:2736], addr_684_7);

wire[31:0] addr_685_7;

Selector_2 s685_7(wires_171_6[1], addr_171_6, addr_positional[2743:2740], addr_685_7);

wire[31:0] addr_686_7;

Selector_2 s686_7(wires_171_6[2], addr_171_6, addr_positional[2747:2744], addr_686_7);

wire[31:0] addr_687_7;

Selector_2 s687_7(wires_171_6[3], addr_171_6, addr_positional[2751:2748], addr_687_7);

wire[31:0] addr_688_7;

Selector_2 s688_7(wires_172_6[0], addr_172_6, addr_positional[2755:2752], addr_688_7);

wire[31:0] addr_689_7;

Selector_2 s689_7(wires_172_6[1], addr_172_6, addr_positional[2759:2756], addr_689_7);

wire[31:0] addr_690_7;

Selector_2 s690_7(wires_172_6[2], addr_172_6, addr_positional[2763:2760], addr_690_7);

wire[31:0] addr_691_7;

Selector_2 s691_7(wires_172_6[3], addr_172_6, addr_positional[2767:2764], addr_691_7);

wire[31:0] addr_692_7;

Selector_2 s692_7(wires_173_6[0], addr_173_6, addr_positional[2771:2768], addr_692_7);

wire[31:0] addr_693_7;

Selector_2 s693_7(wires_173_6[1], addr_173_6, addr_positional[2775:2772], addr_693_7);

wire[31:0] addr_694_7;

Selector_2 s694_7(wires_173_6[2], addr_173_6, addr_positional[2779:2776], addr_694_7);

wire[31:0] addr_695_7;

Selector_2 s695_7(wires_173_6[3], addr_173_6, addr_positional[2783:2780], addr_695_7);

wire[31:0] addr_696_7;

Selector_2 s696_7(wires_174_6[0], addr_174_6, addr_positional[2787:2784], addr_696_7);

wire[31:0] addr_697_7;

Selector_2 s697_7(wires_174_6[1], addr_174_6, addr_positional[2791:2788], addr_697_7);

wire[31:0] addr_698_7;

Selector_2 s698_7(wires_174_6[2], addr_174_6, addr_positional[2795:2792], addr_698_7);

wire[31:0] addr_699_7;

Selector_2 s699_7(wires_174_6[3], addr_174_6, addr_positional[2799:2796], addr_699_7);

wire[31:0] addr_700_7;

Selector_2 s700_7(wires_175_6[0], addr_175_6, addr_positional[2803:2800], addr_700_7);

wire[31:0] addr_701_7;

Selector_2 s701_7(wires_175_6[1], addr_175_6, addr_positional[2807:2804], addr_701_7);

wire[31:0] addr_702_7;

Selector_2 s702_7(wires_175_6[2], addr_175_6, addr_positional[2811:2808], addr_702_7);

wire[31:0] addr_703_7;

Selector_2 s703_7(wires_175_6[3], addr_175_6, addr_positional[2815:2812], addr_703_7);

wire[31:0] addr_704_7;

Selector_2 s704_7(wires_176_6[0], addr_176_6, addr_positional[2819:2816], addr_704_7);

wire[31:0] addr_705_7;

Selector_2 s705_7(wires_176_6[1], addr_176_6, addr_positional[2823:2820], addr_705_7);

wire[31:0] addr_706_7;

Selector_2 s706_7(wires_176_6[2], addr_176_6, addr_positional[2827:2824], addr_706_7);

wire[31:0] addr_707_7;

Selector_2 s707_7(wires_176_6[3], addr_176_6, addr_positional[2831:2828], addr_707_7);

wire[31:0] addr_708_7;

Selector_2 s708_7(wires_177_6[0], addr_177_6, addr_positional[2835:2832], addr_708_7);

wire[31:0] addr_709_7;

Selector_2 s709_7(wires_177_6[1], addr_177_6, addr_positional[2839:2836], addr_709_7);

wire[31:0] addr_710_7;

Selector_2 s710_7(wires_177_6[2], addr_177_6, addr_positional[2843:2840], addr_710_7);

wire[31:0] addr_711_7;

Selector_2 s711_7(wires_177_6[3], addr_177_6, addr_positional[2847:2844], addr_711_7);

wire[31:0] addr_712_7;

Selector_2 s712_7(wires_178_6[0], addr_178_6, addr_positional[2851:2848], addr_712_7);

wire[31:0] addr_713_7;

Selector_2 s713_7(wires_178_6[1], addr_178_6, addr_positional[2855:2852], addr_713_7);

wire[31:0] addr_714_7;

Selector_2 s714_7(wires_178_6[2], addr_178_6, addr_positional[2859:2856], addr_714_7);

wire[31:0] addr_715_7;

Selector_2 s715_7(wires_178_6[3], addr_178_6, addr_positional[2863:2860], addr_715_7);

wire[31:0] addr_716_7;

Selector_2 s716_7(wires_179_6[0], addr_179_6, addr_positional[2867:2864], addr_716_7);

wire[31:0] addr_717_7;

Selector_2 s717_7(wires_179_6[1], addr_179_6, addr_positional[2871:2868], addr_717_7);

wire[31:0] addr_718_7;

Selector_2 s718_7(wires_179_6[2], addr_179_6, addr_positional[2875:2872], addr_718_7);

wire[31:0] addr_719_7;

Selector_2 s719_7(wires_179_6[3], addr_179_6, addr_positional[2879:2876], addr_719_7);

wire[31:0] addr_720_7;

Selector_2 s720_7(wires_180_6[0], addr_180_6, addr_positional[2883:2880], addr_720_7);

wire[31:0] addr_721_7;

Selector_2 s721_7(wires_180_6[1], addr_180_6, addr_positional[2887:2884], addr_721_7);

wire[31:0] addr_722_7;

Selector_2 s722_7(wires_180_6[2], addr_180_6, addr_positional[2891:2888], addr_722_7);

wire[31:0] addr_723_7;

Selector_2 s723_7(wires_180_6[3], addr_180_6, addr_positional[2895:2892], addr_723_7);

wire[31:0] addr_724_7;

Selector_2 s724_7(wires_181_6[0], addr_181_6, addr_positional[2899:2896], addr_724_7);

wire[31:0] addr_725_7;

Selector_2 s725_7(wires_181_6[1], addr_181_6, addr_positional[2903:2900], addr_725_7);

wire[31:0] addr_726_7;

Selector_2 s726_7(wires_181_6[2], addr_181_6, addr_positional[2907:2904], addr_726_7);

wire[31:0] addr_727_7;

Selector_2 s727_7(wires_181_6[3], addr_181_6, addr_positional[2911:2908], addr_727_7);

wire[31:0] addr_728_7;

Selector_2 s728_7(wires_182_6[0], addr_182_6, addr_positional[2915:2912], addr_728_7);

wire[31:0] addr_729_7;

Selector_2 s729_7(wires_182_6[1], addr_182_6, addr_positional[2919:2916], addr_729_7);

wire[31:0] addr_730_7;

Selector_2 s730_7(wires_182_6[2], addr_182_6, addr_positional[2923:2920], addr_730_7);

wire[31:0] addr_731_7;

Selector_2 s731_7(wires_182_6[3], addr_182_6, addr_positional[2927:2924], addr_731_7);

wire[31:0] addr_732_7;

Selector_2 s732_7(wires_183_6[0], addr_183_6, addr_positional[2931:2928], addr_732_7);

wire[31:0] addr_733_7;

Selector_2 s733_7(wires_183_6[1], addr_183_6, addr_positional[2935:2932], addr_733_7);

wire[31:0] addr_734_7;

Selector_2 s734_7(wires_183_6[2], addr_183_6, addr_positional[2939:2936], addr_734_7);

wire[31:0] addr_735_7;

Selector_2 s735_7(wires_183_6[3], addr_183_6, addr_positional[2943:2940], addr_735_7);

wire[31:0] addr_736_7;

Selector_2 s736_7(wires_184_6[0], addr_184_6, addr_positional[2947:2944], addr_736_7);

wire[31:0] addr_737_7;

Selector_2 s737_7(wires_184_6[1], addr_184_6, addr_positional[2951:2948], addr_737_7);

wire[31:0] addr_738_7;

Selector_2 s738_7(wires_184_6[2], addr_184_6, addr_positional[2955:2952], addr_738_7);

wire[31:0] addr_739_7;

Selector_2 s739_7(wires_184_6[3], addr_184_6, addr_positional[2959:2956], addr_739_7);

wire[31:0] addr_740_7;

Selector_2 s740_7(wires_185_6[0], addr_185_6, addr_positional[2963:2960], addr_740_7);

wire[31:0] addr_741_7;

Selector_2 s741_7(wires_185_6[1], addr_185_6, addr_positional[2967:2964], addr_741_7);

wire[31:0] addr_742_7;

Selector_2 s742_7(wires_185_6[2], addr_185_6, addr_positional[2971:2968], addr_742_7);

wire[31:0] addr_743_7;

Selector_2 s743_7(wires_185_6[3], addr_185_6, addr_positional[2975:2972], addr_743_7);

wire[31:0] addr_744_7;

Selector_2 s744_7(wires_186_6[0], addr_186_6, addr_positional[2979:2976], addr_744_7);

wire[31:0] addr_745_7;

Selector_2 s745_7(wires_186_6[1], addr_186_6, addr_positional[2983:2980], addr_745_7);

wire[31:0] addr_746_7;

Selector_2 s746_7(wires_186_6[2], addr_186_6, addr_positional[2987:2984], addr_746_7);

wire[31:0] addr_747_7;

Selector_2 s747_7(wires_186_6[3], addr_186_6, addr_positional[2991:2988], addr_747_7);

wire[31:0] addr_748_7;

Selector_2 s748_7(wires_187_6[0], addr_187_6, addr_positional[2995:2992], addr_748_7);

wire[31:0] addr_749_7;

Selector_2 s749_7(wires_187_6[1], addr_187_6, addr_positional[2999:2996], addr_749_7);

wire[31:0] addr_750_7;

Selector_2 s750_7(wires_187_6[2], addr_187_6, addr_positional[3003:3000], addr_750_7);

wire[31:0] addr_751_7;

Selector_2 s751_7(wires_187_6[3], addr_187_6, addr_positional[3007:3004], addr_751_7);

wire[31:0] addr_752_7;

Selector_2 s752_7(wires_188_6[0], addr_188_6, addr_positional[3011:3008], addr_752_7);

wire[31:0] addr_753_7;

Selector_2 s753_7(wires_188_6[1], addr_188_6, addr_positional[3015:3012], addr_753_7);

wire[31:0] addr_754_7;

Selector_2 s754_7(wires_188_6[2], addr_188_6, addr_positional[3019:3016], addr_754_7);

wire[31:0] addr_755_7;

Selector_2 s755_7(wires_188_6[3], addr_188_6, addr_positional[3023:3020], addr_755_7);

wire[31:0] addr_756_7;

Selector_2 s756_7(wires_189_6[0], addr_189_6, addr_positional[3027:3024], addr_756_7);

wire[31:0] addr_757_7;

Selector_2 s757_7(wires_189_6[1], addr_189_6, addr_positional[3031:3028], addr_757_7);

wire[31:0] addr_758_7;

Selector_2 s758_7(wires_189_6[2], addr_189_6, addr_positional[3035:3032], addr_758_7);

wire[31:0] addr_759_7;

Selector_2 s759_7(wires_189_6[3], addr_189_6, addr_positional[3039:3036], addr_759_7);

wire[31:0] addr_760_7;

Selector_2 s760_7(wires_190_6[0], addr_190_6, addr_positional[3043:3040], addr_760_7);

wire[31:0] addr_761_7;

Selector_2 s761_7(wires_190_6[1], addr_190_6, addr_positional[3047:3044], addr_761_7);

wire[31:0] addr_762_7;

Selector_2 s762_7(wires_190_6[2], addr_190_6, addr_positional[3051:3048], addr_762_7);

wire[31:0] addr_763_7;

Selector_2 s763_7(wires_190_6[3], addr_190_6, addr_positional[3055:3052], addr_763_7);

wire[31:0] addr_764_7;

Selector_2 s764_7(wires_191_6[0], addr_191_6, addr_positional[3059:3056], addr_764_7);

wire[31:0] addr_765_7;

Selector_2 s765_7(wires_191_6[1], addr_191_6, addr_positional[3063:3060], addr_765_7);

wire[31:0] addr_766_7;

Selector_2 s766_7(wires_191_6[2], addr_191_6, addr_positional[3067:3064], addr_766_7);

wire[31:0] addr_767_7;

Selector_2 s767_7(wires_191_6[3], addr_191_6, addr_positional[3071:3068], addr_767_7);

wire[31:0] addr_768_7;

Selector_2 s768_7(wires_192_6[0], addr_192_6, addr_positional[3075:3072], addr_768_7);

wire[31:0] addr_769_7;

Selector_2 s769_7(wires_192_6[1], addr_192_6, addr_positional[3079:3076], addr_769_7);

wire[31:0] addr_770_7;

Selector_2 s770_7(wires_192_6[2], addr_192_6, addr_positional[3083:3080], addr_770_7);

wire[31:0] addr_771_7;

Selector_2 s771_7(wires_192_6[3], addr_192_6, addr_positional[3087:3084], addr_771_7);

wire[31:0] addr_772_7;

Selector_2 s772_7(wires_193_6[0], addr_193_6, addr_positional[3091:3088], addr_772_7);

wire[31:0] addr_773_7;

Selector_2 s773_7(wires_193_6[1], addr_193_6, addr_positional[3095:3092], addr_773_7);

wire[31:0] addr_774_7;

Selector_2 s774_7(wires_193_6[2], addr_193_6, addr_positional[3099:3096], addr_774_7);

wire[31:0] addr_775_7;

Selector_2 s775_7(wires_193_6[3], addr_193_6, addr_positional[3103:3100], addr_775_7);

wire[31:0] addr_776_7;

Selector_2 s776_7(wires_194_6[0], addr_194_6, addr_positional[3107:3104], addr_776_7);

wire[31:0] addr_777_7;

Selector_2 s777_7(wires_194_6[1], addr_194_6, addr_positional[3111:3108], addr_777_7);

wire[31:0] addr_778_7;

Selector_2 s778_7(wires_194_6[2], addr_194_6, addr_positional[3115:3112], addr_778_7);

wire[31:0] addr_779_7;

Selector_2 s779_7(wires_194_6[3], addr_194_6, addr_positional[3119:3116], addr_779_7);

wire[31:0] addr_780_7;

Selector_2 s780_7(wires_195_6[0], addr_195_6, addr_positional[3123:3120], addr_780_7);

wire[31:0] addr_781_7;

Selector_2 s781_7(wires_195_6[1], addr_195_6, addr_positional[3127:3124], addr_781_7);

wire[31:0] addr_782_7;

Selector_2 s782_7(wires_195_6[2], addr_195_6, addr_positional[3131:3128], addr_782_7);

wire[31:0] addr_783_7;

Selector_2 s783_7(wires_195_6[3], addr_195_6, addr_positional[3135:3132], addr_783_7);

wire[31:0] addr_784_7;

Selector_2 s784_7(wires_196_6[0], addr_196_6, addr_positional[3139:3136], addr_784_7);

wire[31:0] addr_785_7;

Selector_2 s785_7(wires_196_6[1], addr_196_6, addr_positional[3143:3140], addr_785_7);

wire[31:0] addr_786_7;

Selector_2 s786_7(wires_196_6[2], addr_196_6, addr_positional[3147:3144], addr_786_7);

wire[31:0] addr_787_7;

Selector_2 s787_7(wires_196_6[3], addr_196_6, addr_positional[3151:3148], addr_787_7);

wire[31:0] addr_788_7;

Selector_2 s788_7(wires_197_6[0], addr_197_6, addr_positional[3155:3152], addr_788_7);

wire[31:0] addr_789_7;

Selector_2 s789_7(wires_197_6[1], addr_197_6, addr_positional[3159:3156], addr_789_7);

wire[31:0] addr_790_7;

Selector_2 s790_7(wires_197_6[2], addr_197_6, addr_positional[3163:3160], addr_790_7);

wire[31:0] addr_791_7;

Selector_2 s791_7(wires_197_6[3], addr_197_6, addr_positional[3167:3164], addr_791_7);

wire[31:0] addr_792_7;

Selector_2 s792_7(wires_198_6[0], addr_198_6, addr_positional[3171:3168], addr_792_7);

wire[31:0] addr_793_7;

Selector_2 s793_7(wires_198_6[1], addr_198_6, addr_positional[3175:3172], addr_793_7);

wire[31:0] addr_794_7;

Selector_2 s794_7(wires_198_6[2], addr_198_6, addr_positional[3179:3176], addr_794_7);

wire[31:0] addr_795_7;

Selector_2 s795_7(wires_198_6[3], addr_198_6, addr_positional[3183:3180], addr_795_7);

wire[31:0] addr_796_7;

Selector_2 s796_7(wires_199_6[0], addr_199_6, addr_positional[3187:3184], addr_796_7);

wire[31:0] addr_797_7;

Selector_2 s797_7(wires_199_6[1], addr_199_6, addr_positional[3191:3188], addr_797_7);

wire[31:0] addr_798_7;

Selector_2 s798_7(wires_199_6[2], addr_199_6, addr_positional[3195:3192], addr_798_7);

wire[31:0] addr_799_7;

Selector_2 s799_7(wires_199_6[3], addr_199_6, addr_positional[3199:3196], addr_799_7);

wire[31:0] addr_800_7;

Selector_2 s800_7(wires_200_6[0], addr_200_6, addr_positional[3203:3200], addr_800_7);

wire[31:0] addr_801_7;

Selector_2 s801_7(wires_200_6[1], addr_200_6, addr_positional[3207:3204], addr_801_7);

wire[31:0] addr_802_7;

Selector_2 s802_7(wires_200_6[2], addr_200_6, addr_positional[3211:3208], addr_802_7);

wire[31:0] addr_803_7;

Selector_2 s803_7(wires_200_6[3], addr_200_6, addr_positional[3215:3212], addr_803_7);

wire[31:0] addr_804_7;

Selector_2 s804_7(wires_201_6[0], addr_201_6, addr_positional[3219:3216], addr_804_7);

wire[31:0] addr_805_7;

Selector_2 s805_7(wires_201_6[1], addr_201_6, addr_positional[3223:3220], addr_805_7);

wire[31:0] addr_806_7;

Selector_2 s806_7(wires_201_6[2], addr_201_6, addr_positional[3227:3224], addr_806_7);

wire[31:0] addr_807_7;

Selector_2 s807_7(wires_201_6[3], addr_201_6, addr_positional[3231:3228], addr_807_7);

wire[31:0] addr_808_7;

Selector_2 s808_7(wires_202_6[0], addr_202_6, addr_positional[3235:3232], addr_808_7);

wire[31:0] addr_809_7;

Selector_2 s809_7(wires_202_6[1], addr_202_6, addr_positional[3239:3236], addr_809_7);

wire[31:0] addr_810_7;

Selector_2 s810_7(wires_202_6[2], addr_202_6, addr_positional[3243:3240], addr_810_7);

wire[31:0] addr_811_7;

Selector_2 s811_7(wires_202_6[3], addr_202_6, addr_positional[3247:3244], addr_811_7);

wire[31:0] addr_812_7;

Selector_2 s812_7(wires_203_6[0], addr_203_6, addr_positional[3251:3248], addr_812_7);

wire[31:0] addr_813_7;

Selector_2 s813_7(wires_203_6[1], addr_203_6, addr_positional[3255:3252], addr_813_7);

wire[31:0] addr_814_7;

Selector_2 s814_7(wires_203_6[2], addr_203_6, addr_positional[3259:3256], addr_814_7);

wire[31:0] addr_815_7;

Selector_2 s815_7(wires_203_6[3], addr_203_6, addr_positional[3263:3260], addr_815_7);

wire[31:0] addr_816_7;

Selector_2 s816_7(wires_204_6[0], addr_204_6, addr_positional[3267:3264], addr_816_7);

wire[31:0] addr_817_7;

Selector_2 s817_7(wires_204_6[1], addr_204_6, addr_positional[3271:3268], addr_817_7);

wire[31:0] addr_818_7;

Selector_2 s818_7(wires_204_6[2], addr_204_6, addr_positional[3275:3272], addr_818_7);

wire[31:0] addr_819_7;

Selector_2 s819_7(wires_204_6[3], addr_204_6, addr_positional[3279:3276], addr_819_7);

wire[31:0] addr_820_7;

Selector_2 s820_7(wires_205_6[0], addr_205_6, addr_positional[3283:3280], addr_820_7);

wire[31:0] addr_821_7;

Selector_2 s821_7(wires_205_6[1], addr_205_6, addr_positional[3287:3284], addr_821_7);

wire[31:0] addr_822_7;

Selector_2 s822_7(wires_205_6[2], addr_205_6, addr_positional[3291:3288], addr_822_7);

wire[31:0] addr_823_7;

Selector_2 s823_7(wires_205_6[3], addr_205_6, addr_positional[3295:3292], addr_823_7);

wire[31:0] addr_824_7;

Selector_2 s824_7(wires_206_6[0], addr_206_6, addr_positional[3299:3296], addr_824_7);

wire[31:0] addr_825_7;

Selector_2 s825_7(wires_206_6[1], addr_206_6, addr_positional[3303:3300], addr_825_7);

wire[31:0] addr_826_7;

Selector_2 s826_7(wires_206_6[2], addr_206_6, addr_positional[3307:3304], addr_826_7);

wire[31:0] addr_827_7;

Selector_2 s827_7(wires_206_6[3], addr_206_6, addr_positional[3311:3308], addr_827_7);

wire[31:0] addr_828_7;

Selector_2 s828_7(wires_207_6[0], addr_207_6, addr_positional[3315:3312], addr_828_7);

wire[31:0] addr_829_7;

Selector_2 s829_7(wires_207_6[1], addr_207_6, addr_positional[3319:3316], addr_829_7);

wire[31:0] addr_830_7;

Selector_2 s830_7(wires_207_6[2], addr_207_6, addr_positional[3323:3320], addr_830_7);

wire[31:0] addr_831_7;

Selector_2 s831_7(wires_207_6[3], addr_207_6, addr_positional[3327:3324], addr_831_7);

wire[31:0] addr_832_7;

Selector_2 s832_7(wires_208_6[0], addr_208_6, addr_positional[3331:3328], addr_832_7);

wire[31:0] addr_833_7;

Selector_2 s833_7(wires_208_6[1], addr_208_6, addr_positional[3335:3332], addr_833_7);

wire[31:0] addr_834_7;

Selector_2 s834_7(wires_208_6[2], addr_208_6, addr_positional[3339:3336], addr_834_7);

wire[31:0] addr_835_7;

Selector_2 s835_7(wires_208_6[3], addr_208_6, addr_positional[3343:3340], addr_835_7);

wire[31:0] addr_836_7;

Selector_2 s836_7(wires_209_6[0], addr_209_6, addr_positional[3347:3344], addr_836_7);

wire[31:0] addr_837_7;

Selector_2 s837_7(wires_209_6[1], addr_209_6, addr_positional[3351:3348], addr_837_7);

wire[31:0] addr_838_7;

Selector_2 s838_7(wires_209_6[2], addr_209_6, addr_positional[3355:3352], addr_838_7);

wire[31:0] addr_839_7;

Selector_2 s839_7(wires_209_6[3], addr_209_6, addr_positional[3359:3356], addr_839_7);

wire[31:0] addr_840_7;

Selector_2 s840_7(wires_210_6[0], addr_210_6, addr_positional[3363:3360], addr_840_7);

wire[31:0] addr_841_7;

Selector_2 s841_7(wires_210_6[1], addr_210_6, addr_positional[3367:3364], addr_841_7);

wire[31:0] addr_842_7;

Selector_2 s842_7(wires_210_6[2], addr_210_6, addr_positional[3371:3368], addr_842_7);

wire[31:0] addr_843_7;

Selector_2 s843_7(wires_210_6[3], addr_210_6, addr_positional[3375:3372], addr_843_7);

wire[31:0] addr_844_7;

Selector_2 s844_7(wires_211_6[0], addr_211_6, addr_positional[3379:3376], addr_844_7);

wire[31:0] addr_845_7;

Selector_2 s845_7(wires_211_6[1], addr_211_6, addr_positional[3383:3380], addr_845_7);

wire[31:0] addr_846_7;

Selector_2 s846_7(wires_211_6[2], addr_211_6, addr_positional[3387:3384], addr_846_7);

wire[31:0] addr_847_7;

Selector_2 s847_7(wires_211_6[3], addr_211_6, addr_positional[3391:3388], addr_847_7);

wire[31:0] addr_848_7;

Selector_2 s848_7(wires_212_6[0], addr_212_6, addr_positional[3395:3392], addr_848_7);

wire[31:0] addr_849_7;

Selector_2 s849_7(wires_212_6[1], addr_212_6, addr_positional[3399:3396], addr_849_7);

wire[31:0] addr_850_7;

Selector_2 s850_7(wires_212_6[2], addr_212_6, addr_positional[3403:3400], addr_850_7);

wire[31:0] addr_851_7;

Selector_2 s851_7(wires_212_6[3], addr_212_6, addr_positional[3407:3404], addr_851_7);

wire[31:0] addr_852_7;

Selector_2 s852_7(wires_213_6[0], addr_213_6, addr_positional[3411:3408], addr_852_7);

wire[31:0] addr_853_7;

Selector_2 s853_7(wires_213_6[1], addr_213_6, addr_positional[3415:3412], addr_853_7);

wire[31:0] addr_854_7;

Selector_2 s854_7(wires_213_6[2], addr_213_6, addr_positional[3419:3416], addr_854_7);

wire[31:0] addr_855_7;

Selector_2 s855_7(wires_213_6[3], addr_213_6, addr_positional[3423:3420], addr_855_7);

wire[31:0] addr_856_7;

Selector_2 s856_7(wires_214_6[0], addr_214_6, addr_positional[3427:3424], addr_856_7);

wire[31:0] addr_857_7;

Selector_2 s857_7(wires_214_6[1], addr_214_6, addr_positional[3431:3428], addr_857_7);

wire[31:0] addr_858_7;

Selector_2 s858_7(wires_214_6[2], addr_214_6, addr_positional[3435:3432], addr_858_7);

wire[31:0] addr_859_7;

Selector_2 s859_7(wires_214_6[3], addr_214_6, addr_positional[3439:3436], addr_859_7);

wire[31:0] addr_860_7;

Selector_2 s860_7(wires_215_6[0], addr_215_6, addr_positional[3443:3440], addr_860_7);

wire[31:0] addr_861_7;

Selector_2 s861_7(wires_215_6[1], addr_215_6, addr_positional[3447:3444], addr_861_7);

wire[31:0] addr_862_7;

Selector_2 s862_7(wires_215_6[2], addr_215_6, addr_positional[3451:3448], addr_862_7);

wire[31:0] addr_863_7;

Selector_2 s863_7(wires_215_6[3], addr_215_6, addr_positional[3455:3452], addr_863_7);

wire[31:0] addr_864_7;

Selector_2 s864_7(wires_216_6[0], addr_216_6, addr_positional[3459:3456], addr_864_7);

wire[31:0] addr_865_7;

Selector_2 s865_7(wires_216_6[1], addr_216_6, addr_positional[3463:3460], addr_865_7);

wire[31:0] addr_866_7;

Selector_2 s866_7(wires_216_6[2], addr_216_6, addr_positional[3467:3464], addr_866_7);

wire[31:0] addr_867_7;

Selector_2 s867_7(wires_216_6[3], addr_216_6, addr_positional[3471:3468], addr_867_7);

wire[31:0] addr_868_7;

Selector_2 s868_7(wires_217_6[0], addr_217_6, addr_positional[3475:3472], addr_868_7);

wire[31:0] addr_869_7;

Selector_2 s869_7(wires_217_6[1], addr_217_6, addr_positional[3479:3476], addr_869_7);

wire[31:0] addr_870_7;

Selector_2 s870_7(wires_217_6[2], addr_217_6, addr_positional[3483:3480], addr_870_7);

wire[31:0] addr_871_7;

Selector_2 s871_7(wires_217_6[3], addr_217_6, addr_positional[3487:3484], addr_871_7);

wire[31:0] addr_872_7;

Selector_2 s872_7(wires_218_6[0], addr_218_6, addr_positional[3491:3488], addr_872_7);

wire[31:0] addr_873_7;

Selector_2 s873_7(wires_218_6[1], addr_218_6, addr_positional[3495:3492], addr_873_7);

wire[31:0] addr_874_7;

Selector_2 s874_7(wires_218_6[2], addr_218_6, addr_positional[3499:3496], addr_874_7);

wire[31:0] addr_875_7;

Selector_2 s875_7(wires_218_6[3], addr_218_6, addr_positional[3503:3500], addr_875_7);

wire[31:0] addr_876_7;

Selector_2 s876_7(wires_219_6[0], addr_219_6, addr_positional[3507:3504], addr_876_7);

wire[31:0] addr_877_7;

Selector_2 s877_7(wires_219_6[1], addr_219_6, addr_positional[3511:3508], addr_877_7);

wire[31:0] addr_878_7;

Selector_2 s878_7(wires_219_6[2], addr_219_6, addr_positional[3515:3512], addr_878_7);

wire[31:0] addr_879_7;

Selector_2 s879_7(wires_219_6[3], addr_219_6, addr_positional[3519:3516], addr_879_7);

wire[31:0] addr_880_7;

Selector_2 s880_7(wires_220_6[0], addr_220_6, addr_positional[3523:3520], addr_880_7);

wire[31:0] addr_881_7;

Selector_2 s881_7(wires_220_6[1], addr_220_6, addr_positional[3527:3524], addr_881_7);

wire[31:0] addr_882_7;

Selector_2 s882_7(wires_220_6[2], addr_220_6, addr_positional[3531:3528], addr_882_7);

wire[31:0] addr_883_7;

Selector_2 s883_7(wires_220_6[3], addr_220_6, addr_positional[3535:3532], addr_883_7);

wire[31:0] addr_884_7;

Selector_2 s884_7(wires_221_6[0], addr_221_6, addr_positional[3539:3536], addr_884_7);

wire[31:0] addr_885_7;

Selector_2 s885_7(wires_221_6[1], addr_221_6, addr_positional[3543:3540], addr_885_7);

wire[31:0] addr_886_7;

Selector_2 s886_7(wires_221_6[2], addr_221_6, addr_positional[3547:3544], addr_886_7);

wire[31:0] addr_887_7;

Selector_2 s887_7(wires_221_6[3], addr_221_6, addr_positional[3551:3548], addr_887_7);

wire[31:0] addr_888_7;

Selector_2 s888_7(wires_222_6[0], addr_222_6, addr_positional[3555:3552], addr_888_7);

wire[31:0] addr_889_7;

Selector_2 s889_7(wires_222_6[1], addr_222_6, addr_positional[3559:3556], addr_889_7);

wire[31:0] addr_890_7;

Selector_2 s890_7(wires_222_6[2], addr_222_6, addr_positional[3563:3560], addr_890_7);

wire[31:0] addr_891_7;

Selector_2 s891_7(wires_222_6[3], addr_222_6, addr_positional[3567:3564], addr_891_7);

wire[31:0] addr_892_7;

Selector_2 s892_7(wires_223_6[0], addr_223_6, addr_positional[3571:3568], addr_892_7);

wire[31:0] addr_893_7;

Selector_2 s893_7(wires_223_6[1], addr_223_6, addr_positional[3575:3572], addr_893_7);

wire[31:0] addr_894_7;

Selector_2 s894_7(wires_223_6[2], addr_223_6, addr_positional[3579:3576], addr_894_7);

wire[31:0] addr_895_7;

Selector_2 s895_7(wires_223_6[3], addr_223_6, addr_positional[3583:3580], addr_895_7);

wire[31:0] addr_896_7;

Selector_2 s896_7(wires_224_6[0], addr_224_6, addr_positional[3587:3584], addr_896_7);

wire[31:0] addr_897_7;

Selector_2 s897_7(wires_224_6[1], addr_224_6, addr_positional[3591:3588], addr_897_7);

wire[31:0] addr_898_7;

Selector_2 s898_7(wires_224_6[2], addr_224_6, addr_positional[3595:3592], addr_898_7);

wire[31:0] addr_899_7;

Selector_2 s899_7(wires_224_6[3], addr_224_6, addr_positional[3599:3596], addr_899_7);

wire[31:0] addr_900_7;

Selector_2 s900_7(wires_225_6[0], addr_225_6, addr_positional[3603:3600], addr_900_7);

wire[31:0] addr_901_7;

Selector_2 s901_7(wires_225_6[1], addr_225_6, addr_positional[3607:3604], addr_901_7);

wire[31:0] addr_902_7;

Selector_2 s902_7(wires_225_6[2], addr_225_6, addr_positional[3611:3608], addr_902_7);

wire[31:0] addr_903_7;

Selector_2 s903_7(wires_225_6[3], addr_225_6, addr_positional[3615:3612], addr_903_7);

wire[31:0] addr_904_7;

Selector_2 s904_7(wires_226_6[0], addr_226_6, addr_positional[3619:3616], addr_904_7);

wire[31:0] addr_905_7;

Selector_2 s905_7(wires_226_6[1], addr_226_6, addr_positional[3623:3620], addr_905_7);

wire[31:0] addr_906_7;

Selector_2 s906_7(wires_226_6[2], addr_226_6, addr_positional[3627:3624], addr_906_7);

wire[31:0] addr_907_7;

Selector_2 s907_7(wires_226_6[3], addr_226_6, addr_positional[3631:3628], addr_907_7);

wire[31:0] addr_908_7;

Selector_2 s908_7(wires_227_6[0], addr_227_6, addr_positional[3635:3632], addr_908_7);

wire[31:0] addr_909_7;

Selector_2 s909_7(wires_227_6[1], addr_227_6, addr_positional[3639:3636], addr_909_7);

wire[31:0] addr_910_7;

Selector_2 s910_7(wires_227_6[2], addr_227_6, addr_positional[3643:3640], addr_910_7);

wire[31:0] addr_911_7;

Selector_2 s911_7(wires_227_6[3], addr_227_6, addr_positional[3647:3644], addr_911_7);

wire[31:0] addr_912_7;

Selector_2 s912_7(wires_228_6[0], addr_228_6, addr_positional[3651:3648], addr_912_7);

wire[31:0] addr_913_7;

Selector_2 s913_7(wires_228_6[1], addr_228_6, addr_positional[3655:3652], addr_913_7);

wire[31:0] addr_914_7;

Selector_2 s914_7(wires_228_6[2], addr_228_6, addr_positional[3659:3656], addr_914_7);

wire[31:0] addr_915_7;

Selector_2 s915_7(wires_228_6[3], addr_228_6, addr_positional[3663:3660], addr_915_7);

wire[31:0] addr_916_7;

Selector_2 s916_7(wires_229_6[0], addr_229_6, addr_positional[3667:3664], addr_916_7);

wire[31:0] addr_917_7;

Selector_2 s917_7(wires_229_6[1], addr_229_6, addr_positional[3671:3668], addr_917_7);

wire[31:0] addr_918_7;

Selector_2 s918_7(wires_229_6[2], addr_229_6, addr_positional[3675:3672], addr_918_7);

wire[31:0] addr_919_7;

Selector_2 s919_7(wires_229_6[3], addr_229_6, addr_positional[3679:3676], addr_919_7);

wire[31:0] addr_920_7;

Selector_2 s920_7(wires_230_6[0], addr_230_6, addr_positional[3683:3680], addr_920_7);

wire[31:0] addr_921_7;

Selector_2 s921_7(wires_230_6[1], addr_230_6, addr_positional[3687:3684], addr_921_7);

wire[31:0] addr_922_7;

Selector_2 s922_7(wires_230_6[2], addr_230_6, addr_positional[3691:3688], addr_922_7);

wire[31:0] addr_923_7;

Selector_2 s923_7(wires_230_6[3], addr_230_6, addr_positional[3695:3692], addr_923_7);

wire[31:0] addr_924_7;

Selector_2 s924_7(wires_231_6[0], addr_231_6, addr_positional[3699:3696], addr_924_7);

wire[31:0] addr_925_7;

Selector_2 s925_7(wires_231_6[1], addr_231_6, addr_positional[3703:3700], addr_925_7);

wire[31:0] addr_926_7;

Selector_2 s926_7(wires_231_6[2], addr_231_6, addr_positional[3707:3704], addr_926_7);

wire[31:0] addr_927_7;

Selector_2 s927_7(wires_231_6[3], addr_231_6, addr_positional[3711:3708], addr_927_7);

wire[31:0] addr_928_7;

Selector_2 s928_7(wires_232_6[0], addr_232_6, addr_positional[3715:3712], addr_928_7);

wire[31:0] addr_929_7;

Selector_2 s929_7(wires_232_6[1], addr_232_6, addr_positional[3719:3716], addr_929_7);

wire[31:0] addr_930_7;

Selector_2 s930_7(wires_232_6[2], addr_232_6, addr_positional[3723:3720], addr_930_7);

wire[31:0] addr_931_7;

Selector_2 s931_7(wires_232_6[3], addr_232_6, addr_positional[3727:3724], addr_931_7);

wire[31:0] addr_932_7;

Selector_2 s932_7(wires_233_6[0], addr_233_6, addr_positional[3731:3728], addr_932_7);

wire[31:0] addr_933_7;

Selector_2 s933_7(wires_233_6[1], addr_233_6, addr_positional[3735:3732], addr_933_7);

wire[31:0] addr_934_7;

Selector_2 s934_7(wires_233_6[2], addr_233_6, addr_positional[3739:3736], addr_934_7);

wire[31:0] addr_935_7;

Selector_2 s935_7(wires_233_6[3], addr_233_6, addr_positional[3743:3740], addr_935_7);

wire[31:0] addr_936_7;

Selector_2 s936_7(wires_234_6[0], addr_234_6, addr_positional[3747:3744], addr_936_7);

wire[31:0] addr_937_7;

Selector_2 s937_7(wires_234_6[1], addr_234_6, addr_positional[3751:3748], addr_937_7);

wire[31:0] addr_938_7;

Selector_2 s938_7(wires_234_6[2], addr_234_6, addr_positional[3755:3752], addr_938_7);

wire[31:0] addr_939_7;

Selector_2 s939_7(wires_234_6[3], addr_234_6, addr_positional[3759:3756], addr_939_7);

wire[31:0] addr_940_7;

Selector_2 s940_7(wires_235_6[0], addr_235_6, addr_positional[3763:3760], addr_940_7);

wire[31:0] addr_941_7;

Selector_2 s941_7(wires_235_6[1], addr_235_6, addr_positional[3767:3764], addr_941_7);

wire[31:0] addr_942_7;

Selector_2 s942_7(wires_235_6[2], addr_235_6, addr_positional[3771:3768], addr_942_7);

wire[31:0] addr_943_7;

Selector_2 s943_7(wires_235_6[3], addr_235_6, addr_positional[3775:3772], addr_943_7);

wire[31:0] addr_944_7;

Selector_2 s944_7(wires_236_6[0], addr_236_6, addr_positional[3779:3776], addr_944_7);

wire[31:0] addr_945_7;

Selector_2 s945_7(wires_236_6[1], addr_236_6, addr_positional[3783:3780], addr_945_7);

wire[31:0] addr_946_7;

Selector_2 s946_7(wires_236_6[2], addr_236_6, addr_positional[3787:3784], addr_946_7);

wire[31:0] addr_947_7;

Selector_2 s947_7(wires_236_6[3], addr_236_6, addr_positional[3791:3788], addr_947_7);

wire[31:0] addr_948_7;

Selector_2 s948_7(wires_237_6[0], addr_237_6, addr_positional[3795:3792], addr_948_7);

wire[31:0] addr_949_7;

Selector_2 s949_7(wires_237_6[1], addr_237_6, addr_positional[3799:3796], addr_949_7);

wire[31:0] addr_950_7;

Selector_2 s950_7(wires_237_6[2], addr_237_6, addr_positional[3803:3800], addr_950_7);

wire[31:0] addr_951_7;

Selector_2 s951_7(wires_237_6[3], addr_237_6, addr_positional[3807:3804], addr_951_7);

wire[31:0] addr_952_7;

Selector_2 s952_7(wires_238_6[0], addr_238_6, addr_positional[3811:3808], addr_952_7);

wire[31:0] addr_953_7;

Selector_2 s953_7(wires_238_6[1], addr_238_6, addr_positional[3815:3812], addr_953_7);

wire[31:0] addr_954_7;

Selector_2 s954_7(wires_238_6[2], addr_238_6, addr_positional[3819:3816], addr_954_7);

wire[31:0] addr_955_7;

Selector_2 s955_7(wires_238_6[3], addr_238_6, addr_positional[3823:3820], addr_955_7);

wire[31:0] addr_956_7;

Selector_2 s956_7(wires_239_6[0], addr_239_6, addr_positional[3827:3824], addr_956_7);

wire[31:0] addr_957_7;

Selector_2 s957_7(wires_239_6[1], addr_239_6, addr_positional[3831:3828], addr_957_7);

wire[31:0] addr_958_7;

Selector_2 s958_7(wires_239_6[2], addr_239_6, addr_positional[3835:3832], addr_958_7);

wire[31:0] addr_959_7;

Selector_2 s959_7(wires_239_6[3], addr_239_6, addr_positional[3839:3836], addr_959_7);

wire[31:0] addr_960_7;

Selector_2 s960_7(wires_240_6[0], addr_240_6, addr_positional[3843:3840], addr_960_7);

wire[31:0] addr_961_7;

Selector_2 s961_7(wires_240_6[1], addr_240_6, addr_positional[3847:3844], addr_961_7);

wire[31:0] addr_962_7;

Selector_2 s962_7(wires_240_6[2], addr_240_6, addr_positional[3851:3848], addr_962_7);

wire[31:0] addr_963_7;

Selector_2 s963_7(wires_240_6[3], addr_240_6, addr_positional[3855:3852], addr_963_7);

wire[31:0] addr_964_7;

Selector_2 s964_7(wires_241_6[0], addr_241_6, addr_positional[3859:3856], addr_964_7);

wire[31:0] addr_965_7;

Selector_2 s965_7(wires_241_6[1], addr_241_6, addr_positional[3863:3860], addr_965_7);

wire[31:0] addr_966_7;

Selector_2 s966_7(wires_241_6[2], addr_241_6, addr_positional[3867:3864], addr_966_7);

wire[31:0] addr_967_7;

Selector_2 s967_7(wires_241_6[3], addr_241_6, addr_positional[3871:3868], addr_967_7);

wire[31:0] addr_968_7;

Selector_2 s968_7(wires_242_6[0], addr_242_6, addr_positional[3875:3872], addr_968_7);

wire[31:0] addr_969_7;

Selector_2 s969_7(wires_242_6[1], addr_242_6, addr_positional[3879:3876], addr_969_7);

wire[31:0] addr_970_7;

Selector_2 s970_7(wires_242_6[2], addr_242_6, addr_positional[3883:3880], addr_970_7);

wire[31:0] addr_971_7;

Selector_2 s971_7(wires_242_6[3], addr_242_6, addr_positional[3887:3884], addr_971_7);

wire[31:0] addr_972_7;

Selector_2 s972_7(wires_243_6[0], addr_243_6, addr_positional[3891:3888], addr_972_7);

wire[31:0] addr_973_7;

Selector_2 s973_7(wires_243_6[1], addr_243_6, addr_positional[3895:3892], addr_973_7);

wire[31:0] addr_974_7;

Selector_2 s974_7(wires_243_6[2], addr_243_6, addr_positional[3899:3896], addr_974_7);

wire[31:0] addr_975_7;

Selector_2 s975_7(wires_243_6[3], addr_243_6, addr_positional[3903:3900], addr_975_7);

wire[31:0] addr_976_7;

Selector_2 s976_7(wires_244_6[0], addr_244_6, addr_positional[3907:3904], addr_976_7);

wire[31:0] addr_977_7;

Selector_2 s977_7(wires_244_6[1], addr_244_6, addr_positional[3911:3908], addr_977_7);

wire[31:0] addr_978_7;

Selector_2 s978_7(wires_244_6[2], addr_244_6, addr_positional[3915:3912], addr_978_7);

wire[31:0] addr_979_7;

Selector_2 s979_7(wires_244_6[3], addr_244_6, addr_positional[3919:3916], addr_979_7);

wire[31:0] addr_980_7;

Selector_2 s980_7(wires_245_6[0], addr_245_6, addr_positional[3923:3920], addr_980_7);

wire[31:0] addr_981_7;

Selector_2 s981_7(wires_245_6[1], addr_245_6, addr_positional[3927:3924], addr_981_7);

wire[31:0] addr_982_7;

Selector_2 s982_7(wires_245_6[2], addr_245_6, addr_positional[3931:3928], addr_982_7);

wire[31:0] addr_983_7;

Selector_2 s983_7(wires_245_6[3], addr_245_6, addr_positional[3935:3932], addr_983_7);

wire[31:0] addr_984_7;

Selector_2 s984_7(wires_246_6[0], addr_246_6, addr_positional[3939:3936], addr_984_7);

wire[31:0] addr_985_7;

Selector_2 s985_7(wires_246_6[1], addr_246_6, addr_positional[3943:3940], addr_985_7);

wire[31:0] addr_986_7;

Selector_2 s986_7(wires_246_6[2], addr_246_6, addr_positional[3947:3944], addr_986_7);

wire[31:0] addr_987_7;

Selector_2 s987_7(wires_246_6[3], addr_246_6, addr_positional[3951:3948], addr_987_7);

wire[31:0] addr_988_7;

Selector_2 s988_7(wires_247_6[0], addr_247_6, addr_positional[3955:3952], addr_988_7);

wire[31:0] addr_989_7;

Selector_2 s989_7(wires_247_6[1], addr_247_6, addr_positional[3959:3956], addr_989_7);

wire[31:0] addr_990_7;

Selector_2 s990_7(wires_247_6[2], addr_247_6, addr_positional[3963:3960], addr_990_7);

wire[31:0] addr_991_7;

Selector_2 s991_7(wires_247_6[3], addr_247_6, addr_positional[3967:3964], addr_991_7);

wire[31:0] addr_992_7;

Selector_2 s992_7(wires_248_6[0], addr_248_6, addr_positional[3971:3968], addr_992_7);

wire[31:0] addr_993_7;

Selector_2 s993_7(wires_248_6[1], addr_248_6, addr_positional[3975:3972], addr_993_7);

wire[31:0] addr_994_7;

Selector_2 s994_7(wires_248_6[2], addr_248_6, addr_positional[3979:3976], addr_994_7);

wire[31:0] addr_995_7;

Selector_2 s995_7(wires_248_6[3], addr_248_6, addr_positional[3983:3980], addr_995_7);

wire[31:0] addr_996_7;

Selector_2 s996_7(wires_249_6[0], addr_249_6, addr_positional[3987:3984], addr_996_7);

wire[31:0] addr_997_7;

Selector_2 s997_7(wires_249_6[1], addr_249_6, addr_positional[3991:3988], addr_997_7);

wire[31:0] addr_998_7;

Selector_2 s998_7(wires_249_6[2], addr_249_6, addr_positional[3995:3992], addr_998_7);

wire[31:0] addr_999_7;

Selector_2 s999_7(wires_249_6[3], addr_249_6, addr_positional[3999:3996], addr_999_7);

wire[31:0] addr_1000_7;

Selector_2 s1000_7(wires_250_6[0], addr_250_6, addr_positional[4003:4000], addr_1000_7);

wire[31:0] addr_1001_7;

Selector_2 s1001_7(wires_250_6[1], addr_250_6, addr_positional[4007:4004], addr_1001_7);

wire[31:0] addr_1002_7;

Selector_2 s1002_7(wires_250_6[2], addr_250_6, addr_positional[4011:4008], addr_1002_7);

wire[31:0] addr_1003_7;

Selector_2 s1003_7(wires_250_6[3], addr_250_6, addr_positional[4015:4012], addr_1003_7);

wire[31:0] addr_1004_7;

Selector_2 s1004_7(wires_251_6[0], addr_251_6, addr_positional[4019:4016], addr_1004_7);

wire[31:0] addr_1005_7;

Selector_2 s1005_7(wires_251_6[1], addr_251_6, addr_positional[4023:4020], addr_1005_7);

wire[31:0] addr_1006_7;

Selector_2 s1006_7(wires_251_6[2], addr_251_6, addr_positional[4027:4024], addr_1006_7);

wire[31:0] addr_1007_7;

Selector_2 s1007_7(wires_251_6[3], addr_251_6, addr_positional[4031:4028], addr_1007_7);

wire[31:0] addr_1008_7;

Selector_2 s1008_7(wires_252_6[0], addr_252_6, addr_positional[4035:4032], addr_1008_7);

wire[31:0] addr_1009_7;

Selector_2 s1009_7(wires_252_6[1], addr_252_6, addr_positional[4039:4036], addr_1009_7);

wire[31:0] addr_1010_7;

Selector_2 s1010_7(wires_252_6[2], addr_252_6, addr_positional[4043:4040], addr_1010_7);

wire[31:0] addr_1011_7;

Selector_2 s1011_7(wires_252_6[3], addr_252_6, addr_positional[4047:4044], addr_1011_7);

wire[31:0] addr_1012_7;

Selector_2 s1012_7(wires_253_6[0], addr_253_6, addr_positional[4051:4048], addr_1012_7);

wire[31:0] addr_1013_7;

Selector_2 s1013_7(wires_253_6[1], addr_253_6, addr_positional[4055:4052], addr_1013_7);

wire[31:0] addr_1014_7;

Selector_2 s1014_7(wires_253_6[2], addr_253_6, addr_positional[4059:4056], addr_1014_7);

wire[31:0] addr_1015_7;

Selector_2 s1015_7(wires_253_6[3], addr_253_6, addr_positional[4063:4060], addr_1015_7);

wire[31:0] addr_1016_7;

Selector_2 s1016_7(wires_254_6[0], addr_254_6, addr_positional[4067:4064], addr_1016_7);

wire[31:0] addr_1017_7;

Selector_2 s1017_7(wires_254_6[1], addr_254_6, addr_positional[4071:4068], addr_1017_7);

wire[31:0] addr_1018_7;

Selector_2 s1018_7(wires_254_6[2], addr_254_6, addr_positional[4075:4072], addr_1018_7);

wire[31:0] addr_1019_7;

Selector_2 s1019_7(wires_254_6[3], addr_254_6, addr_positional[4079:4076], addr_1019_7);

wire[31:0] addr_1020_7;

Selector_2 s1020_7(wires_255_6[0], addr_255_6, addr_positional[4083:4080], addr_1020_7);

wire[31:0] addr_1021_7;

Selector_2 s1021_7(wires_255_6[1], addr_255_6, addr_positional[4087:4084], addr_1021_7);

wire[31:0] addr_1022_7;

Selector_2 s1022_7(wires_255_6[2], addr_255_6, addr_positional[4091:4088], addr_1022_7);

wire[31:0] addr_1023_7;

Selector_2 s1023_7(wires_255_6[3], addr_255_6, addr_positional[4095:4092], addr_1023_7);

wire[31:0] addr_1024_7;

Selector_2 s1024_7(wires_256_6[0], addr_256_6, addr_positional[4099:4096], addr_1024_7);

wire[31:0] addr_1025_7;

Selector_2 s1025_7(wires_256_6[1], addr_256_6, addr_positional[4103:4100], addr_1025_7);

wire[31:0] addr_1026_7;

Selector_2 s1026_7(wires_256_6[2], addr_256_6, addr_positional[4107:4104], addr_1026_7);

wire[31:0] addr_1027_7;

Selector_2 s1027_7(wires_256_6[3], addr_256_6, addr_positional[4111:4108], addr_1027_7);

wire[31:0] addr_1028_7;

Selector_2 s1028_7(wires_257_6[0], addr_257_6, addr_positional[4115:4112], addr_1028_7);

wire[31:0] addr_1029_7;

Selector_2 s1029_7(wires_257_6[1], addr_257_6, addr_positional[4119:4116], addr_1029_7);

wire[31:0] addr_1030_7;

Selector_2 s1030_7(wires_257_6[2], addr_257_6, addr_positional[4123:4120], addr_1030_7);

wire[31:0] addr_1031_7;

Selector_2 s1031_7(wires_257_6[3], addr_257_6, addr_positional[4127:4124], addr_1031_7);

wire[31:0] addr_1032_7;

Selector_2 s1032_7(wires_258_6[0], addr_258_6, addr_positional[4131:4128], addr_1032_7);

wire[31:0] addr_1033_7;

Selector_2 s1033_7(wires_258_6[1], addr_258_6, addr_positional[4135:4132], addr_1033_7);

wire[31:0] addr_1034_7;

Selector_2 s1034_7(wires_258_6[2], addr_258_6, addr_positional[4139:4136], addr_1034_7);

wire[31:0] addr_1035_7;

Selector_2 s1035_7(wires_258_6[3], addr_258_6, addr_positional[4143:4140], addr_1035_7);

wire[31:0] addr_1036_7;

Selector_2 s1036_7(wires_259_6[0], addr_259_6, addr_positional[4147:4144], addr_1036_7);

wire[31:0] addr_1037_7;

Selector_2 s1037_7(wires_259_6[1], addr_259_6, addr_positional[4151:4148], addr_1037_7);

wire[31:0] addr_1038_7;

Selector_2 s1038_7(wires_259_6[2], addr_259_6, addr_positional[4155:4152], addr_1038_7);

wire[31:0] addr_1039_7;

Selector_2 s1039_7(wires_259_6[3], addr_259_6, addr_positional[4159:4156], addr_1039_7);

wire[31:0] addr_1040_7;

Selector_2 s1040_7(wires_260_6[0], addr_260_6, addr_positional[4163:4160], addr_1040_7);

wire[31:0] addr_1041_7;

Selector_2 s1041_7(wires_260_6[1], addr_260_6, addr_positional[4167:4164], addr_1041_7);

wire[31:0] addr_1042_7;

Selector_2 s1042_7(wires_260_6[2], addr_260_6, addr_positional[4171:4168], addr_1042_7);

wire[31:0] addr_1043_7;

Selector_2 s1043_7(wires_260_6[3], addr_260_6, addr_positional[4175:4172], addr_1043_7);

wire[31:0] addr_1044_7;

Selector_2 s1044_7(wires_261_6[0], addr_261_6, addr_positional[4179:4176], addr_1044_7);

wire[31:0] addr_1045_7;

Selector_2 s1045_7(wires_261_6[1], addr_261_6, addr_positional[4183:4180], addr_1045_7);

wire[31:0] addr_1046_7;

Selector_2 s1046_7(wires_261_6[2], addr_261_6, addr_positional[4187:4184], addr_1046_7);

wire[31:0] addr_1047_7;

Selector_2 s1047_7(wires_261_6[3], addr_261_6, addr_positional[4191:4188], addr_1047_7);

wire[31:0] addr_1048_7;

Selector_2 s1048_7(wires_262_6[0], addr_262_6, addr_positional[4195:4192], addr_1048_7);

wire[31:0] addr_1049_7;

Selector_2 s1049_7(wires_262_6[1], addr_262_6, addr_positional[4199:4196], addr_1049_7);

wire[31:0] addr_1050_7;

Selector_2 s1050_7(wires_262_6[2], addr_262_6, addr_positional[4203:4200], addr_1050_7);

wire[31:0] addr_1051_7;

Selector_2 s1051_7(wires_262_6[3], addr_262_6, addr_positional[4207:4204], addr_1051_7);

wire[31:0] addr_1052_7;

Selector_2 s1052_7(wires_263_6[0], addr_263_6, addr_positional[4211:4208], addr_1052_7);

wire[31:0] addr_1053_7;

Selector_2 s1053_7(wires_263_6[1], addr_263_6, addr_positional[4215:4212], addr_1053_7);

wire[31:0] addr_1054_7;

Selector_2 s1054_7(wires_263_6[2], addr_263_6, addr_positional[4219:4216], addr_1054_7);

wire[31:0] addr_1055_7;

Selector_2 s1055_7(wires_263_6[3], addr_263_6, addr_positional[4223:4220], addr_1055_7);

wire[31:0] addr_1056_7;

Selector_2 s1056_7(wires_264_6[0], addr_264_6, addr_positional[4227:4224], addr_1056_7);

wire[31:0] addr_1057_7;

Selector_2 s1057_7(wires_264_6[1], addr_264_6, addr_positional[4231:4228], addr_1057_7);

wire[31:0] addr_1058_7;

Selector_2 s1058_7(wires_264_6[2], addr_264_6, addr_positional[4235:4232], addr_1058_7);

wire[31:0] addr_1059_7;

Selector_2 s1059_7(wires_264_6[3], addr_264_6, addr_positional[4239:4236], addr_1059_7);

wire[31:0] addr_1060_7;

Selector_2 s1060_7(wires_265_6[0], addr_265_6, addr_positional[4243:4240], addr_1060_7);

wire[31:0] addr_1061_7;

Selector_2 s1061_7(wires_265_6[1], addr_265_6, addr_positional[4247:4244], addr_1061_7);

wire[31:0] addr_1062_7;

Selector_2 s1062_7(wires_265_6[2], addr_265_6, addr_positional[4251:4248], addr_1062_7);

wire[31:0] addr_1063_7;

Selector_2 s1063_7(wires_265_6[3], addr_265_6, addr_positional[4255:4252], addr_1063_7);

wire[31:0] addr_1064_7;

Selector_2 s1064_7(wires_266_6[0], addr_266_6, addr_positional[4259:4256], addr_1064_7);

wire[31:0] addr_1065_7;

Selector_2 s1065_7(wires_266_6[1], addr_266_6, addr_positional[4263:4260], addr_1065_7);

wire[31:0] addr_1066_7;

Selector_2 s1066_7(wires_266_6[2], addr_266_6, addr_positional[4267:4264], addr_1066_7);

wire[31:0] addr_1067_7;

Selector_2 s1067_7(wires_266_6[3], addr_266_6, addr_positional[4271:4268], addr_1067_7);

wire[31:0] addr_1068_7;

Selector_2 s1068_7(wires_267_6[0], addr_267_6, addr_positional[4275:4272], addr_1068_7);

wire[31:0] addr_1069_7;

Selector_2 s1069_7(wires_267_6[1], addr_267_6, addr_positional[4279:4276], addr_1069_7);

wire[31:0] addr_1070_7;

Selector_2 s1070_7(wires_267_6[2], addr_267_6, addr_positional[4283:4280], addr_1070_7);

wire[31:0] addr_1071_7;

Selector_2 s1071_7(wires_267_6[3], addr_267_6, addr_positional[4287:4284], addr_1071_7);

wire[31:0] addr_1072_7;

Selector_2 s1072_7(wires_268_6[0], addr_268_6, addr_positional[4291:4288], addr_1072_7);

wire[31:0] addr_1073_7;

Selector_2 s1073_7(wires_268_6[1], addr_268_6, addr_positional[4295:4292], addr_1073_7);

wire[31:0] addr_1074_7;

Selector_2 s1074_7(wires_268_6[2], addr_268_6, addr_positional[4299:4296], addr_1074_7);

wire[31:0] addr_1075_7;

Selector_2 s1075_7(wires_268_6[3], addr_268_6, addr_positional[4303:4300], addr_1075_7);

wire[31:0] addr_1076_7;

Selector_2 s1076_7(wires_269_6[0], addr_269_6, addr_positional[4307:4304], addr_1076_7);

wire[31:0] addr_1077_7;

Selector_2 s1077_7(wires_269_6[1], addr_269_6, addr_positional[4311:4308], addr_1077_7);

wire[31:0] addr_1078_7;

Selector_2 s1078_7(wires_269_6[2], addr_269_6, addr_positional[4315:4312], addr_1078_7);

wire[31:0] addr_1079_7;

Selector_2 s1079_7(wires_269_6[3], addr_269_6, addr_positional[4319:4316], addr_1079_7);

wire[31:0] addr_1080_7;

Selector_2 s1080_7(wires_270_6[0], addr_270_6, addr_positional[4323:4320], addr_1080_7);

wire[31:0] addr_1081_7;

Selector_2 s1081_7(wires_270_6[1], addr_270_6, addr_positional[4327:4324], addr_1081_7);

wire[31:0] addr_1082_7;

Selector_2 s1082_7(wires_270_6[2], addr_270_6, addr_positional[4331:4328], addr_1082_7);

wire[31:0] addr_1083_7;

Selector_2 s1083_7(wires_270_6[3], addr_270_6, addr_positional[4335:4332], addr_1083_7);

wire[31:0] addr_1084_7;

Selector_2 s1084_7(wires_271_6[0], addr_271_6, addr_positional[4339:4336], addr_1084_7);

wire[31:0] addr_1085_7;

Selector_2 s1085_7(wires_271_6[1], addr_271_6, addr_positional[4343:4340], addr_1085_7);

wire[31:0] addr_1086_7;

Selector_2 s1086_7(wires_271_6[2], addr_271_6, addr_positional[4347:4344], addr_1086_7);

wire[31:0] addr_1087_7;

Selector_2 s1087_7(wires_271_6[3], addr_271_6, addr_positional[4351:4348], addr_1087_7);

wire[31:0] addr_1088_7;

Selector_2 s1088_7(wires_272_6[0], addr_272_6, addr_positional[4355:4352], addr_1088_7);

wire[31:0] addr_1089_7;

Selector_2 s1089_7(wires_272_6[1], addr_272_6, addr_positional[4359:4356], addr_1089_7);

wire[31:0] addr_1090_7;

Selector_2 s1090_7(wires_272_6[2], addr_272_6, addr_positional[4363:4360], addr_1090_7);

wire[31:0] addr_1091_7;

Selector_2 s1091_7(wires_272_6[3], addr_272_6, addr_positional[4367:4364], addr_1091_7);

wire[31:0] addr_1092_7;

Selector_2 s1092_7(wires_273_6[0], addr_273_6, addr_positional[4371:4368], addr_1092_7);

wire[31:0] addr_1093_7;

Selector_2 s1093_7(wires_273_6[1], addr_273_6, addr_positional[4375:4372], addr_1093_7);

wire[31:0] addr_1094_7;

Selector_2 s1094_7(wires_273_6[2], addr_273_6, addr_positional[4379:4376], addr_1094_7);

wire[31:0] addr_1095_7;

Selector_2 s1095_7(wires_273_6[3], addr_273_6, addr_positional[4383:4380], addr_1095_7);

wire[31:0] addr_1096_7;

Selector_2 s1096_7(wires_274_6[0], addr_274_6, addr_positional[4387:4384], addr_1096_7);

wire[31:0] addr_1097_7;

Selector_2 s1097_7(wires_274_6[1], addr_274_6, addr_positional[4391:4388], addr_1097_7);

wire[31:0] addr_1098_7;

Selector_2 s1098_7(wires_274_6[2], addr_274_6, addr_positional[4395:4392], addr_1098_7);

wire[31:0] addr_1099_7;

Selector_2 s1099_7(wires_274_6[3], addr_274_6, addr_positional[4399:4396], addr_1099_7);

wire[31:0] addr_1100_7;

Selector_2 s1100_7(wires_275_6[0], addr_275_6, addr_positional[4403:4400], addr_1100_7);

wire[31:0] addr_1101_7;

Selector_2 s1101_7(wires_275_6[1], addr_275_6, addr_positional[4407:4404], addr_1101_7);

wire[31:0] addr_1102_7;

Selector_2 s1102_7(wires_275_6[2], addr_275_6, addr_positional[4411:4408], addr_1102_7);

wire[31:0] addr_1103_7;

Selector_2 s1103_7(wires_275_6[3], addr_275_6, addr_positional[4415:4412], addr_1103_7);

wire[31:0] addr_1104_7;

Selector_2 s1104_7(wires_276_6[0], addr_276_6, addr_positional[4419:4416], addr_1104_7);

wire[31:0] addr_1105_7;

Selector_2 s1105_7(wires_276_6[1], addr_276_6, addr_positional[4423:4420], addr_1105_7);

wire[31:0] addr_1106_7;

Selector_2 s1106_7(wires_276_6[2], addr_276_6, addr_positional[4427:4424], addr_1106_7);

wire[31:0] addr_1107_7;

Selector_2 s1107_7(wires_276_6[3], addr_276_6, addr_positional[4431:4428], addr_1107_7);

wire[31:0] addr_1108_7;

Selector_2 s1108_7(wires_277_6[0], addr_277_6, addr_positional[4435:4432], addr_1108_7);

wire[31:0] addr_1109_7;

Selector_2 s1109_7(wires_277_6[1], addr_277_6, addr_positional[4439:4436], addr_1109_7);

wire[31:0] addr_1110_7;

Selector_2 s1110_7(wires_277_6[2], addr_277_6, addr_positional[4443:4440], addr_1110_7);

wire[31:0] addr_1111_7;

Selector_2 s1111_7(wires_277_6[3], addr_277_6, addr_positional[4447:4444], addr_1111_7);

wire[31:0] addr_1112_7;

Selector_2 s1112_7(wires_278_6[0], addr_278_6, addr_positional[4451:4448], addr_1112_7);

wire[31:0] addr_1113_7;

Selector_2 s1113_7(wires_278_6[1], addr_278_6, addr_positional[4455:4452], addr_1113_7);

wire[31:0] addr_1114_7;

Selector_2 s1114_7(wires_278_6[2], addr_278_6, addr_positional[4459:4456], addr_1114_7);

wire[31:0] addr_1115_7;

Selector_2 s1115_7(wires_278_6[3], addr_278_6, addr_positional[4463:4460], addr_1115_7);

wire[31:0] addr_1116_7;

Selector_2 s1116_7(wires_279_6[0], addr_279_6, addr_positional[4467:4464], addr_1116_7);

wire[31:0] addr_1117_7;

Selector_2 s1117_7(wires_279_6[1], addr_279_6, addr_positional[4471:4468], addr_1117_7);

wire[31:0] addr_1118_7;

Selector_2 s1118_7(wires_279_6[2], addr_279_6, addr_positional[4475:4472], addr_1118_7);

wire[31:0] addr_1119_7;

Selector_2 s1119_7(wires_279_6[3], addr_279_6, addr_positional[4479:4476], addr_1119_7);

wire[31:0] addr_1120_7;

Selector_2 s1120_7(wires_280_6[0], addr_280_6, addr_positional[4483:4480], addr_1120_7);

wire[31:0] addr_1121_7;

Selector_2 s1121_7(wires_280_6[1], addr_280_6, addr_positional[4487:4484], addr_1121_7);

wire[31:0] addr_1122_7;

Selector_2 s1122_7(wires_280_6[2], addr_280_6, addr_positional[4491:4488], addr_1122_7);

wire[31:0] addr_1123_7;

Selector_2 s1123_7(wires_280_6[3], addr_280_6, addr_positional[4495:4492], addr_1123_7);

wire[31:0] addr_1124_7;

Selector_2 s1124_7(wires_281_6[0], addr_281_6, addr_positional[4499:4496], addr_1124_7);

wire[31:0] addr_1125_7;

Selector_2 s1125_7(wires_281_6[1], addr_281_6, addr_positional[4503:4500], addr_1125_7);

wire[31:0] addr_1126_7;

Selector_2 s1126_7(wires_281_6[2], addr_281_6, addr_positional[4507:4504], addr_1126_7);

wire[31:0] addr_1127_7;

Selector_2 s1127_7(wires_281_6[3], addr_281_6, addr_positional[4511:4508], addr_1127_7);

wire[31:0] addr_1128_7;

Selector_2 s1128_7(wires_282_6[0], addr_282_6, addr_positional[4515:4512], addr_1128_7);

wire[31:0] addr_1129_7;

Selector_2 s1129_7(wires_282_6[1], addr_282_6, addr_positional[4519:4516], addr_1129_7);

wire[31:0] addr_1130_7;

Selector_2 s1130_7(wires_282_6[2], addr_282_6, addr_positional[4523:4520], addr_1130_7);

wire[31:0] addr_1131_7;

Selector_2 s1131_7(wires_282_6[3], addr_282_6, addr_positional[4527:4524], addr_1131_7);

wire[31:0] addr_1132_7;

Selector_2 s1132_7(wires_283_6[0], addr_283_6, addr_positional[4531:4528], addr_1132_7);

wire[31:0] addr_1133_7;

Selector_2 s1133_7(wires_283_6[1], addr_283_6, addr_positional[4535:4532], addr_1133_7);

wire[31:0] addr_1134_7;

Selector_2 s1134_7(wires_283_6[2], addr_283_6, addr_positional[4539:4536], addr_1134_7);

wire[31:0] addr_1135_7;

Selector_2 s1135_7(wires_283_6[3], addr_283_6, addr_positional[4543:4540], addr_1135_7);

wire[31:0] addr_1136_7;

Selector_2 s1136_7(wires_284_6[0], addr_284_6, addr_positional[4547:4544], addr_1136_7);

wire[31:0] addr_1137_7;

Selector_2 s1137_7(wires_284_6[1], addr_284_6, addr_positional[4551:4548], addr_1137_7);

wire[31:0] addr_1138_7;

Selector_2 s1138_7(wires_284_6[2], addr_284_6, addr_positional[4555:4552], addr_1138_7);

wire[31:0] addr_1139_7;

Selector_2 s1139_7(wires_284_6[3], addr_284_6, addr_positional[4559:4556], addr_1139_7);

wire[31:0] addr_1140_7;

Selector_2 s1140_7(wires_285_6[0], addr_285_6, addr_positional[4563:4560], addr_1140_7);

wire[31:0] addr_1141_7;

Selector_2 s1141_7(wires_285_6[1], addr_285_6, addr_positional[4567:4564], addr_1141_7);

wire[31:0] addr_1142_7;

Selector_2 s1142_7(wires_285_6[2], addr_285_6, addr_positional[4571:4568], addr_1142_7);

wire[31:0] addr_1143_7;

Selector_2 s1143_7(wires_285_6[3], addr_285_6, addr_positional[4575:4572], addr_1143_7);

wire[31:0] addr_1144_7;

Selector_2 s1144_7(wires_286_6[0], addr_286_6, addr_positional[4579:4576], addr_1144_7);

wire[31:0] addr_1145_7;

Selector_2 s1145_7(wires_286_6[1], addr_286_6, addr_positional[4583:4580], addr_1145_7);

wire[31:0] addr_1146_7;

Selector_2 s1146_7(wires_286_6[2], addr_286_6, addr_positional[4587:4584], addr_1146_7);

wire[31:0] addr_1147_7;

Selector_2 s1147_7(wires_286_6[3], addr_286_6, addr_positional[4591:4588], addr_1147_7);

wire[31:0] addr_1148_7;

Selector_2 s1148_7(wires_287_6[0], addr_287_6, addr_positional[4595:4592], addr_1148_7);

wire[31:0] addr_1149_7;

Selector_2 s1149_7(wires_287_6[1], addr_287_6, addr_positional[4599:4596], addr_1149_7);

wire[31:0] addr_1150_7;

Selector_2 s1150_7(wires_287_6[2], addr_287_6, addr_positional[4603:4600], addr_1150_7);

wire[31:0] addr_1151_7;

Selector_2 s1151_7(wires_287_6[3], addr_287_6, addr_positional[4607:4604], addr_1151_7);

wire[31:0] addr_1152_7;

Selector_2 s1152_7(wires_288_6[0], addr_288_6, addr_positional[4611:4608], addr_1152_7);

wire[31:0] addr_1153_7;

Selector_2 s1153_7(wires_288_6[1], addr_288_6, addr_positional[4615:4612], addr_1153_7);

wire[31:0] addr_1154_7;

Selector_2 s1154_7(wires_288_6[2], addr_288_6, addr_positional[4619:4616], addr_1154_7);

wire[31:0] addr_1155_7;

Selector_2 s1155_7(wires_288_6[3], addr_288_6, addr_positional[4623:4620], addr_1155_7);

wire[31:0] addr_1156_7;

Selector_2 s1156_7(wires_289_6[0], addr_289_6, addr_positional[4627:4624], addr_1156_7);

wire[31:0] addr_1157_7;

Selector_2 s1157_7(wires_289_6[1], addr_289_6, addr_positional[4631:4628], addr_1157_7);

wire[31:0] addr_1158_7;

Selector_2 s1158_7(wires_289_6[2], addr_289_6, addr_positional[4635:4632], addr_1158_7);

wire[31:0] addr_1159_7;

Selector_2 s1159_7(wires_289_6[3], addr_289_6, addr_positional[4639:4636], addr_1159_7);

wire[31:0] addr_1160_7;

Selector_2 s1160_7(wires_290_6[0], addr_290_6, addr_positional[4643:4640], addr_1160_7);

wire[31:0] addr_1161_7;

Selector_2 s1161_7(wires_290_6[1], addr_290_6, addr_positional[4647:4644], addr_1161_7);

wire[31:0] addr_1162_7;

Selector_2 s1162_7(wires_290_6[2], addr_290_6, addr_positional[4651:4648], addr_1162_7);

wire[31:0] addr_1163_7;

Selector_2 s1163_7(wires_290_6[3], addr_290_6, addr_positional[4655:4652], addr_1163_7);

wire[31:0] addr_1164_7;

Selector_2 s1164_7(wires_291_6[0], addr_291_6, addr_positional[4659:4656], addr_1164_7);

wire[31:0] addr_1165_7;

Selector_2 s1165_7(wires_291_6[1], addr_291_6, addr_positional[4663:4660], addr_1165_7);

wire[31:0] addr_1166_7;

Selector_2 s1166_7(wires_291_6[2], addr_291_6, addr_positional[4667:4664], addr_1166_7);

wire[31:0] addr_1167_7;

Selector_2 s1167_7(wires_291_6[3], addr_291_6, addr_positional[4671:4668], addr_1167_7);

wire[31:0] addr_1168_7;

Selector_2 s1168_7(wires_292_6[0], addr_292_6, addr_positional[4675:4672], addr_1168_7);

wire[31:0] addr_1169_7;

Selector_2 s1169_7(wires_292_6[1], addr_292_6, addr_positional[4679:4676], addr_1169_7);

wire[31:0] addr_1170_7;

Selector_2 s1170_7(wires_292_6[2], addr_292_6, addr_positional[4683:4680], addr_1170_7);

wire[31:0] addr_1171_7;

Selector_2 s1171_7(wires_292_6[3], addr_292_6, addr_positional[4687:4684], addr_1171_7);

wire[31:0] addr_1172_7;

Selector_2 s1172_7(wires_293_6[0], addr_293_6, addr_positional[4691:4688], addr_1172_7);

wire[31:0] addr_1173_7;

Selector_2 s1173_7(wires_293_6[1], addr_293_6, addr_positional[4695:4692], addr_1173_7);

wire[31:0] addr_1174_7;

Selector_2 s1174_7(wires_293_6[2], addr_293_6, addr_positional[4699:4696], addr_1174_7);

wire[31:0] addr_1175_7;

Selector_2 s1175_7(wires_293_6[3], addr_293_6, addr_positional[4703:4700], addr_1175_7);

wire[31:0] addr_1176_7;

Selector_2 s1176_7(wires_294_6[0], addr_294_6, addr_positional[4707:4704], addr_1176_7);

wire[31:0] addr_1177_7;

Selector_2 s1177_7(wires_294_6[1], addr_294_6, addr_positional[4711:4708], addr_1177_7);

wire[31:0] addr_1178_7;

Selector_2 s1178_7(wires_294_6[2], addr_294_6, addr_positional[4715:4712], addr_1178_7);

wire[31:0] addr_1179_7;

Selector_2 s1179_7(wires_294_6[3], addr_294_6, addr_positional[4719:4716], addr_1179_7);

wire[31:0] addr_1180_7;

Selector_2 s1180_7(wires_295_6[0], addr_295_6, addr_positional[4723:4720], addr_1180_7);

wire[31:0] addr_1181_7;

Selector_2 s1181_7(wires_295_6[1], addr_295_6, addr_positional[4727:4724], addr_1181_7);

wire[31:0] addr_1182_7;

Selector_2 s1182_7(wires_295_6[2], addr_295_6, addr_positional[4731:4728], addr_1182_7);

wire[31:0] addr_1183_7;

Selector_2 s1183_7(wires_295_6[3], addr_295_6, addr_positional[4735:4732], addr_1183_7);

wire[31:0] addr_1184_7;

Selector_2 s1184_7(wires_296_6[0], addr_296_6, addr_positional[4739:4736], addr_1184_7);

wire[31:0] addr_1185_7;

Selector_2 s1185_7(wires_296_6[1], addr_296_6, addr_positional[4743:4740], addr_1185_7);

wire[31:0] addr_1186_7;

Selector_2 s1186_7(wires_296_6[2], addr_296_6, addr_positional[4747:4744], addr_1186_7);

wire[31:0] addr_1187_7;

Selector_2 s1187_7(wires_296_6[3], addr_296_6, addr_positional[4751:4748], addr_1187_7);

wire[31:0] addr_1188_7;

Selector_2 s1188_7(wires_297_6[0], addr_297_6, addr_positional[4755:4752], addr_1188_7);

wire[31:0] addr_1189_7;

Selector_2 s1189_7(wires_297_6[1], addr_297_6, addr_positional[4759:4756], addr_1189_7);

wire[31:0] addr_1190_7;

Selector_2 s1190_7(wires_297_6[2], addr_297_6, addr_positional[4763:4760], addr_1190_7);

wire[31:0] addr_1191_7;

Selector_2 s1191_7(wires_297_6[3], addr_297_6, addr_positional[4767:4764], addr_1191_7);

wire[31:0] addr_1192_7;

Selector_2 s1192_7(wires_298_6[0], addr_298_6, addr_positional[4771:4768], addr_1192_7);

wire[31:0] addr_1193_7;

Selector_2 s1193_7(wires_298_6[1], addr_298_6, addr_positional[4775:4772], addr_1193_7);

wire[31:0] addr_1194_7;

Selector_2 s1194_7(wires_298_6[2], addr_298_6, addr_positional[4779:4776], addr_1194_7);

wire[31:0] addr_1195_7;

Selector_2 s1195_7(wires_298_6[3], addr_298_6, addr_positional[4783:4780], addr_1195_7);

wire[31:0] addr_1196_7;

Selector_2 s1196_7(wires_299_6[0], addr_299_6, addr_positional[4787:4784], addr_1196_7);

wire[31:0] addr_1197_7;

Selector_2 s1197_7(wires_299_6[1], addr_299_6, addr_positional[4791:4788], addr_1197_7);

wire[31:0] addr_1198_7;

Selector_2 s1198_7(wires_299_6[2], addr_299_6, addr_positional[4795:4792], addr_1198_7);

wire[31:0] addr_1199_7;

Selector_2 s1199_7(wires_299_6[3], addr_299_6, addr_positional[4799:4796], addr_1199_7);

wire[31:0] addr_1200_7;

Selector_2 s1200_7(wires_300_6[0], addr_300_6, addr_positional[4803:4800], addr_1200_7);

wire[31:0] addr_1201_7;

Selector_2 s1201_7(wires_300_6[1], addr_300_6, addr_positional[4807:4804], addr_1201_7);

wire[31:0] addr_1202_7;

Selector_2 s1202_7(wires_300_6[2], addr_300_6, addr_positional[4811:4808], addr_1202_7);

wire[31:0] addr_1203_7;

Selector_2 s1203_7(wires_300_6[3], addr_300_6, addr_positional[4815:4812], addr_1203_7);

wire[31:0] addr_1204_7;

Selector_2 s1204_7(wires_301_6[0], addr_301_6, addr_positional[4819:4816], addr_1204_7);

wire[31:0] addr_1205_7;

Selector_2 s1205_7(wires_301_6[1], addr_301_6, addr_positional[4823:4820], addr_1205_7);

wire[31:0] addr_1206_7;

Selector_2 s1206_7(wires_301_6[2], addr_301_6, addr_positional[4827:4824], addr_1206_7);

wire[31:0] addr_1207_7;

Selector_2 s1207_7(wires_301_6[3], addr_301_6, addr_positional[4831:4828], addr_1207_7);

wire[31:0] addr_1208_7;

Selector_2 s1208_7(wires_302_6[0], addr_302_6, addr_positional[4835:4832], addr_1208_7);

wire[31:0] addr_1209_7;

Selector_2 s1209_7(wires_302_6[1], addr_302_6, addr_positional[4839:4836], addr_1209_7);

wire[31:0] addr_1210_7;

Selector_2 s1210_7(wires_302_6[2], addr_302_6, addr_positional[4843:4840], addr_1210_7);

wire[31:0] addr_1211_7;

Selector_2 s1211_7(wires_302_6[3], addr_302_6, addr_positional[4847:4844], addr_1211_7);

wire[31:0] addr_1212_7;

Selector_2 s1212_7(wires_303_6[0], addr_303_6, addr_positional[4851:4848], addr_1212_7);

wire[31:0] addr_1213_7;

Selector_2 s1213_7(wires_303_6[1], addr_303_6, addr_positional[4855:4852], addr_1213_7);

wire[31:0] addr_1214_7;

Selector_2 s1214_7(wires_303_6[2], addr_303_6, addr_positional[4859:4856], addr_1214_7);

wire[31:0] addr_1215_7;

Selector_2 s1215_7(wires_303_6[3], addr_303_6, addr_positional[4863:4860], addr_1215_7);

wire[31:0] addr_1216_7;

Selector_2 s1216_7(wires_304_6[0], addr_304_6, addr_positional[4867:4864], addr_1216_7);

wire[31:0] addr_1217_7;

Selector_2 s1217_7(wires_304_6[1], addr_304_6, addr_positional[4871:4868], addr_1217_7);

wire[31:0] addr_1218_7;

Selector_2 s1218_7(wires_304_6[2], addr_304_6, addr_positional[4875:4872], addr_1218_7);

wire[31:0] addr_1219_7;

Selector_2 s1219_7(wires_304_6[3], addr_304_6, addr_positional[4879:4876], addr_1219_7);

wire[31:0] addr_1220_7;

Selector_2 s1220_7(wires_305_6[0], addr_305_6, addr_positional[4883:4880], addr_1220_7);

wire[31:0] addr_1221_7;

Selector_2 s1221_7(wires_305_6[1], addr_305_6, addr_positional[4887:4884], addr_1221_7);

wire[31:0] addr_1222_7;

Selector_2 s1222_7(wires_305_6[2], addr_305_6, addr_positional[4891:4888], addr_1222_7);

wire[31:0] addr_1223_7;

Selector_2 s1223_7(wires_305_6[3], addr_305_6, addr_positional[4895:4892], addr_1223_7);

wire[31:0] addr_1224_7;

Selector_2 s1224_7(wires_306_6[0], addr_306_6, addr_positional[4899:4896], addr_1224_7);

wire[31:0] addr_1225_7;

Selector_2 s1225_7(wires_306_6[1], addr_306_6, addr_positional[4903:4900], addr_1225_7);

wire[31:0] addr_1226_7;

Selector_2 s1226_7(wires_306_6[2], addr_306_6, addr_positional[4907:4904], addr_1226_7);

wire[31:0] addr_1227_7;

Selector_2 s1227_7(wires_306_6[3], addr_306_6, addr_positional[4911:4908], addr_1227_7);

wire[31:0] addr_1228_7;

Selector_2 s1228_7(wires_307_6[0], addr_307_6, addr_positional[4915:4912], addr_1228_7);

wire[31:0] addr_1229_7;

Selector_2 s1229_7(wires_307_6[1], addr_307_6, addr_positional[4919:4916], addr_1229_7);

wire[31:0] addr_1230_7;

Selector_2 s1230_7(wires_307_6[2], addr_307_6, addr_positional[4923:4920], addr_1230_7);

wire[31:0] addr_1231_7;

Selector_2 s1231_7(wires_307_6[3], addr_307_6, addr_positional[4927:4924], addr_1231_7);

wire[31:0] addr_1232_7;

Selector_2 s1232_7(wires_308_6[0], addr_308_6, addr_positional[4931:4928], addr_1232_7);

wire[31:0] addr_1233_7;

Selector_2 s1233_7(wires_308_6[1], addr_308_6, addr_positional[4935:4932], addr_1233_7);

wire[31:0] addr_1234_7;

Selector_2 s1234_7(wires_308_6[2], addr_308_6, addr_positional[4939:4936], addr_1234_7);

wire[31:0] addr_1235_7;

Selector_2 s1235_7(wires_308_6[3], addr_308_6, addr_positional[4943:4940], addr_1235_7);

wire[31:0] addr_1236_7;

Selector_2 s1236_7(wires_309_6[0], addr_309_6, addr_positional[4947:4944], addr_1236_7);

wire[31:0] addr_1237_7;

Selector_2 s1237_7(wires_309_6[1], addr_309_6, addr_positional[4951:4948], addr_1237_7);

wire[31:0] addr_1238_7;

Selector_2 s1238_7(wires_309_6[2], addr_309_6, addr_positional[4955:4952], addr_1238_7);

wire[31:0] addr_1239_7;

Selector_2 s1239_7(wires_309_6[3], addr_309_6, addr_positional[4959:4956], addr_1239_7);

wire[31:0] addr_1240_7;

Selector_2 s1240_7(wires_310_6[0], addr_310_6, addr_positional[4963:4960], addr_1240_7);

wire[31:0] addr_1241_7;

Selector_2 s1241_7(wires_310_6[1], addr_310_6, addr_positional[4967:4964], addr_1241_7);

wire[31:0] addr_1242_7;

Selector_2 s1242_7(wires_310_6[2], addr_310_6, addr_positional[4971:4968], addr_1242_7);

wire[31:0] addr_1243_7;

Selector_2 s1243_7(wires_310_6[3], addr_310_6, addr_positional[4975:4972], addr_1243_7);

wire[31:0] addr_1244_7;

Selector_2 s1244_7(wires_311_6[0], addr_311_6, addr_positional[4979:4976], addr_1244_7);

wire[31:0] addr_1245_7;

Selector_2 s1245_7(wires_311_6[1], addr_311_6, addr_positional[4983:4980], addr_1245_7);

wire[31:0] addr_1246_7;

Selector_2 s1246_7(wires_311_6[2], addr_311_6, addr_positional[4987:4984], addr_1246_7);

wire[31:0] addr_1247_7;

Selector_2 s1247_7(wires_311_6[3], addr_311_6, addr_positional[4991:4988], addr_1247_7);

wire[31:0] addr_1248_7;

Selector_2 s1248_7(wires_312_6[0], addr_312_6, addr_positional[4995:4992], addr_1248_7);

wire[31:0] addr_1249_7;

Selector_2 s1249_7(wires_312_6[1], addr_312_6, addr_positional[4999:4996], addr_1249_7);

wire[31:0] addr_1250_7;

Selector_2 s1250_7(wires_312_6[2], addr_312_6, addr_positional[5003:5000], addr_1250_7);

wire[31:0] addr_1251_7;

Selector_2 s1251_7(wires_312_6[3], addr_312_6, addr_positional[5007:5004], addr_1251_7);

wire[31:0] addr_1252_7;

Selector_2 s1252_7(wires_313_6[0], addr_313_6, addr_positional[5011:5008], addr_1252_7);

wire[31:0] addr_1253_7;

Selector_2 s1253_7(wires_313_6[1], addr_313_6, addr_positional[5015:5012], addr_1253_7);

wire[31:0] addr_1254_7;

Selector_2 s1254_7(wires_313_6[2], addr_313_6, addr_positional[5019:5016], addr_1254_7);

wire[31:0] addr_1255_7;

Selector_2 s1255_7(wires_313_6[3], addr_313_6, addr_positional[5023:5020], addr_1255_7);

wire[31:0] addr_1256_7;

Selector_2 s1256_7(wires_314_6[0], addr_314_6, addr_positional[5027:5024], addr_1256_7);

wire[31:0] addr_1257_7;

Selector_2 s1257_7(wires_314_6[1], addr_314_6, addr_positional[5031:5028], addr_1257_7);

wire[31:0] addr_1258_7;

Selector_2 s1258_7(wires_314_6[2], addr_314_6, addr_positional[5035:5032], addr_1258_7);

wire[31:0] addr_1259_7;

Selector_2 s1259_7(wires_314_6[3], addr_314_6, addr_positional[5039:5036], addr_1259_7);

wire[31:0] addr_1260_7;

Selector_2 s1260_7(wires_315_6[0], addr_315_6, addr_positional[5043:5040], addr_1260_7);

wire[31:0] addr_1261_7;

Selector_2 s1261_7(wires_315_6[1], addr_315_6, addr_positional[5047:5044], addr_1261_7);

wire[31:0] addr_1262_7;

Selector_2 s1262_7(wires_315_6[2], addr_315_6, addr_positional[5051:5048], addr_1262_7);

wire[31:0] addr_1263_7;

Selector_2 s1263_7(wires_315_6[3], addr_315_6, addr_positional[5055:5052], addr_1263_7);

wire[31:0] addr_1264_7;

Selector_2 s1264_7(wires_316_6[0], addr_316_6, addr_positional[5059:5056], addr_1264_7);

wire[31:0] addr_1265_7;

Selector_2 s1265_7(wires_316_6[1], addr_316_6, addr_positional[5063:5060], addr_1265_7);

wire[31:0] addr_1266_7;

Selector_2 s1266_7(wires_316_6[2], addr_316_6, addr_positional[5067:5064], addr_1266_7);

wire[31:0] addr_1267_7;

Selector_2 s1267_7(wires_316_6[3], addr_316_6, addr_positional[5071:5068], addr_1267_7);

wire[31:0] addr_1268_7;

Selector_2 s1268_7(wires_317_6[0], addr_317_6, addr_positional[5075:5072], addr_1268_7);

wire[31:0] addr_1269_7;

Selector_2 s1269_7(wires_317_6[1], addr_317_6, addr_positional[5079:5076], addr_1269_7);

wire[31:0] addr_1270_7;

Selector_2 s1270_7(wires_317_6[2], addr_317_6, addr_positional[5083:5080], addr_1270_7);

wire[31:0] addr_1271_7;

Selector_2 s1271_7(wires_317_6[3], addr_317_6, addr_positional[5087:5084], addr_1271_7);

wire[31:0] addr_1272_7;

Selector_2 s1272_7(wires_318_6[0], addr_318_6, addr_positional[5091:5088], addr_1272_7);

wire[31:0] addr_1273_7;

Selector_2 s1273_7(wires_318_6[1], addr_318_6, addr_positional[5095:5092], addr_1273_7);

wire[31:0] addr_1274_7;

Selector_2 s1274_7(wires_318_6[2], addr_318_6, addr_positional[5099:5096], addr_1274_7);

wire[31:0] addr_1275_7;

Selector_2 s1275_7(wires_318_6[3], addr_318_6, addr_positional[5103:5100], addr_1275_7);

wire[31:0] addr_1276_7;

Selector_2 s1276_7(wires_319_6[0], addr_319_6, addr_positional[5107:5104], addr_1276_7);

wire[31:0] addr_1277_7;

Selector_2 s1277_7(wires_319_6[1], addr_319_6, addr_positional[5111:5108], addr_1277_7);

wire[31:0] addr_1278_7;

Selector_2 s1278_7(wires_319_6[2], addr_319_6, addr_positional[5115:5112], addr_1278_7);

wire[31:0] addr_1279_7;

Selector_2 s1279_7(wires_319_6[3], addr_319_6, addr_positional[5119:5116], addr_1279_7);

wire[31:0] addr_1280_7;

Selector_2 s1280_7(wires_320_6[0], addr_320_6, addr_positional[5123:5120], addr_1280_7);

wire[31:0] addr_1281_7;

Selector_2 s1281_7(wires_320_6[1], addr_320_6, addr_positional[5127:5124], addr_1281_7);

wire[31:0] addr_1282_7;

Selector_2 s1282_7(wires_320_6[2], addr_320_6, addr_positional[5131:5128], addr_1282_7);

wire[31:0] addr_1283_7;

Selector_2 s1283_7(wires_320_6[3], addr_320_6, addr_positional[5135:5132], addr_1283_7);

wire[31:0] addr_1284_7;

Selector_2 s1284_7(wires_321_6[0], addr_321_6, addr_positional[5139:5136], addr_1284_7);

wire[31:0] addr_1285_7;

Selector_2 s1285_7(wires_321_6[1], addr_321_6, addr_positional[5143:5140], addr_1285_7);

wire[31:0] addr_1286_7;

Selector_2 s1286_7(wires_321_6[2], addr_321_6, addr_positional[5147:5144], addr_1286_7);

wire[31:0] addr_1287_7;

Selector_2 s1287_7(wires_321_6[3], addr_321_6, addr_positional[5151:5148], addr_1287_7);

wire[31:0] addr_1288_7;

Selector_2 s1288_7(wires_322_6[0], addr_322_6, addr_positional[5155:5152], addr_1288_7);

wire[31:0] addr_1289_7;

Selector_2 s1289_7(wires_322_6[1], addr_322_6, addr_positional[5159:5156], addr_1289_7);

wire[31:0] addr_1290_7;

Selector_2 s1290_7(wires_322_6[2], addr_322_6, addr_positional[5163:5160], addr_1290_7);

wire[31:0] addr_1291_7;

Selector_2 s1291_7(wires_322_6[3], addr_322_6, addr_positional[5167:5164], addr_1291_7);

wire[31:0] addr_1292_7;

Selector_2 s1292_7(wires_323_6[0], addr_323_6, addr_positional[5171:5168], addr_1292_7);

wire[31:0] addr_1293_7;

Selector_2 s1293_7(wires_323_6[1], addr_323_6, addr_positional[5175:5172], addr_1293_7);

wire[31:0] addr_1294_7;

Selector_2 s1294_7(wires_323_6[2], addr_323_6, addr_positional[5179:5176], addr_1294_7);

wire[31:0] addr_1295_7;

Selector_2 s1295_7(wires_323_6[3], addr_323_6, addr_positional[5183:5180], addr_1295_7);

wire[31:0] addr_1296_7;

Selector_2 s1296_7(wires_324_6[0], addr_324_6, addr_positional[5187:5184], addr_1296_7);

wire[31:0] addr_1297_7;

Selector_2 s1297_7(wires_324_6[1], addr_324_6, addr_positional[5191:5188], addr_1297_7);

wire[31:0] addr_1298_7;

Selector_2 s1298_7(wires_324_6[2], addr_324_6, addr_positional[5195:5192], addr_1298_7);

wire[31:0] addr_1299_7;

Selector_2 s1299_7(wires_324_6[3], addr_324_6, addr_positional[5199:5196], addr_1299_7);

wire[31:0] addr_1300_7;

Selector_2 s1300_7(wires_325_6[0], addr_325_6, addr_positional[5203:5200], addr_1300_7);

wire[31:0] addr_1301_7;

Selector_2 s1301_7(wires_325_6[1], addr_325_6, addr_positional[5207:5204], addr_1301_7);

wire[31:0] addr_1302_7;

Selector_2 s1302_7(wires_325_6[2], addr_325_6, addr_positional[5211:5208], addr_1302_7);

wire[31:0] addr_1303_7;

Selector_2 s1303_7(wires_325_6[3], addr_325_6, addr_positional[5215:5212], addr_1303_7);

wire[31:0] addr_1304_7;

Selector_2 s1304_7(wires_326_6[0], addr_326_6, addr_positional[5219:5216], addr_1304_7);

wire[31:0] addr_1305_7;

Selector_2 s1305_7(wires_326_6[1], addr_326_6, addr_positional[5223:5220], addr_1305_7);

wire[31:0] addr_1306_7;

Selector_2 s1306_7(wires_326_6[2], addr_326_6, addr_positional[5227:5224], addr_1306_7);

wire[31:0] addr_1307_7;

Selector_2 s1307_7(wires_326_6[3], addr_326_6, addr_positional[5231:5228], addr_1307_7);

wire[31:0] addr_1308_7;

Selector_2 s1308_7(wires_327_6[0], addr_327_6, addr_positional[5235:5232], addr_1308_7);

wire[31:0] addr_1309_7;

Selector_2 s1309_7(wires_327_6[1], addr_327_6, addr_positional[5239:5236], addr_1309_7);

wire[31:0] addr_1310_7;

Selector_2 s1310_7(wires_327_6[2], addr_327_6, addr_positional[5243:5240], addr_1310_7);

wire[31:0] addr_1311_7;

Selector_2 s1311_7(wires_327_6[3], addr_327_6, addr_positional[5247:5244], addr_1311_7);

wire[31:0] addr_1312_7;

Selector_2 s1312_7(wires_328_6[0], addr_328_6, addr_positional[5251:5248], addr_1312_7);

wire[31:0] addr_1313_7;

Selector_2 s1313_7(wires_328_6[1], addr_328_6, addr_positional[5255:5252], addr_1313_7);

wire[31:0] addr_1314_7;

Selector_2 s1314_7(wires_328_6[2], addr_328_6, addr_positional[5259:5256], addr_1314_7);

wire[31:0] addr_1315_7;

Selector_2 s1315_7(wires_328_6[3], addr_328_6, addr_positional[5263:5260], addr_1315_7);

wire[31:0] addr_1316_7;

Selector_2 s1316_7(wires_329_6[0], addr_329_6, addr_positional[5267:5264], addr_1316_7);

wire[31:0] addr_1317_7;

Selector_2 s1317_7(wires_329_6[1], addr_329_6, addr_positional[5271:5268], addr_1317_7);

wire[31:0] addr_1318_7;

Selector_2 s1318_7(wires_329_6[2], addr_329_6, addr_positional[5275:5272], addr_1318_7);

wire[31:0] addr_1319_7;

Selector_2 s1319_7(wires_329_6[3], addr_329_6, addr_positional[5279:5276], addr_1319_7);

wire[31:0] addr_1320_7;

Selector_2 s1320_7(wires_330_6[0], addr_330_6, addr_positional[5283:5280], addr_1320_7);

wire[31:0] addr_1321_7;

Selector_2 s1321_7(wires_330_6[1], addr_330_6, addr_positional[5287:5284], addr_1321_7);

wire[31:0] addr_1322_7;

Selector_2 s1322_7(wires_330_6[2], addr_330_6, addr_positional[5291:5288], addr_1322_7);

wire[31:0] addr_1323_7;

Selector_2 s1323_7(wires_330_6[3], addr_330_6, addr_positional[5295:5292], addr_1323_7);

wire[31:0] addr_1324_7;

Selector_2 s1324_7(wires_331_6[0], addr_331_6, addr_positional[5299:5296], addr_1324_7);

wire[31:0] addr_1325_7;

Selector_2 s1325_7(wires_331_6[1], addr_331_6, addr_positional[5303:5300], addr_1325_7);

wire[31:0] addr_1326_7;

Selector_2 s1326_7(wires_331_6[2], addr_331_6, addr_positional[5307:5304], addr_1326_7);

wire[31:0] addr_1327_7;

Selector_2 s1327_7(wires_331_6[3], addr_331_6, addr_positional[5311:5308], addr_1327_7);

wire[31:0] addr_1328_7;

Selector_2 s1328_7(wires_332_6[0], addr_332_6, addr_positional[5315:5312], addr_1328_7);

wire[31:0] addr_1329_7;

Selector_2 s1329_7(wires_332_6[1], addr_332_6, addr_positional[5319:5316], addr_1329_7);

wire[31:0] addr_1330_7;

Selector_2 s1330_7(wires_332_6[2], addr_332_6, addr_positional[5323:5320], addr_1330_7);

wire[31:0] addr_1331_7;

Selector_2 s1331_7(wires_332_6[3], addr_332_6, addr_positional[5327:5324], addr_1331_7);

wire[31:0] addr_1332_7;

Selector_2 s1332_7(wires_333_6[0], addr_333_6, addr_positional[5331:5328], addr_1332_7);

wire[31:0] addr_1333_7;

Selector_2 s1333_7(wires_333_6[1], addr_333_6, addr_positional[5335:5332], addr_1333_7);

wire[31:0] addr_1334_7;

Selector_2 s1334_7(wires_333_6[2], addr_333_6, addr_positional[5339:5336], addr_1334_7);

wire[31:0] addr_1335_7;

Selector_2 s1335_7(wires_333_6[3], addr_333_6, addr_positional[5343:5340], addr_1335_7);

wire[31:0] addr_1336_7;

Selector_2 s1336_7(wires_334_6[0], addr_334_6, addr_positional[5347:5344], addr_1336_7);

wire[31:0] addr_1337_7;

Selector_2 s1337_7(wires_334_6[1], addr_334_6, addr_positional[5351:5348], addr_1337_7);

wire[31:0] addr_1338_7;

Selector_2 s1338_7(wires_334_6[2], addr_334_6, addr_positional[5355:5352], addr_1338_7);

wire[31:0] addr_1339_7;

Selector_2 s1339_7(wires_334_6[3], addr_334_6, addr_positional[5359:5356], addr_1339_7);

wire[31:0] addr_1340_7;

Selector_2 s1340_7(wires_335_6[0], addr_335_6, addr_positional[5363:5360], addr_1340_7);

wire[31:0] addr_1341_7;

Selector_2 s1341_7(wires_335_6[1], addr_335_6, addr_positional[5367:5364], addr_1341_7);

wire[31:0] addr_1342_7;

Selector_2 s1342_7(wires_335_6[2], addr_335_6, addr_positional[5371:5368], addr_1342_7);

wire[31:0] addr_1343_7;

Selector_2 s1343_7(wires_335_6[3], addr_335_6, addr_positional[5375:5372], addr_1343_7);

wire[31:0] addr_1344_7;

Selector_2 s1344_7(wires_336_6[0], addr_336_6, addr_positional[5379:5376], addr_1344_7);

wire[31:0] addr_1345_7;

Selector_2 s1345_7(wires_336_6[1], addr_336_6, addr_positional[5383:5380], addr_1345_7);

wire[31:0] addr_1346_7;

Selector_2 s1346_7(wires_336_6[2], addr_336_6, addr_positional[5387:5384], addr_1346_7);

wire[31:0] addr_1347_7;

Selector_2 s1347_7(wires_336_6[3], addr_336_6, addr_positional[5391:5388], addr_1347_7);

wire[31:0] addr_1348_7;

Selector_2 s1348_7(wires_337_6[0], addr_337_6, addr_positional[5395:5392], addr_1348_7);

wire[31:0] addr_1349_7;

Selector_2 s1349_7(wires_337_6[1], addr_337_6, addr_positional[5399:5396], addr_1349_7);

wire[31:0] addr_1350_7;

Selector_2 s1350_7(wires_337_6[2], addr_337_6, addr_positional[5403:5400], addr_1350_7);

wire[31:0] addr_1351_7;

Selector_2 s1351_7(wires_337_6[3], addr_337_6, addr_positional[5407:5404], addr_1351_7);

wire[31:0] addr_1352_7;

Selector_2 s1352_7(wires_338_6[0], addr_338_6, addr_positional[5411:5408], addr_1352_7);

wire[31:0] addr_1353_7;

Selector_2 s1353_7(wires_338_6[1], addr_338_6, addr_positional[5415:5412], addr_1353_7);

wire[31:0] addr_1354_7;

Selector_2 s1354_7(wires_338_6[2], addr_338_6, addr_positional[5419:5416], addr_1354_7);

wire[31:0] addr_1355_7;

Selector_2 s1355_7(wires_338_6[3], addr_338_6, addr_positional[5423:5420], addr_1355_7);

wire[31:0] addr_1356_7;

Selector_2 s1356_7(wires_339_6[0], addr_339_6, addr_positional[5427:5424], addr_1356_7);

wire[31:0] addr_1357_7;

Selector_2 s1357_7(wires_339_6[1], addr_339_6, addr_positional[5431:5428], addr_1357_7);

wire[31:0] addr_1358_7;

Selector_2 s1358_7(wires_339_6[2], addr_339_6, addr_positional[5435:5432], addr_1358_7);

wire[31:0] addr_1359_7;

Selector_2 s1359_7(wires_339_6[3], addr_339_6, addr_positional[5439:5436], addr_1359_7);

wire[31:0] addr_1360_7;

Selector_2 s1360_7(wires_340_6[0], addr_340_6, addr_positional[5443:5440], addr_1360_7);

wire[31:0] addr_1361_7;

Selector_2 s1361_7(wires_340_6[1], addr_340_6, addr_positional[5447:5444], addr_1361_7);

wire[31:0] addr_1362_7;

Selector_2 s1362_7(wires_340_6[2], addr_340_6, addr_positional[5451:5448], addr_1362_7);

wire[31:0] addr_1363_7;

Selector_2 s1363_7(wires_340_6[3], addr_340_6, addr_positional[5455:5452], addr_1363_7);

wire[31:0] addr_1364_7;

Selector_2 s1364_7(wires_341_6[0], addr_341_6, addr_positional[5459:5456], addr_1364_7);

wire[31:0] addr_1365_7;

Selector_2 s1365_7(wires_341_6[1], addr_341_6, addr_positional[5463:5460], addr_1365_7);

wire[31:0] addr_1366_7;

Selector_2 s1366_7(wires_341_6[2], addr_341_6, addr_positional[5467:5464], addr_1366_7);

wire[31:0] addr_1367_7;

Selector_2 s1367_7(wires_341_6[3], addr_341_6, addr_positional[5471:5468], addr_1367_7);

wire[31:0] addr_1368_7;

Selector_2 s1368_7(wires_342_6[0], addr_342_6, addr_positional[5475:5472], addr_1368_7);

wire[31:0] addr_1369_7;

Selector_2 s1369_7(wires_342_6[1], addr_342_6, addr_positional[5479:5476], addr_1369_7);

wire[31:0] addr_1370_7;

Selector_2 s1370_7(wires_342_6[2], addr_342_6, addr_positional[5483:5480], addr_1370_7);

wire[31:0] addr_1371_7;

Selector_2 s1371_7(wires_342_6[3], addr_342_6, addr_positional[5487:5484], addr_1371_7);

wire[31:0] addr_1372_7;

Selector_2 s1372_7(wires_343_6[0], addr_343_6, addr_positional[5491:5488], addr_1372_7);

wire[31:0] addr_1373_7;

Selector_2 s1373_7(wires_343_6[1], addr_343_6, addr_positional[5495:5492], addr_1373_7);

wire[31:0] addr_1374_7;

Selector_2 s1374_7(wires_343_6[2], addr_343_6, addr_positional[5499:5496], addr_1374_7);

wire[31:0] addr_1375_7;

Selector_2 s1375_7(wires_343_6[3], addr_343_6, addr_positional[5503:5500], addr_1375_7);

wire[31:0] addr_1376_7;

Selector_2 s1376_7(wires_344_6[0], addr_344_6, addr_positional[5507:5504], addr_1376_7);

wire[31:0] addr_1377_7;

Selector_2 s1377_7(wires_344_6[1], addr_344_6, addr_positional[5511:5508], addr_1377_7);

wire[31:0] addr_1378_7;

Selector_2 s1378_7(wires_344_6[2], addr_344_6, addr_positional[5515:5512], addr_1378_7);

wire[31:0] addr_1379_7;

Selector_2 s1379_7(wires_344_6[3], addr_344_6, addr_positional[5519:5516], addr_1379_7);

wire[31:0] addr_1380_7;

Selector_2 s1380_7(wires_345_6[0], addr_345_6, addr_positional[5523:5520], addr_1380_7);

wire[31:0] addr_1381_7;

Selector_2 s1381_7(wires_345_6[1], addr_345_6, addr_positional[5527:5524], addr_1381_7);

wire[31:0] addr_1382_7;

Selector_2 s1382_7(wires_345_6[2], addr_345_6, addr_positional[5531:5528], addr_1382_7);

wire[31:0] addr_1383_7;

Selector_2 s1383_7(wires_345_6[3], addr_345_6, addr_positional[5535:5532], addr_1383_7);

wire[31:0] addr_1384_7;

Selector_2 s1384_7(wires_346_6[0], addr_346_6, addr_positional[5539:5536], addr_1384_7);

wire[31:0] addr_1385_7;

Selector_2 s1385_7(wires_346_6[1], addr_346_6, addr_positional[5543:5540], addr_1385_7);

wire[31:0] addr_1386_7;

Selector_2 s1386_7(wires_346_6[2], addr_346_6, addr_positional[5547:5544], addr_1386_7);

wire[31:0] addr_1387_7;

Selector_2 s1387_7(wires_346_6[3], addr_346_6, addr_positional[5551:5548], addr_1387_7);

wire[31:0] addr_1388_7;

Selector_2 s1388_7(wires_347_6[0], addr_347_6, addr_positional[5555:5552], addr_1388_7);

wire[31:0] addr_1389_7;

Selector_2 s1389_7(wires_347_6[1], addr_347_6, addr_positional[5559:5556], addr_1389_7);

wire[31:0] addr_1390_7;

Selector_2 s1390_7(wires_347_6[2], addr_347_6, addr_positional[5563:5560], addr_1390_7);

wire[31:0] addr_1391_7;

Selector_2 s1391_7(wires_347_6[3], addr_347_6, addr_positional[5567:5564], addr_1391_7);

wire[31:0] addr_1392_7;

Selector_2 s1392_7(wires_348_6[0], addr_348_6, addr_positional[5571:5568], addr_1392_7);

wire[31:0] addr_1393_7;

Selector_2 s1393_7(wires_348_6[1], addr_348_6, addr_positional[5575:5572], addr_1393_7);

wire[31:0] addr_1394_7;

Selector_2 s1394_7(wires_348_6[2], addr_348_6, addr_positional[5579:5576], addr_1394_7);

wire[31:0] addr_1395_7;

Selector_2 s1395_7(wires_348_6[3], addr_348_6, addr_positional[5583:5580], addr_1395_7);

wire[31:0] addr_1396_7;

Selector_2 s1396_7(wires_349_6[0], addr_349_6, addr_positional[5587:5584], addr_1396_7);

wire[31:0] addr_1397_7;

Selector_2 s1397_7(wires_349_6[1], addr_349_6, addr_positional[5591:5588], addr_1397_7);

wire[31:0] addr_1398_7;

Selector_2 s1398_7(wires_349_6[2], addr_349_6, addr_positional[5595:5592], addr_1398_7);

wire[31:0] addr_1399_7;

Selector_2 s1399_7(wires_349_6[3], addr_349_6, addr_positional[5599:5596], addr_1399_7);

wire[31:0] addr_1400_7;

Selector_2 s1400_7(wires_350_6[0], addr_350_6, addr_positional[5603:5600], addr_1400_7);

wire[31:0] addr_1401_7;

Selector_2 s1401_7(wires_350_6[1], addr_350_6, addr_positional[5607:5604], addr_1401_7);

wire[31:0] addr_1402_7;

Selector_2 s1402_7(wires_350_6[2], addr_350_6, addr_positional[5611:5608], addr_1402_7);

wire[31:0] addr_1403_7;

Selector_2 s1403_7(wires_350_6[3], addr_350_6, addr_positional[5615:5612], addr_1403_7);

wire[31:0] addr_1404_7;

Selector_2 s1404_7(wires_351_6[0], addr_351_6, addr_positional[5619:5616], addr_1404_7);

wire[31:0] addr_1405_7;

Selector_2 s1405_7(wires_351_6[1], addr_351_6, addr_positional[5623:5620], addr_1405_7);

wire[31:0] addr_1406_7;

Selector_2 s1406_7(wires_351_6[2], addr_351_6, addr_positional[5627:5624], addr_1406_7);

wire[31:0] addr_1407_7;

Selector_2 s1407_7(wires_351_6[3], addr_351_6, addr_positional[5631:5628], addr_1407_7);

wire[31:0] addr_1408_7;

Selector_2 s1408_7(wires_352_6[0], addr_352_6, addr_positional[5635:5632], addr_1408_7);

wire[31:0] addr_1409_7;

Selector_2 s1409_7(wires_352_6[1], addr_352_6, addr_positional[5639:5636], addr_1409_7);

wire[31:0] addr_1410_7;

Selector_2 s1410_7(wires_352_6[2], addr_352_6, addr_positional[5643:5640], addr_1410_7);

wire[31:0] addr_1411_7;

Selector_2 s1411_7(wires_352_6[3], addr_352_6, addr_positional[5647:5644], addr_1411_7);

wire[31:0] addr_1412_7;

Selector_2 s1412_7(wires_353_6[0], addr_353_6, addr_positional[5651:5648], addr_1412_7);

wire[31:0] addr_1413_7;

Selector_2 s1413_7(wires_353_6[1], addr_353_6, addr_positional[5655:5652], addr_1413_7);

wire[31:0] addr_1414_7;

Selector_2 s1414_7(wires_353_6[2], addr_353_6, addr_positional[5659:5656], addr_1414_7);

wire[31:0] addr_1415_7;

Selector_2 s1415_7(wires_353_6[3], addr_353_6, addr_positional[5663:5660], addr_1415_7);

wire[31:0] addr_1416_7;

Selector_2 s1416_7(wires_354_6[0], addr_354_6, addr_positional[5667:5664], addr_1416_7);

wire[31:0] addr_1417_7;

Selector_2 s1417_7(wires_354_6[1], addr_354_6, addr_positional[5671:5668], addr_1417_7);

wire[31:0] addr_1418_7;

Selector_2 s1418_7(wires_354_6[2], addr_354_6, addr_positional[5675:5672], addr_1418_7);

wire[31:0] addr_1419_7;

Selector_2 s1419_7(wires_354_6[3], addr_354_6, addr_positional[5679:5676], addr_1419_7);

wire[31:0] addr_1420_7;

Selector_2 s1420_7(wires_355_6[0], addr_355_6, addr_positional[5683:5680], addr_1420_7);

wire[31:0] addr_1421_7;

Selector_2 s1421_7(wires_355_6[1], addr_355_6, addr_positional[5687:5684], addr_1421_7);

wire[31:0] addr_1422_7;

Selector_2 s1422_7(wires_355_6[2], addr_355_6, addr_positional[5691:5688], addr_1422_7);

wire[31:0] addr_1423_7;

Selector_2 s1423_7(wires_355_6[3], addr_355_6, addr_positional[5695:5692], addr_1423_7);

wire[31:0] addr_1424_7;

Selector_2 s1424_7(wires_356_6[0], addr_356_6, addr_positional[5699:5696], addr_1424_7);

wire[31:0] addr_1425_7;

Selector_2 s1425_7(wires_356_6[1], addr_356_6, addr_positional[5703:5700], addr_1425_7);

wire[31:0] addr_1426_7;

Selector_2 s1426_7(wires_356_6[2], addr_356_6, addr_positional[5707:5704], addr_1426_7);

wire[31:0] addr_1427_7;

Selector_2 s1427_7(wires_356_6[3], addr_356_6, addr_positional[5711:5708], addr_1427_7);

wire[31:0] addr_1428_7;

Selector_2 s1428_7(wires_357_6[0], addr_357_6, addr_positional[5715:5712], addr_1428_7);

wire[31:0] addr_1429_7;

Selector_2 s1429_7(wires_357_6[1], addr_357_6, addr_positional[5719:5716], addr_1429_7);

wire[31:0] addr_1430_7;

Selector_2 s1430_7(wires_357_6[2], addr_357_6, addr_positional[5723:5720], addr_1430_7);

wire[31:0] addr_1431_7;

Selector_2 s1431_7(wires_357_6[3], addr_357_6, addr_positional[5727:5724], addr_1431_7);

wire[31:0] addr_1432_7;

Selector_2 s1432_7(wires_358_6[0], addr_358_6, addr_positional[5731:5728], addr_1432_7);

wire[31:0] addr_1433_7;

Selector_2 s1433_7(wires_358_6[1], addr_358_6, addr_positional[5735:5732], addr_1433_7);

wire[31:0] addr_1434_7;

Selector_2 s1434_7(wires_358_6[2], addr_358_6, addr_positional[5739:5736], addr_1434_7);

wire[31:0] addr_1435_7;

Selector_2 s1435_7(wires_358_6[3], addr_358_6, addr_positional[5743:5740], addr_1435_7);

wire[31:0] addr_1436_7;

Selector_2 s1436_7(wires_359_6[0], addr_359_6, addr_positional[5747:5744], addr_1436_7);

wire[31:0] addr_1437_7;

Selector_2 s1437_7(wires_359_6[1], addr_359_6, addr_positional[5751:5748], addr_1437_7);

wire[31:0] addr_1438_7;

Selector_2 s1438_7(wires_359_6[2], addr_359_6, addr_positional[5755:5752], addr_1438_7);

wire[31:0] addr_1439_7;

Selector_2 s1439_7(wires_359_6[3], addr_359_6, addr_positional[5759:5756], addr_1439_7);

wire[31:0] addr_1440_7;

Selector_2 s1440_7(wires_360_6[0], addr_360_6, addr_positional[5763:5760], addr_1440_7);

wire[31:0] addr_1441_7;

Selector_2 s1441_7(wires_360_6[1], addr_360_6, addr_positional[5767:5764], addr_1441_7);

wire[31:0] addr_1442_7;

Selector_2 s1442_7(wires_360_6[2], addr_360_6, addr_positional[5771:5768], addr_1442_7);

wire[31:0] addr_1443_7;

Selector_2 s1443_7(wires_360_6[3], addr_360_6, addr_positional[5775:5772], addr_1443_7);

wire[31:0] addr_1444_7;

Selector_2 s1444_7(wires_361_6[0], addr_361_6, addr_positional[5779:5776], addr_1444_7);

wire[31:0] addr_1445_7;

Selector_2 s1445_7(wires_361_6[1], addr_361_6, addr_positional[5783:5780], addr_1445_7);

wire[31:0] addr_1446_7;

Selector_2 s1446_7(wires_361_6[2], addr_361_6, addr_positional[5787:5784], addr_1446_7);

wire[31:0] addr_1447_7;

Selector_2 s1447_7(wires_361_6[3], addr_361_6, addr_positional[5791:5788], addr_1447_7);

wire[31:0] addr_1448_7;

Selector_2 s1448_7(wires_362_6[0], addr_362_6, addr_positional[5795:5792], addr_1448_7);

wire[31:0] addr_1449_7;

Selector_2 s1449_7(wires_362_6[1], addr_362_6, addr_positional[5799:5796], addr_1449_7);

wire[31:0] addr_1450_7;

Selector_2 s1450_7(wires_362_6[2], addr_362_6, addr_positional[5803:5800], addr_1450_7);

wire[31:0] addr_1451_7;

Selector_2 s1451_7(wires_362_6[3], addr_362_6, addr_positional[5807:5804], addr_1451_7);

wire[31:0] addr_1452_7;

Selector_2 s1452_7(wires_363_6[0], addr_363_6, addr_positional[5811:5808], addr_1452_7);

wire[31:0] addr_1453_7;

Selector_2 s1453_7(wires_363_6[1], addr_363_6, addr_positional[5815:5812], addr_1453_7);

wire[31:0] addr_1454_7;

Selector_2 s1454_7(wires_363_6[2], addr_363_6, addr_positional[5819:5816], addr_1454_7);

wire[31:0] addr_1455_7;

Selector_2 s1455_7(wires_363_6[3], addr_363_6, addr_positional[5823:5820], addr_1455_7);

wire[31:0] addr_1456_7;

Selector_2 s1456_7(wires_364_6[0], addr_364_6, addr_positional[5827:5824], addr_1456_7);

wire[31:0] addr_1457_7;

Selector_2 s1457_7(wires_364_6[1], addr_364_6, addr_positional[5831:5828], addr_1457_7);

wire[31:0] addr_1458_7;

Selector_2 s1458_7(wires_364_6[2], addr_364_6, addr_positional[5835:5832], addr_1458_7);

wire[31:0] addr_1459_7;

Selector_2 s1459_7(wires_364_6[3], addr_364_6, addr_positional[5839:5836], addr_1459_7);

wire[31:0] addr_1460_7;

Selector_2 s1460_7(wires_365_6[0], addr_365_6, addr_positional[5843:5840], addr_1460_7);

wire[31:0] addr_1461_7;

Selector_2 s1461_7(wires_365_6[1], addr_365_6, addr_positional[5847:5844], addr_1461_7);

wire[31:0] addr_1462_7;

Selector_2 s1462_7(wires_365_6[2], addr_365_6, addr_positional[5851:5848], addr_1462_7);

wire[31:0] addr_1463_7;

Selector_2 s1463_7(wires_365_6[3], addr_365_6, addr_positional[5855:5852], addr_1463_7);

wire[31:0] addr_1464_7;

Selector_2 s1464_7(wires_366_6[0], addr_366_6, addr_positional[5859:5856], addr_1464_7);

wire[31:0] addr_1465_7;

Selector_2 s1465_7(wires_366_6[1], addr_366_6, addr_positional[5863:5860], addr_1465_7);

wire[31:0] addr_1466_7;

Selector_2 s1466_7(wires_366_6[2], addr_366_6, addr_positional[5867:5864], addr_1466_7);

wire[31:0] addr_1467_7;

Selector_2 s1467_7(wires_366_6[3], addr_366_6, addr_positional[5871:5868], addr_1467_7);

wire[31:0] addr_1468_7;

Selector_2 s1468_7(wires_367_6[0], addr_367_6, addr_positional[5875:5872], addr_1468_7);

wire[31:0] addr_1469_7;

Selector_2 s1469_7(wires_367_6[1], addr_367_6, addr_positional[5879:5876], addr_1469_7);

wire[31:0] addr_1470_7;

Selector_2 s1470_7(wires_367_6[2], addr_367_6, addr_positional[5883:5880], addr_1470_7);

wire[31:0] addr_1471_7;

Selector_2 s1471_7(wires_367_6[3], addr_367_6, addr_positional[5887:5884], addr_1471_7);

wire[31:0] addr_1472_7;

Selector_2 s1472_7(wires_368_6[0], addr_368_6, addr_positional[5891:5888], addr_1472_7);

wire[31:0] addr_1473_7;

Selector_2 s1473_7(wires_368_6[1], addr_368_6, addr_positional[5895:5892], addr_1473_7);

wire[31:0] addr_1474_7;

Selector_2 s1474_7(wires_368_6[2], addr_368_6, addr_positional[5899:5896], addr_1474_7);

wire[31:0] addr_1475_7;

Selector_2 s1475_7(wires_368_6[3], addr_368_6, addr_positional[5903:5900], addr_1475_7);

wire[31:0] addr_1476_7;

Selector_2 s1476_7(wires_369_6[0], addr_369_6, addr_positional[5907:5904], addr_1476_7);

wire[31:0] addr_1477_7;

Selector_2 s1477_7(wires_369_6[1], addr_369_6, addr_positional[5911:5908], addr_1477_7);

wire[31:0] addr_1478_7;

Selector_2 s1478_7(wires_369_6[2], addr_369_6, addr_positional[5915:5912], addr_1478_7);

wire[31:0] addr_1479_7;

Selector_2 s1479_7(wires_369_6[3], addr_369_6, addr_positional[5919:5916], addr_1479_7);

wire[31:0] addr_1480_7;

Selector_2 s1480_7(wires_370_6[0], addr_370_6, addr_positional[5923:5920], addr_1480_7);

wire[31:0] addr_1481_7;

Selector_2 s1481_7(wires_370_6[1], addr_370_6, addr_positional[5927:5924], addr_1481_7);

wire[31:0] addr_1482_7;

Selector_2 s1482_7(wires_370_6[2], addr_370_6, addr_positional[5931:5928], addr_1482_7);

wire[31:0] addr_1483_7;

Selector_2 s1483_7(wires_370_6[3], addr_370_6, addr_positional[5935:5932], addr_1483_7);

wire[31:0] addr_1484_7;

Selector_2 s1484_7(wires_371_6[0], addr_371_6, addr_positional[5939:5936], addr_1484_7);

wire[31:0] addr_1485_7;

Selector_2 s1485_7(wires_371_6[1], addr_371_6, addr_positional[5943:5940], addr_1485_7);

wire[31:0] addr_1486_7;

Selector_2 s1486_7(wires_371_6[2], addr_371_6, addr_positional[5947:5944], addr_1486_7);

wire[31:0] addr_1487_7;

Selector_2 s1487_7(wires_371_6[3], addr_371_6, addr_positional[5951:5948], addr_1487_7);

wire[31:0] addr_1488_7;

Selector_2 s1488_7(wires_372_6[0], addr_372_6, addr_positional[5955:5952], addr_1488_7);

wire[31:0] addr_1489_7;

Selector_2 s1489_7(wires_372_6[1], addr_372_6, addr_positional[5959:5956], addr_1489_7);

wire[31:0] addr_1490_7;

Selector_2 s1490_7(wires_372_6[2], addr_372_6, addr_positional[5963:5960], addr_1490_7);

wire[31:0] addr_1491_7;

Selector_2 s1491_7(wires_372_6[3], addr_372_6, addr_positional[5967:5964], addr_1491_7);

wire[31:0] addr_1492_7;

Selector_2 s1492_7(wires_373_6[0], addr_373_6, addr_positional[5971:5968], addr_1492_7);

wire[31:0] addr_1493_7;

Selector_2 s1493_7(wires_373_6[1], addr_373_6, addr_positional[5975:5972], addr_1493_7);

wire[31:0] addr_1494_7;

Selector_2 s1494_7(wires_373_6[2], addr_373_6, addr_positional[5979:5976], addr_1494_7);

wire[31:0] addr_1495_7;

Selector_2 s1495_7(wires_373_6[3], addr_373_6, addr_positional[5983:5980], addr_1495_7);

wire[31:0] addr_1496_7;

Selector_2 s1496_7(wires_374_6[0], addr_374_6, addr_positional[5987:5984], addr_1496_7);

wire[31:0] addr_1497_7;

Selector_2 s1497_7(wires_374_6[1], addr_374_6, addr_positional[5991:5988], addr_1497_7);

wire[31:0] addr_1498_7;

Selector_2 s1498_7(wires_374_6[2], addr_374_6, addr_positional[5995:5992], addr_1498_7);

wire[31:0] addr_1499_7;

Selector_2 s1499_7(wires_374_6[3], addr_374_6, addr_positional[5999:5996], addr_1499_7);

wire[31:0] addr_1500_7;

Selector_2 s1500_7(wires_375_6[0], addr_375_6, addr_positional[6003:6000], addr_1500_7);

wire[31:0] addr_1501_7;

Selector_2 s1501_7(wires_375_6[1], addr_375_6, addr_positional[6007:6004], addr_1501_7);

wire[31:0] addr_1502_7;

Selector_2 s1502_7(wires_375_6[2], addr_375_6, addr_positional[6011:6008], addr_1502_7);

wire[31:0] addr_1503_7;

Selector_2 s1503_7(wires_375_6[3], addr_375_6, addr_positional[6015:6012], addr_1503_7);

wire[31:0] addr_1504_7;

Selector_2 s1504_7(wires_376_6[0], addr_376_6, addr_positional[6019:6016], addr_1504_7);

wire[31:0] addr_1505_7;

Selector_2 s1505_7(wires_376_6[1], addr_376_6, addr_positional[6023:6020], addr_1505_7);

wire[31:0] addr_1506_7;

Selector_2 s1506_7(wires_376_6[2], addr_376_6, addr_positional[6027:6024], addr_1506_7);

wire[31:0] addr_1507_7;

Selector_2 s1507_7(wires_376_6[3], addr_376_6, addr_positional[6031:6028], addr_1507_7);

wire[31:0] addr_1508_7;

Selector_2 s1508_7(wires_377_6[0], addr_377_6, addr_positional[6035:6032], addr_1508_7);

wire[31:0] addr_1509_7;

Selector_2 s1509_7(wires_377_6[1], addr_377_6, addr_positional[6039:6036], addr_1509_7);

wire[31:0] addr_1510_7;

Selector_2 s1510_7(wires_377_6[2], addr_377_6, addr_positional[6043:6040], addr_1510_7);

wire[31:0] addr_1511_7;

Selector_2 s1511_7(wires_377_6[3], addr_377_6, addr_positional[6047:6044], addr_1511_7);

wire[31:0] addr_1512_7;

Selector_2 s1512_7(wires_378_6[0], addr_378_6, addr_positional[6051:6048], addr_1512_7);

wire[31:0] addr_1513_7;

Selector_2 s1513_7(wires_378_6[1], addr_378_6, addr_positional[6055:6052], addr_1513_7);

wire[31:0] addr_1514_7;

Selector_2 s1514_7(wires_378_6[2], addr_378_6, addr_positional[6059:6056], addr_1514_7);

wire[31:0] addr_1515_7;

Selector_2 s1515_7(wires_378_6[3], addr_378_6, addr_positional[6063:6060], addr_1515_7);

wire[31:0] addr_1516_7;

Selector_2 s1516_7(wires_379_6[0], addr_379_6, addr_positional[6067:6064], addr_1516_7);

wire[31:0] addr_1517_7;

Selector_2 s1517_7(wires_379_6[1], addr_379_6, addr_positional[6071:6068], addr_1517_7);

wire[31:0] addr_1518_7;

Selector_2 s1518_7(wires_379_6[2], addr_379_6, addr_positional[6075:6072], addr_1518_7);

wire[31:0] addr_1519_7;

Selector_2 s1519_7(wires_379_6[3], addr_379_6, addr_positional[6079:6076], addr_1519_7);

wire[31:0] addr_1520_7;

Selector_2 s1520_7(wires_380_6[0], addr_380_6, addr_positional[6083:6080], addr_1520_7);

wire[31:0] addr_1521_7;

Selector_2 s1521_7(wires_380_6[1], addr_380_6, addr_positional[6087:6084], addr_1521_7);

wire[31:0] addr_1522_7;

Selector_2 s1522_7(wires_380_6[2], addr_380_6, addr_positional[6091:6088], addr_1522_7);

wire[31:0] addr_1523_7;

Selector_2 s1523_7(wires_380_6[3], addr_380_6, addr_positional[6095:6092], addr_1523_7);

wire[31:0] addr_1524_7;

Selector_2 s1524_7(wires_381_6[0], addr_381_6, addr_positional[6099:6096], addr_1524_7);

wire[31:0] addr_1525_7;

Selector_2 s1525_7(wires_381_6[1], addr_381_6, addr_positional[6103:6100], addr_1525_7);

wire[31:0] addr_1526_7;

Selector_2 s1526_7(wires_381_6[2], addr_381_6, addr_positional[6107:6104], addr_1526_7);

wire[31:0] addr_1527_7;

Selector_2 s1527_7(wires_381_6[3], addr_381_6, addr_positional[6111:6108], addr_1527_7);

wire[31:0] addr_1528_7;

Selector_2 s1528_7(wires_382_6[0], addr_382_6, addr_positional[6115:6112], addr_1528_7);

wire[31:0] addr_1529_7;

Selector_2 s1529_7(wires_382_6[1], addr_382_6, addr_positional[6119:6116], addr_1529_7);

wire[31:0] addr_1530_7;

Selector_2 s1530_7(wires_382_6[2], addr_382_6, addr_positional[6123:6120], addr_1530_7);

wire[31:0] addr_1531_7;

Selector_2 s1531_7(wires_382_6[3], addr_382_6, addr_positional[6127:6124], addr_1531_7);

wire[31:0] addr_1532_7;

Selector_2 s1532_7(wires_383_6[0], addr_383_6, addr_positional[6131:6128], addr_1532_7);

wire[31:0] addr_1533_7;

Selector_2 s1533_7(wires_383_6[1], addr_383_6, addr_positional[6135:6132], addr_1533_7);

wire[31:0] addr_1534_7;

Selector_2 s1534_7(wires_383_6[2], addr_383_6, addr_positional[6139:6136], addr_1534_7);

wire[31:0] addr_1535_7;

Selector_2 s1535_7(wires_383_6[3], addr_383_6, addr_positional[6143:6140], addr_1535_7);

wire[31:0] addr_1536_7;

Selector_2 s1536_7(wires_384_6[0], addr_384_6, addr_positional[6147:6144], addr_1536_7);

wire[31:0] addr_1537_7;

Selector_2 s1537_7(wires_384_6[1], addr_384_6, addr_positional[6151:6148], addr_1537_7);

wire[31:0] addr_1538_7;

Selector_2 s1538_7(wires_384_6[2], addr_384_6, addr_positional[6155:6152], addr_1538_7);

wire[31:0] addr_1539_7;

Selector_2 s1539_7(wires_384_6[3], addr_384_6, addr_positional[6159:6156], addr_1539_7);

wire[31:0] addr_1540_7;

Selector_2 s1540_7(wires_385_6[0], addr_385_6, addr_positional[6163:6160], addr_1540_7);

wire[31:0] addr_1541_7;

Selector_2 s1541_7(wires_385_6[1], addr_385_6, addr_positional[6167:6164], addr_1541_7);

wire[31:0] addr_1542_7;

Selector_2 s1542_7(wires_385_6[2], addr_385_6, addr_positional[6171:6168], addr_1542_7);

wire[31:0] addr_1543_7;

Selector_2 s1543_7(wires_385_6[3], addr_385_6, addr_positional[6175:6172], addr_1543_7);

wire[31:0] addr_1544_7;

Selector_2 s1544_7(wires_386_6[0], addr_386_6, addr_positional[6179:6176], addr_1544_7);

wire[31:0] addr_1545_7;

Selector_2 s1545_7(wires_386_6[1], addr_386_6, addr_positional[6183:6180], addr_1545_7);

wire[31:0] addr_1546_7;

Selector_2 s1546_7(wires_386_6[2], addr_386_6, addr_positional[6187:6184], addr_1546_7);

wire[31:0] addr_1547_7;

Selector_2 s1547_7(wires_386_6[3], addr_386_6, addr_positional[6191:6188], addr_1547_7);

wire[31:0] addr_1548_7;

Selector_2 s1548_7(wires_387_6[0], addr_387_6, addr_positional[6195:6192], addr_1548_7);

wire[31:0] addr_1549_7;

Selector_2 s1549_7(wires_387_6[1], addr_387_6, addr_positional[6199:6196], addr_1549_7);

wire[31:0] addr_1550_7;

Selector_2 s1550_7(wires_387_6[2], addr_387_6, addr_positional[6203:6200], addr_1550_7);

wire[31:0] addr_1551_7;

Selector_2 s1551_7(wires_387_6[3], addr_387_6, addr_positional[6207:6204], addr_1551_7);

wire[31:0] addr_1552_7;

Selector_2 s1552_7(wires_388_6[0], addr_388_6, addr_positional[6211:6208], addr_1552_7);

wire[31:0] addr_1553_7;

Selector_2 s1553_7(wires_388_6[1], addr_388_6, addr_positional[6215:6212], addr_1553_7);

wire[31:0] addr_1554_7;

Selector_2 s1554_7(wires_388_6[2], addr_388_6, addr_positional[6219:6216], addr_1554_7);

wire[31:0] addr_1555_7;

Selector_2 s1555_7(wires_388_6[3], addr_388_6, addr_positional[6223:6220], addr_1555_7);

wire[31:0] addr_1556_7;

Selector_2 s1556_7(wires_389_6[0], addr_389_6, addr_positional[6227:6224], addr_1556_7);

wire[31:0] addr_1557_7;

Selector_2 s1557_7(wires_389_6[1], addr_389_6, addr_positional[6231:6228], addr_1557_7);

wire[31:0] addr_1558_7;

Selector_2 s1558_7(wires_389_6[2], addr_389_6, addr_positional[6235:6232], addr_1558_7);

wire[31:0] addr_1559_7;

Selector_2 s1559_7(wires_389_6[3], addr_389_6, addr_positional[6239:6236], addr_1559_7);

wire[31:0] addr_1560_7;

Selector_2 s1560_7(wires_390_6[0], addr_390_6, addr_positional[6243:6240], addr_1560_7);

wire[31:0] addr_1561_7;

Selector_2 s1561_7(wires_390_6[1], addr_390_6, addr_positional[6247:6244], addr_1561_7);

wire[31:0] addr_1562_7;

Selector_2 s1562_7(wires_390_6[2], addr_390_6, addr_positional[6251:6248], addr_1562_7);

wire[31:0] addr_1563_7;

Selector_2 s1563_7(wires_390_6[3], addr_390_6, addr_positional[6255:6252], addr_1563_7);

wire[31:0] addr_1564_7;

Selector_2 s1564_7(wires_391_6[0], addr_391_6, addr_positional[6259:6256], addr_1564_7);

wire[31:0] addr_1565_7;

Selector_2 s1565_7(wires_391_6[1], addr_391_6, addr_positional[6263:6260], addr_1565_7);

wire[31:0] addr_1566_7;

Selector_2 s1566_7(wires_391_6[2], addr_391_6, addr_positional[6267:6264], addr_1566_7);

wire[31:0] addr_1567_7;

Selector_2 s1567_7(wires_391_6[3], addr_391_6, addr_positional[6271:6268], addr_1567_7);

wire[31:0] addr_1568_7;

Selector_2 s1568_7(wires_392_6[0], addr_392_6, addr_positional[6275:6272], addr_1568_7);

wire[31:0] addr_1569_7;

Selector_2 s1569_7(wires_392_6[1], addr_392_6, addr_positional[6279:6276], addr_1569_7);

wire[31:0] addr_1570_7;

Selector_2 s1570_7(wires_392_6[2], addr_392_6, addr_positional[6283:6280], addr_1570_7);

wire[31:0] addr_1571_7;

Selector_2 s1571_7(wires_392_6[3], addr_392_6, addr_positional[6287:6284], addr_1571_7);

wire[31:0] addr_1572_7;

Selector_2 s1572_7(wires_393_6[0], addr_393_6, addr_positional[6291:6288], addr_1572_7);

wire[31:0] addr_1573_7;

Selector_2 s1573_7(wires_393_6[1], addr_393_6, addr_positional[6295:6292], addr_1573_7);

wire[31:0] addr_1574_7;

Selector_2 s1574_7(wires_393_6[2], addr_393_6, addr_positional[6299:6296], addr_1574_7);

wire[31:0] addr_1575_7;

Selector_2 s1575_7(wires_393_6[3], addr_393_6, addr_positional[6303:6300], addr_1575_7);

wire[31:0] addr_1576_7;

Selector_2 s1576_7(wires_394_6[0], addr_394_6, addr_positional[6307:6304], addr_1576_7);

wire[31:0] addr_1577_7;

Selector_2 s1577_7(wires_394_6[1], addr_394_6, addr_positional[6311:6308], addr_1577_7);

wire[31:0] addr_1578_7;

Selector_2 s1578_7(wires_394_6[2], addr_394_6, addr_positional[6315:6312], addr_1578_7);

wire[31:0] addr_1579_7;

Selector_2 s1579_7(wires_394_6[3], addr_394_6, addr_positional[6319:6316], addr_1579_7);

wire[31:0] addr_1580_7;

Selector_2 s1580_7(wires_395_6[0], addr_395_6, addr_positional[6323:6320], addr_1580_7);

wire[31:0] addr_1581_7;

Selector_2 s1581_7(wires_395_6[1], addr_395_6, addr_positional[6327:6324], addr_1581_7);

wire[31:0] addr_1582_7;

Selector_2 s1582_7(wires_395_6[2], addr_395_6, addr_positional[6331:6328], addr_1582_7);

wire[31:0] addr_1583_7;

Selector_2 s1583_7(wires_395_6[3], addr_395_6, addr_positional[6335:6332], addr_1583_7);

wire[31:0] addr_1584_7;

Selector_2 s1584_7(wires_396_6[0], addr_396_6, addr_positional[6339:6336], addr_1584_7);

wire[31:0] addr_1585_7;

Selector_2 s1585_7(wires_396_6[1], addr_396_6, addr_positional[6343:6340], addr_1585_7);

wire[31:0] addr_1586_7;

Selector_2 s1586_7(wires_396_6[2], addr_396_6, addr_positional[6347:6344], addr_1586_7);

wire[31:0] addr_1587_7;

Selector_2 s1587_7(wires_396_6[3], addr_396_6, addr_positional[6351:6348], addr_1587_7);

wire[31:0] addr_1588_7;

Selector_2 s1588_7(wires_397_6[0], addr_397_6, addr_positional[6355:6352], addr_1588_7);

wire[31:0] addr_1589_7;

Selector_2 s1589_7(wires_397_6[1], addr_397_6, addr_positional[6359:6356], addr_1589_7);

wire[31:0] addr_1590_7;

Selector_2 s1590_7(wires_397_6[2], addr_397_6, addr_positional[6363:6360], addr_1590_7);

wire[31:0] addr_1591_7;

Selector_2 s1591_7(wires_397_6[3], addr_397_6, addr_positional[6367:6364], addr_1591_7);

wire[31:0] addr_1592_7;

Selector_2 s1592_7(wires_398_6[0], addr_398_6, addr_positional[6371:6368], addr_1592_7);

wire[31:0] addr_1593_7;

Selector_2 s1593_7(wires_398_6[1], addr_398_6, addr_positional[6375:6372], addr_1593_7);

wire[31:0] addr_1594_7;

Selector_2 s1594_7(wires_398_6[2], addr_398_6, addr_positional[6379:6376], addr_1594_7);

wire[31:0] addr_1595_7;

Selector_2 s1595_7(wires_398_6[3], addr_398_6, addr_positional[6383:6380], addr_1595_7);

wire[31:0] addr_1596_7;

Selector_2 s1596_7(wires_399_6[0], addr_399_6, addr_positional[6387:6384], addr_1596_7);

wire[31:0] addr_1597_7;

Selector_2 s1597_7(wires_399_6[1], addr_399_6, addr_positional[6391:6388], addr_1597_7);

wire[31:0] addr_1598_7;

Selector_2 s1598_7(wires_399_6[2], addr_399_6, addr_positional[6395:6392], addr_1598_7);

wire[31:0] addr_1599_7;

Selector_2 s1599_7(wires_399_6[3], addr_399_6, addr_positional[6399:6396], addr_1599_7);

wire[31:0] addr_1600_7;

Selector_2 s1600_7(wires_400_6[0], addr_400_6, addr_positional[6403:6400], addr_1600_7);

wire[31:0] addr_1601_7;

Selector_2 s1601_7(wires_400_6[1], addr_400_6, addr_positional[6407:6404], addr_1601_7);

wire[31:0] addr_1602_7;

Selector_2 s1602_7(wires_400_6[2], addr_400_6, addr_positional[6411:6408], addr_1602_7);

wire[31:0] addr_1603_7;

Selector_2 s1603_7(wires_400_6[3], addr_400_6, addr_positional[6415:6412], addr_1603_7);

wire[31:0] addr_1604_7;

Selector_2 s1604_7(wires_401_6[0], addr_401_6, addr_positional[6419:6416], addr_1604_7);

wire[31:0] addr_1605_7;

Selector_2 s1605_7(wires_401_6[1], addr_401_6, addr_positional[6423:6420], addr_1605_7);

wire[31:0] addr_1606_7;

Selector_2 s1606_7(wires_401_6[2], addr_401_6, addr_positional[6427:6424], addr_1606_7);

wire[31:0] addr_1607_7;

Selector_2 s1607_7(wires_401_6[3], addr_401_6, addr_positional[6431:6428], addr_1607_7);

wire[31:0] addr_1608_7;

Selector_2 s1608_7(wires_402_6[0], addr_402_6, addr_positional[6435:6432], addr_1608_7);

wire[31:0] addr_1609_7;

Selector_2 s1609_7(wires_402_6[1], addr_402_6, addr_positional[6439:6436], addr_1609_7);

wire[31:0] addr_1610_7;

Selector_2 s1610_7(wires_402_6[2], addr_402_6, addr_positional[6443:6440], addr_1610_7);

wire[31:0] addr_1611_7;

Selector_2 s1611_7(wires_402_6[3], addr_402_6, addr_positional[6447:6444], addr_1611_7);

wire[31:0] addr_1612_7;

Selector_2 s1612_7(wires_403_6[0], addr_403_6, addr_positional[6451:6448], addr_1612_7);

wire[31:0] addr_1613_7;

Selector_2 s1613_7(wires_403_6[1], addr_403_6, addr_positional[6455:6452], addr_1613_7);

wire[31:0] addr_1614_7;

Selector_2 s1614_7(wires_403_6[2], addr_403_6, addr_positional[6459:6456], addr_1614_7);

wire[31:0] addr_1615_7;

Selector_2 s1615_7(wires_403_6[3], addr_403_6, addr_positional[6463:6460], addr_1615_7);

wire[31:0] addr_1616_7;

Selector_2 s1616_7(wires_404_6[0], addr_404_6, addr_positional[6467:6464], addr_1616_7);

wire[31:0] addr_1617_7;

Selector_2 s1617_7(wires_404_6[1], addr_404_6, addr_positional[6471:6468], addr_1617_7);

wire[31:0] addr_1618_7;

Selector_2 s1618_7(wires_404_6[2], addr_404_6, addr_positional[6475:6472], addr_1618_7);

wire[31:0] addr_1619_7;

Selector_2 s1619_7(wires_404_6[3], addr_404_6, addr_positional[6479:6476], addr_1619_7);

wire[31:0] addr_1620_7;

Selector_2 s1620_7(wires_405_6[0], addr_405_6, addr_positional[6483:6480], addr_1620_7);

wire[31:0] addr_1621_7;

Selector_2 s1621_7(wires_405_6[1], addr_405_6, addr_positional[6487:6484], addr_1621_7);

wire[31:0] addr_1622_7;

Selector_2 s1622_7(wires_405_6[2], addr_405_6, addr_positional[6491:6488], addr_1622_7);

wire[31:0] addr_1623_7;

Selector_2 s1623_7(wires_405_6[3], addr_405_6, addr_positional[6495:6492], addr_1623_7);

wire[31:0] addr_1624_7;

Selector_2 s1624_7(wires_406_6[0], addr_406_6, addr_positional[6499:6496], addr_1624_7);

wire[31:0] addr_1625_7;

Selector_2 s1625_7(wires_406_6[1], addr_406_6, addr_positional[6503:6500], addr_1625_7);

wire[31:0] addr_1626_7;

Selector_2 s1626_7(wires_406_6[2], addr_406_6, addr_positional[6507:6504], addr_1626_7);

wire[31:0] addr_1627_7;

Selector_2 s1627_7(wires_406_6[3], addr_406_6, addr_positional[6511:6508], addr_1627_7);

wire[31:0] addr_1628_7;

Selector_2 s1628_7(wires_407_6[0], addr_407_6, addr_positional[6515:6512], addr_1628_7);

wire[31:0] addr_1629_7;

Selector_2 s1629_7(wires_407_6[1], addr_407_6, addr_positional[6519:6516], addr_1629_7);

wire[31:0] addr_1630_7;

Selector_2 s1630_7(wires_407_6[2], addr_407_6, addr_positional[6523:6520], addr_1630_7);

wire[31:0] addr_1631_7;

Selector_2 s1631_7(wires_407_6[3], addr_407_6, addr_positional[6527:6524], addr_1631_7);

wire[31:0] addr_1632_7;

Selector_2 s1632_7(wires_408_6[0], addr_408_6, addr_positional[6531:6528], addr_1632_7);

wire[31:0] addr_1633_7;

Selector_2 s1633_7(wires_408_6[1], addr_408_6, addr_positional[6535:6532], addr_1633_7);

wire[31:0] addr_1634_7;

Selector_2 s1634_7(wires_408_6[2], addr_408_6, addr_positional[6539:6536], addr_1634_7);

wire[31:0] addr_1635_7;

Selector_2 s1635_7(wires_408_6[3], addr_408_6, addr_positional[6543:6540], addr_1635_7);

wire[31:0] addr_1636_7;

Selector_2 s1636_7(wires_409_6[0], addr_409_6, addr_positional[6547:6544], addr_1636_7);

wire[31:0] addr_1637_7;

Selector_2 s1637_7(wires_409_6[1], addr_409_6, addr_positional[6551:6548], addr_1637_7);

wire[31:0] addr_1638_7;

Selector_2 s1638_7(wires_409_6[2], addr_409_6, addr_positional[6555:6552], addr_1638_7);

wire[31:0] addr_1639_7;

Selector_2 s1639_7(wires_409_6[3], addr_409_6, addr_positional[6559:6556], addr_1639_7);

wire[31:0] addr_1640_7;

Selector_2 s1640_7(wires_410_6[0], addr_410_6, addr_positional[6563:6560], addr_1640_7);

wire[31:0] addr_1641_7;

Selector_2 s1641_7(wires_410_6[1], addr_410_6, addr_positional[6567:6564], addr_1641_7);

wire[31:0] addr_1642_7;

Selector_2 s1642_7(wires_410_6[2], addr_410_6, addr_positional[6571:6568], addr_1642_7);

wire[31:0] addr_1643_7;

Selector_2 s1643_7(wires_410_6[3], addr_410_6, addr_positional[6575:6572], addr_1643_7);

wire[31:0] addr_1644_7;

Selector_2 s1644_7(wires_411_6[0], addr_411_6, addr_positional[6579:6576], addr_1644_7);

wire[31:0] addr_1645_7;

Selector_2 s1645_7(wires_411_6[1], addr_411_6, addr_positional[6583:6580], addr_1645_7);

wire[31:0] addr_1646_7;

Selector_2 s1646_7(wires_411_6[2], addr_411_6, addr_positional[6587:6584], addr_1646_7);

wire[31:0] addr_1647_7;

Selector_2 s1647_7(wires_411_6[3], addr_411_6, addr_positional[6591:6588], addr_1647_7);

wire[31:0] addr_1648_7;

Selector_2 s1648_7(wires_412_6[0], addr_412_6, addr_positional[6595:6592], addr_1648_7);

wire[31:0] addr_1649_7;

Selector_2 s1649_7(wires_412_6[1], addr_412_6, addr_positional[6599:6596], addr_1649_7);

wire[31:0] addr_1650_7;

Selector_2 s1650_7(wires_412_6[2], addr_412_6, addr_positional[6603:6600], addr_1650_7);

wire[31:0] addr_1651_7;

Selector_2 s1651_7(wires_412_6[3], addr_412_6, addr_positional[6607:6604], addr_1651_7);

wire[31:0] addr_1652_7;

Selector_2 s1652_7(wires_413_6[0], addr_413_6, addr_positional[6611:6608], addr_1652_7);

wire[31:0] addr_1653_7;

Selector_2 s1653_7(wires_413_6[1], addr_413_6, addr_positional[6615:6612], addr_1653_7);

wire[31:0] addr_1654_7;

Selector_2 s1654_7(wires_413_6[2], addr_413_6, addr_positional[6619:6616], addr_1654_7);

wire[31:0] addr_1655_7;

Selector_2 s1655_7(wires_413_6[3], addr_413_6, addr_positional[6623:6620], addr_1655_7);

wire[31:0] addr_1656_7;

Selector_2 s1656_7(wires_414_6[0], addr_414_6, addr_positional[6627:6624], addr_1656_7);

wire[31:0] addr_1657_7;

Selector_2 s1657_7(wires_414_6[1], addr_414_6, addr_positional[6631:6628], addr_1657_7);

wire[31:0] addr_1658_7;

Selector_2 s1658_7(wires_414_6[2], addr_414_6, addr_positional[6635:6632], addr_1658_7);

wire[31:0] addr_1659_7;

Selector_2 s1659_7(wires_414_6[3], addr_414_6, addr_positional[6639:6636], addr_1659_7);

wire[31:0] addr_1660_7;

Selector_2 s1660_7(wires_415_6[0], addr_415_6, addr_positional[6643:6640], addr_1660_7);

wire[31:0] addr_1661_7;

Selector_2 s1661_7(wires_415_6[1], addr_415_6, addr_positional[6647:6644], addr_1661_7);

wire[31:0] addr_1662_7;

Selector_2 s1662_7(wires_415_6[2], addr_415_6, addr_positional[6651:6648], addr_1662_7);

wire[31:0] addr_1663_7;

Selector_2 s1663_7(wires_415_6[3], addr_415_6, addr_positional[6655:6652], addr_1663_7);

wire[31:0] addr_1664_7;

Selector_2 s1664_7(wires_416_6[0], addr_416_6, addr_positional[6659:6656], addr_1664_7);

wire[31:0] addr_1665_7;

Selector_2 s1665_7(wires_416_6[1], addr_416_6, addr_positional[6663:6660], addr_1665_7);

wire[31:0] addr_1666_7;

Selector_2 s1666_7(wires_416_6[2], addr_416_6, addr_positional[6667:6664], addr_1666_7);

wire[31:0] addr_1667_7;

Selector_2 s1667_7(wires_416_6[3], addr_416_6, addr_positional[6671:6668], addr_1667_7);

wire[31:0] addr_1668_7;

Selector_2 s1668_7(wires_417_6[0], addr_417_6, addr_positional[6675:6672], addr_1668_7);

wire[31:0] addr_1669_7;

Selector_2 s1669_7(wires_417_6[1], addr_417_6, addr_positional[6679:6676], addr_1669_7);

wire[31:0] addr_1670_7;

Selector_2 s1670_7(wires_417_6[2], addr_417_6, addr_positional[6683:6680], addr_1670_7);

wire[31:0] addr_1671_7;

Selector_2 s1671_7(wires_417_6[3], addr_417_6, addr_positional[6687:6684], addr_1671_7);

wire[31:0] addr_1672_7;

Selector_2 s1672_7(wires_418_6[0], addr_418_6, addr_positional[6691:6688], addr_1672_7);

wire[31:0] addr_1673_7;

Selector_2 s1673_7(wires_418_6[1], addr_418_6, addr_positional[6695:6692], addr_1673_7);

wire[31:0] addr_1674_7;

Selector_2 s1674_7(wires_418_6[2], addr_418_6, addr_positional[6699:6696], addr_1674_7);

wire[31:0] addr_1675_7;

Selector_2 s1675_7(wires_418_6[3], addr_418_6, addr_positional[6703:6700], addr_1675_7);

wire[31:0] addr_1676_7;

Selector_2 s1676_7(wires_419_6[0], addr_419_6, addr_positional[6707:6704], addr_1676_7);

wire[31:0] addr_1677_7;

Selector_2 s1677_7(wires_419_6[1], addr_419_6, addr_positional[6711:6708], addr_1677_7);

wire[31:0] addr_1678_7;

Selector_2 s1678_7(wires_419_6[2], addr_419_6, addr_positional[6715:6712], addr_1678_7);

wire[31:0] addr_1679_7;

Selector_2 s1679_7(wires_419_6[3], addr_419_6, addr_positional[6719:6716], addr_1679_7);

wire[31:0] addr_1680_7;

Selector_2 s1680_7(wires_420_6[0], addr_420_6, addr_positional[6723:6720], addr_1680_7);

wire[31:0] addr_1681_7;

Selector_2 s1681_7(wires_420_6[1], addr_420_6, addr_positional[6727:6724], addr_1681_7);

wire[31:0] addr_1682_7;

Selector_2 s1682_7(wires_420_6[2], addr_420_6, addr_positional[6731:6728], addr_1682_7);

wire[31:0] addr_1683_7;

Selector_2 s1683_7(wires_420_6[3], addr_420_6, addr_positional[6735:6732], addr_1683_7);

wire[31:0] addr_1684_7;

Selector_2 s1684_7(wires_421_6[0], addr_421_6, addr_positional[6739:6736], addr_1684_7);

wire[31:0] addr_1685_7;

Selector_2 s1685_7(wires_421_6[1], addr_421_6, addr_positional[6743:6740], addr_1685_7);

wire[31:0] addr_1686_7;

Selector_2 s1686_7(wires_421_6[2], addr_421_6, addr_positional[6747:6744], addr_1686_7);

wire[31:0] addr_1687_7;

Selector_2 s1687_7(wires_421_6[3], addr_421_6, addr_positional[6751:6748], addr_1687_7);

wire[31:0] addr_1688_7;

Selector_2 s1688_7(wires_422_6[0], addr_422_6, addr_positional[6755:6752], addr_1688_7);

wire[31:0] addr_1689_7;

Selector_2 s1689_7(wires_422_6[1], addr_422_6, addr_positional[6759:6756], addr_1689_7);

wire[31:0] addr_1690_7;

Selector_2 s1690_7(wires_422_6[2], addr_422_6, addr_positional[6763:6760], addr_1690_7);

wire[31:0] addr_1691_7;

Selector_2 s1691_7(wires_422_6[3], addr_422_6, addr_positional[6767:6764], addr_1691_7);

wire[31:0] addr_1692_7;

Selector_2 s1692_7(wires_423_6[0], addr_423_6, addr_positional[6771:6768], addr_1692_7);

wire[31:0] addr_1693_7;

Selector_2 s1693_7(wires_423_6[1], addr_423_6, addr_positional[6775:6772], addr_1693_7);

wire[31:0] addr_1694_7;

Selector_2 s1694_7(wires_423_6[2], addr_423_6, addr_positional[6779:6776], addr_1694_7);

wire[31:0] addr_1695_7;

Selector_2 s1695_7(wires_423_6[3], addr_423_6, addr_positional[6783:6780], addr_1695_7);

wire[31:0] addr_1696_7;

Selector_2 s1696_7(wires_424_6[0], addr_424_6, addr_positional[6787:6784], addr_1696_7);

wire[31:0] addr_1697_7;

Selector_2 s1697_7(wires_424_6[1], addr_424_6, addr_positional[6791:6788], addr_1697_7);

wire[31:0] addr_1698_7;

Selector_2 s1698_7(wires_424_6[2], addr_424_6, addr_positional[6795:6792], addr_1698_7);

wire[31:0] addr_1699_7;

Selector_2 s1699_7(wires_424_6[3], addr_424_6, addr_positional[6799:6796], addr_1699_7);

wire[31:0] addr_1700_7;

Selector_2 s1700_7(wires_425_6[0], addr_425_6, addr_positional[6803:6800], addr_1700_7);

wire[31:0] addr_1701_7;

Selector_2 s1701_7(wires_425_6[1], addr_425_6, addr_positional[6807:6804], addr_1701_7);

wire[31:0] addr_1702_7;

Selector_2 s1702_7(wires_425_6[2], addr_425_6, addr_positional[6811:6808], addr_1702_7);

wire[31:0] addr_1703_7;

Selector_2 s1703_7(wires_425_6[3], addr_425_6, addr_positional[6815:6812], addr_1703_7);

wire[31:0] addr_1704_7;

Selector_2 s1704_7(wires_426_6[0], addr_426_6, addr_positional[6819:6816], addr_1704_7);

wire[31:0] addr_1705_7;

Selector_2 s1705_7(wires_426_6[1], addr_426_6, addr_positional[6823:6820], addr_1705_7);

wire[31:0] addr_1706_7;

Selector_2 s1706_7(wires_426_6[2], addr_426_6, addr_positional[6827:6824], addr_1706_7);

wire[31:0] addr_1707_7;

Selector_2 s1707_7(wires_426_6[3], addr_426_6, addr_positional[6831:6828], addr_1707_7);

wire[31:0] addr_1708_7;

Selector_2 s1708_7(wires_427_6[0], addr_427_6, addr_positional[6835:6832], addr_1708_7);

wire[31:0] addr_1709_7;

Selector_2 s1709_7(wires_427_6[1], addr_427_6, addr_positional[6839:6836], addr_1709_7);

wire[31:0] addr_1710_7;

Selector_2 s1710_7(wires_427_6[2], addr_427_6, addr_positional[6843:6840], addr_1710_7);

wire[31:0] addr_1711_7;

Selector_2 s1711_7(wires_427_6[3], addr_427_6, addr_positional[6847:6844], addr_1711_7);

wire[31:0] addr_1712_7;

Selector_2 s1712_7(wires_428_6[0], addr_428_6, addr_positional[6851:6848], addr_1712_7);

wire[31:0] addr_1713_7;

Selector_2 s1713_7(wires_428_6[1], addr_428_6, addr_positional[6855:6852], addr_1713_7);

wire[31:0] addr_1714_7;

Selector_2 s1714_7(wires_428_6[2], addr_428_6, addr_positional[6859:6856], addr_1714_7);

wire[31:0] addr_1715_7;

Selector_2 s1715_7(wires_428_6[3], addr_428_6, addr_positional[6863:6860], addr_1715_7);

wire[31:0] addr_1716_7;

Selector_2 s1716_7(wires_429_6[0], addr_429_6, addr_positional[6867:6864], addr_1716_7);

wire[31:0] addr_1717_7;

Selector_2 s1717_7(wires_429_6[1], addr_429_6, addr_positional[6871:6868], addr_1717_7);

wire[31:0] addr_1718_7;

Selector_2 s1718_7(wires_429_6[2], addr_429_6, addr_positional[6875:6872], addr_1718_7);

wire[31:0] addr_1719_7;

Selector_2 s1719_7(wires_429_6[3], addr_429_6, addr_positional[6879:6876], addr_1719_7);

wire[31:0] addr_1720_7;

Selector_2 s1720_7(wires_430_6[0], addr_430_6, addr_positional[6883:6880], addr_1720_7);

wire[31:0] addr_1721_7;

Selector_2 s1721_7(wires_430_6[1], addr_430_6, addr_positional[6887:6884], addr_1721_7);

wire[31:0] addr_1722_7;

Selector_2 s1722_7(wires_430_6[2], addr_430_6, addr_positional[6891:6888], addr_1722_7);

wire[31:0] addr_1723_7;

Selector_2 s1723_7(wires_430_6[3], addr_430_6, addr_positional[6895:6892], addr_1723_7);

wire[31:0] addr_1724_7;

Selector_2 s1724_7(wires_431_6[0], addr_431_6, addr_positional[6899:6896], addr_1724_7);

wire[31:0] addr_1725_7;

Selector_2 s1725_7(wires_431_6[1], addr_431_6, addr_positional[6903:6900], addr_1725_7);

wire[31:0] addr_1726_7;

Selector_2 s1726_7(wires_431_6[2], addr_431_6, addr_positional[6907:6904], addr_1726_7);

wire[31:0] addr_1727_7;

Selector_2 s1727_7(wires_431_6[3], addr_431_6, addr_positional[6911:6908], addr_1727_7);

wire[31:0] addr_1728_7;

Selector_2 s1728_7(wires_432_6[0], addr_432_6, addr_positional[6915:6912], addr_1728_7);

wire[31:0] addr_1729_7;

Selector_2 s1729_7(wires_432_6[1], addr_432_6, addr_positional[6919:6916], addr_1729_7);

wire[31:0] addr_1730_7;

Selector_2 s1730_7(wires_432_6[2], addr_432_6, addr_positional[6923:6920], addr_1730_7);

wire[31:0] addr_1731_7;

Selector_2 s1731_7(wires_432_6[3], addr_432_6, addr_positional[6927:6924], addr_1731_7);

wire[31:0] addr_1732_7;

Selector_2 s1732_7(wires_433_6[0], addr_433_6, addr_positional[6931:6928], addr_1732_7);

wire[31:0] addr_1733_7;

Selector_2 s1733_7(wires_433_6[1], addr_433_6, addr_positional[6935:6932], addr_1733_7);

wire[31:0] addr_1734_7;

Selector_2 s1734_7(wires_433_6[2], addr_433_6, addr_positional[6939:6936], addr_1734_7);

wire[31:0] addr_1735_7;

Selector_2 s1735_7(wires_433_6[3], addr_433_6, addr_positional[6943:6940], addr_1735_7);

wire[31:0] addr_1736_7;

Selector_2 s1736_7(wires_434_6[0], addr_434_6, addr_positional[6947:6944], addr_1736_7);

wire[31:0] addr_1737_7;

Selector_2 s1737_7(wires_434_6[1], addr_434_6, addr_positional[6951:6948], addr_1737_7);

wire[31:0] addr_1738_7;

Selector_2 s1738_7(wires_434_6[2], addr_434_6, addr_positional[6955:6952], addr_1738_7);

wire[31:0] addr_1739_7;

Selector_2 s1739_7(wires_434_6[3], addr_434_6, addr_positional[6959:6956], addr_1739_7);

wire[31:0] addr_1740_7;

Selector_2 s1740_7(wires_435_6[0], addr_435_6, addr_positional[6963:6960], addr_1740_7);

wire[31:0] addr_1741_7;

Selector_2 s1741_7(wires_435_6[1], addr_435_6, addr_positional[6967:6964], addr_1741_7);

wire[31:0] addr_1742_7;

Selector_2 s1742_7(wires_435_6[2], addr_435_6, addr_positional[6971:6968], addr_1742_7);

wire[31:0] addr_1743_7;

Selector_2 s1743_7(wires_435_6[3], addr_435_6, addr_positional[6975:6972], addr_1743_7);

wire[31:0] addr_1744_7;

Selector_2 s1744_7(wires_436_6[0], addr_436_6, addr_positional[6979:6976], addr_1744_7);

wire[31:0] addr_1745_7;

Selector_2 s1745_7(wires_436_6[1], addr_436_6, addr_positional[6983:6980], addr_1745_7);

wire[31:0] addr_1746_7;

Selector_2 s1746_7(wires_436_6[2], addr_436_6, addr_positional[6987:6984], addr_1746_7);

wire[31:0] addr_1747_7;

Selector_2 s1747_7(wires_436_6[3], addr_436_6, addr_positional[6991:6988], addr_1747_7);

wire[31:0] addr_1748_7;

Selector_2 s1748_7(wires_437_6[0], addr_437_6, addr_positional[6995:6992], addr_1748_7);

wire[31:0] addr_1749_7;

Selector_2 s1749_7(wires_437_6[1], addr_437_6, addr_positional[6999:6996], addr_1749_7);

wire[31:0] addr_1750_7;

Selector_2 s1750_7(wires_437_6[2], addr_437_6, addr_positional[7003:7000], addr_1750_7);

wire[31:0] addr_1751_7;

Selector_2 s1751_7(wires_437_6[3], addr_437_6, addr_positional[7007:7004], addr_1751_7);

wire[31:0] addr_1752_7;

Selector_2 s1752_7(wires_438_6[0], addr_438_6, addr_positional[7011:7008], addr_1752_7);

wire[31:0] addr_1753_7;

Selector_2 s1753_7(wires_438_6[1], addr_438_6, addr_positional[7015:7012], addr_1753_7);

wire[31:0] addr_1754_7;

Selector_2 s1754_7(wires_438_6[2], addr_438_6, addr_positional[7019:7016], addr_1754_7);

wire[31:0] addr_1755_7;

Selector_2 s1755_7(wires_438_6[3], addr_438_6, addr_positional[7023:7020], addr_1755_7);

wire[31:0] addr_1756_7;

Selector_2 s1756_7(wires_439_6[0], addr_439_6, addr_positional[7027:7024], addr_1756_7);

wire[31:0] addr_1757_7;

Selector_2 s1757_7(wires_439_6[1], addr_439_6, addr_positional[7031:7028], addr_1757_7);

wire[31:0] addr_1758_7;

Selector_2 s1758_7(wires_439_6[2], addr_439_6, addr_positional[7035:7032], addr_1758_7);

wire[31:0] addr_1759_7;

Selector_2 s1759_7(wires_439_6[3], addr_439_6, addr_positional[7039:7036], addr_1759_7);

wire[31:0] addr_1760_7;

Selector_2 s1760_7(wires_440_6[0], addr_440_6, addr_positional[7043:7040], addr_1760_7);

wire[31:0] addr_1761_7;

Selector_2 s1761_7(wires_440_6[1], addr_440_6, addr_positional[7047:7044], addr_1761_7);

wire[31:0] addr_1762_7;

Selector_2 s1762_7(wires_440_6[2], addr_440_6, addr_positional[7051:7048], addr_1762_7);

wire[31:0] addr_1763_7;

Selector_2 s1763_7(wires_440_6[3], addr_440_6, addr_positional[7055:7052], addr_1763_7);

wire[31:0] addr_1764_7;

Selector_2 s1764_7(wires_441_6[0], addr_441_6, addr_positional[7059:7056], addr_1764_7);

wire[31:0] addr_1765_7;

Selector_2 s1765_7(wires_441_6[1], addr_441_6, addr_positional[7063:7060], addr_1765_7);

wire[31:0] addr_1766_7;

Selector_2 s1766_7(wires_441_6[2], addr_441_6, addr_positional[7067:7064], addr_1766_7);

wire[31:0] addr_1767_7;

Selector_2 s1767_7(wires_441_6[3], addr_441_6, addr_positional[7071:7068], addr_1767_7);

wire[31:0] addr_1768_7;

Selector_2 s1768_7(wires_442_6[0], addr_442_6, addr_positional[7075:7072], addr_1768_7);

wire[31:0] addr_1769_7;

Selector_2 s1769_7(wires_442_6[1], addr_442_6, addr_positional[7079:7076], addr_1769_7);

wire[31:0] addr_1770_7;

Selector_2 s1770_7(wires_442_6[2], addr_442_6, addr_positional[7083:7080], addr_1770_7);

wire[31:0] addr_1771_7;

Selector_2 s1771_7(wires_442_6[3], addr_442_6, addr_positional[7087:7084], addr_1771_7);

wire[31:0] addr_1772_7;

Selector_2 s1772_7(wires_443_6[0], addr_443_6, addr_positional[7091:7088], addr_1772_7);

wire[31:0] addr_1773_7;

Selector_2 s1773_7(wires_443_6[1], addr_443_6, addr_positional[7095:7092], addr_1773_7);

wire[31:0] addr_1774_7;

Selector_2 s1774_7(wires_443_6[2], addr_443_6, addr_positional[7099:7096], addr_1774_7);

wire[31:0] addr_1775_7;

Selector_2 s1775_7(wires_443_6[3], addr_443_6, addr_positional[7103:7100], addr_1775_7);

wire[31:0] addr_1776_7;

Selector_2 s1776_7(wires_444_6[0], addr_444_6, addr_positional[7107:7104], addr_1776_7);

wire[31:0] addr_1777_7;

Selector_2 s1777_7(wires_444_6[1], addr_444_6, addr_positional[7111:7108], addr_1777_7);

wire[31:0] addr_1778_7;

Selector_2 s1778_7(wires_444_6[2], addr_444_6, addr_positional[7115:7112], addr_1778_7);

wire[31:0] addr_1779_7;

Selector_2 s1779_7(wires_444_6[3], addr_444_6, addr_positional[7119:7116], addr_1779_7);

wire[31:0] addr_1780_7;

Selector_2 s1780_7(wires_445_6[0], addr_445_6, addr_positional[7123:7120], addr_1780_7);

wire[31:0] addr_1781_7;

Selector_2 s1781_7(wires_445_6[1], addr_445_6, addr_positional[7127:7124], addr_1781_7);

wire[31:0] addr_1782_7;

Selector_2 s1782_7(wires_445_6[2], addr_445_6, addr_positional[7131:7128], addr_1782_7);

wire[31:0] addr_1783_7;

Selector_2 s1783_7(wires_445_6[3], addr_445_6, addr_positional[7135:7132], addr_1783_7);

wire[31:0] addr_1784_7;

Selector_2 s1784_7(wires_446_6[0], addr_446_6, addr_positional[7139:7136], addr_1784_7);

wire[31:0] addr_1785_7;

Selector_2 s1785_7(wires_446_6[1], addr_446_6, addr_positional[7143:7140], addr_1785_7);

wire[31:0] addr_1786_7;

Selector_2 s1786_7(wires_446_6[2], addr_446_6, addr_positional[7147:7144], addr_1786_7);

wire[31:0] addr_1787_7;

Selector_2 s1787_7(wires_446_6[3], addr_446_6, addr_positional[7151:7148], addr_1787_7);

wire[31:0] addr_1788_7;

Selector_2 s1788_7(wires_447_6[0], addr_447_6, addr_positional[7155:7152], addr_1788_7);

wire[31:0] addr_1789_7;

Selector_2 s1789_7(wires_447_6[1], addr_447_6, addr_positional[7159:7156], addr_1789_7);

wire[31:0] addr_1790_7;

Selector_2 s1790_7(wires_447_6[2], addr_447_6, addr_positional[7163:7160], addr_1790_7);

wire[31:0] addr_1791_7;

Selector_2 s1791_7(wires_447_6[3], addr_447_6, addr_positional[7167:7164], addr_1791_7);

wire[31:0] addr_1792_7;

Selector_2 s1792_7(wires_448_6[0], addr_448_6, addr_positional[7171:7168], addr_1792_7);

wire[31:0] addr_1793_7;

Selector_2 s1793_7(wires_448_6[1], addr_448_6, addr_positional[7175:7172], addr_1793_7);

wire[31:0] addr_1794_7;

Selector_2 s1794_7(wires_448_6[2], addr_448_6, addr_positional[7179:7176], addr_1794_7);

wire[31:0] addr_1795_7;

Selector_2 s1795_7(wires_448_6[3], addr_448_6, addr_positional[7183:7180], addr_1795_7);

wire[31:0] addr_1796_7;

Selector_2 s1796_7(wires_449_6[0], addr_449_6, addr_positional[7187:7184], addr_1796_7);

wire[31:0] addr_1797_7;

Selector_2 s1797_7(wires_449_6[1], addr_449_6, addr_positional[7191:7188], addr_1797_7);

wire[31:0] addr_1798_7;

Selector_2 s1798_7(wires_449_6[2], addr_449_6, addr_positional[7195:7192], addr_1798_7);

wire[31:0] addr_1799_7;

Selector_2 s1799_7(wires_449_6[3], addr_449_6, addr_positional[7199:7196], addr_1799_7);

wire[31:0] addr_1800_7;

Selector_2 s1800_7(wires_450_6[0], addr_450_6, addr_positional[7203:7200], addr_1800_7);

wire[31:0] addr_1801_7;

Selector_2 s1801_7(wires_450_6[1], addr_450_6, addr_positional[7207:7204], addr_1801_7);

wire[31:0] addr_1802_7;

Selector_2 s1802_7(wires_450_6[2], addr_450_6, addr_positional[7211:7208], addr_1802_7);

wire[31:0] addr_1803_7;

Selector_2 s1803_7(wires_450_6[3], addr_450_6, addr_positional[7215:7212], addr_1803_7);

wire[31:0] addr_1804_7;

Selector_2 s1804_7(wires_451_6[0], addr_451_6, addr_positional[7219:7216], addr_1804_7);

wire[31:0] addr_1805_7;

Selector_2 s1805_7(wires_451_6[1], addr_451_6, addr_positional[7223:7220], addr_1805_7);

wire[31:0] addr_1806_7;

Selector_2 s1806_7(wires_451_6[2], addr_451_6, addr_positional[7227:7224], addr_1806_7);

wire[31:0] addr_1807_7;

Selector_2 s1807_7(wires_451_6[3], addr_451_6, addr_positional[7231:7228], addr_1807_7);

wire[31:0] addr_1808_7;

Selector_2 s1808_7(wires_452_6[0], addr_452_6, addr_positional[7235:7232], addr_1808_7);

wire[31:0] addr_1809_7;

Selector_2 s1809_7(wires_452_6[1], addr_452_6, addr_positional[7239:7236], addr_1809_7);

wire[31:0] addr_1810_7;

Selector_2 s1810_7(wires_452_6[2], addr_452_6, addr_positional[7243:7240], addr_1810_7);

wire[31:0] addr_1811_7;

Selector_2 s1811_7(wires_452_6[3], addr_452_6, addr_positional[7247:7244], addr_1811_7);

wire[31:0] addr_1812_7;

Selector_2 s1812_7(wires_453_6[0], addr_453_6, addr_positional[7251:7248], addr_1812_7);

wire[31:0] addr_1813_7;

Selector_2 s1813_7(wires_453_6[1], addr_453_6, addr_positional[7255:7252], addr_1813_7);

wire[31:0] addr_1814_7;

Selector_2 s1814_7(wires_453_6[2], addr_453_6, addr_positional[7259:7256], addr_1814_7);

wire[31:0] addr_1815_7;

Selector_2 s1815_7(wires_453_6[3], addr_453_6, addr_positional[7263:7260], addr_1815_7);

wire[31:0] addr_1816_7;

Selector_2 s1816_7(wires_454_6[0], addr_454_6, addr_positional[7267:7264], addr_1816_7);

wire[31:0] addr_1817_7;

Selector_2 s1817_7(wires_454_6[1], addr_454_6, addr_positional[7271:7268], addr_1817_7);

wire[31:0] addr_1818_7;

Selector_2 s1818_7(wires_454_6[2], addr_454_6, addr_positional[7275:7272], addr_1818_7);

wire[31:0] addr_1819_7;

Selector_2 s1819_7(wires_454_6[3], addr_454_6, addr_positional[7279:7276], addr_1819_7);

wire[31:0] addr_1820_7;

Selector_2 s1820_7(wires_455_6[0], addr_455_6, addr_positional[7283:7280], addr_1820_7);

wire[31:0] addr_1821_7;

Selector_2 s1821_7(wires_455_6[1], addr_455_6, addr_positional[7287:7284], addr_1821_7);

wire[31:0] addr_1822_7;

Selector_2 s1822_7(wires_455_6[2], addr_455_6, addr_positional[7291:7288], addr_1822_7);

wire[31:0] addr_1823_7;

Selector_2 s1823_7(wires_455_6[3], addr_455_6, addr_positional[7295:7292], addr_1823_7);

wire[31:0] addr_1824_7;

Selector_2 s1824_7(wires_456_6[0], addr_456_6, addr_positional[7299:7296], addr_1824_7);

wire[31:0] addr_1825_7;

Selector_2 s1825_7(wires_456_6[1], addr_456_6, addr_positional[7303:7300], addr_1825_7);

wire[31:0] addr_1826_7;

Selector_2 s1826_7(wires_456_6[2], addr_456_6, addr_positional[7307:7304], addr_1826_7);

wire[31:0] addr_1827_7;

Selector_2 s1827_7(wires_456_6[3], addr_456_6, addr_positional[7311:7308], addr_1827_7);

wire[31:0] addr_1828_7;

Selector_2 s1828_7(wires_457_6[0], addr_457_6, addr_positional[7315:7312], addr_1828_7);

wire[31:0] addr_1829_7;

Selector_2 s1829_7(wires_457_6[1], addr_457_6, addr_positional[7319:7316], addr_1829_7);

wire[31:0] addr_1830_7;

Selector_2 s1830_7(wires_457_6[2], addr_457_6, addr_positional[7323:7320], addr_1830_7);

wire[31:0] addr_1831_7;

Selector_2 s1831_7(wires_457_6[3], addr_457_6, addr_positional[7327:7324], addr_1831_7);

wire[31:0] addr_1832_7;

Selector_2 s1832_7(wires_458_6[0], addr_458_6, addr_positional[7331:7328], addr_1832_7);

wire[31:0] addr_1833_7;

Selector_2 s1833_7(wires_458_6[1], addr_458_6, addr_positional[7335:7332], addr_1833_7);

wire[31:0] addr_1834_7;

Selector_2 s1834_7(wires_458_6[2], addr_458_6, addr_positional[7339:7336], addr_1834_7);

wire[31:0] addr_1835_7;

Selector_2 s1835_7(wires_458_6[3], addr_458_6, addr_positional[7343:7340], addr_1835_7);

wire[31:0] addr_1836_7;

Selector_2 s1836_7(wires_459_6[0], addr_459_6, addr_positional[7347:7344], addr_1836_7);

wire[31:0] addr_1837_7;

Selector_2 s1837_7(wires_459_6[1], addr_459_6, addr_positional[7351:7348], addr_1837_7);

wire[31:0] addr_1838_7;

Selector_2 s1838_7(wires_459_6[2], addr_459_6, addr_positional[7355:7352], addr_1838_7);

wire[31:0] addr_1839_7;

Selector_2 s1839_7(wires_459_6[3], addr_459_6, addr_positional[7359:7356], addr_1839_7);

wire[31:0] addr_1840_7;

Selector_2 s1840_7(wires_460_6[0], addr_460_6, addr_positional[7363:7360], addr_1840_7);

wire[31:0] addr_1841_7;

Selector_2 s1841_7(wires_460_6[1], addr_460_6, addr_positional[7367:7364], addr_1841_7);

wire[31:0] addr_1842_7;

Selector_2 s1842_7(wires_460_6[2], addr_460_6, addr_positional[7371:7368], addr_1842_7);

wire[31:0] addr_1843_7;

Selector_2 s1843_7(wires_460_6[3], addr_460_6, addr_positional[7375:7372], addr_1843_7);

wire[31:0] addr_1844_7;

Selector_2 s1844_7(wires_461_6[0], addr_461_6, addr_positional[7379:7376], addr_1844_7);

wire[31:0] addr_1845_7;

Selector_2 s1845_7(wires_461_6[1], addr_461_6, addr_positional[7383:7380], addr_1845_7);

wire[31:0] addr_1846_7;

Selector_2 s1846_7(wires_461_6[2], addr_461_6, addr_positional[7387:7384], addr_1846_7);

wire[31:0] addr_1847_7;

Selector_2 s1847_7(wires_461_6[3], addr_461_6, addr_positional[7391:7388], addr_1847_7);

wire[31:0] addr_1848_7;

Selector_2 s1848_7(wires_462_6[0], addr_462_6, addr_positional[7395:7392], addr_1848_7);

wire[31:0] addr_1849_7;

Selector_2 s1849_7(wires_462_6[1], addr_462_6, addr_positional[7399:7396], addr_1849_7);

wire[31:0] addr_1850_7;

Selector_2 s1850_7(wires_462_6[2], addr_462_6, addr_positional[7403:7400], addr_1850_7);

wire[31:0] addr_1851_7;

Selector_2 s1851_7(wires_462_6[3], addr_462_6, addr_positional[7407:7404], addr_1851_7);

wire[31:0] addr_1852_7;

Selector_2 s1852_7(wires_463_6[0], addr_463_6, addr_positional[7411:7408], addr_1852_7);

wire[31:0] addr_1853_7;

Selector_2 s1853_7(wires_463_6[1], addr_463_6, addr_positional[7415:7412], addr_1853_7);

wire[31:0] addr_1854_7;

Selector_2 s1854_7(wires_463_6[2], addr_463_6, addr_positional[7419:7416], addr_1854_7);

wire[31:0] addr_1855_7;

Selector_2 s1855_7(wires_463_6[3], addr_463_6, addr_positional[7423:7420], addr_1855_7);

wire[31:0] addr_1856_7;

Selector_2 s1856_7(wires_464_6[0], addr_464_6, addr_positional[7427:7424], addr_1856_7);

wire[31:0] addr_1857_7;

Selector_2 s1857_7(wires_464_6[1], addr_464_6, addr_positional[7431:7428], addr_1857_7);

wire[31:0] addr_1858_7;

Selector_2 s1858_7(wires_464_6[2], addr_464_6, addr_positional[7435:7432], addr_1858_7);

wire[31:0] addr_1859_7;

Selector_2 s1859_7(wires_464_6[3], addr_464_6, addr_positional[7439:7436], addr_1859_7);

wire[31:0] addr_1860_7;

Selector_2 s1860_7(wires_465_6[0], addr_465_6, addr_positional[7443:7440], addr_1860_7);

wire[31:0] addr_1861_7;

Selector_2 s1861_7(wires_465_6[1], addr_465_6, addr_positional[7447:7444], addr_1861_7);

wire[31:0] addr_1862_7;

Selector_2 s1862_7(wires_465_6[2], addr_465_6, addr_positional[7451:7448], addr_1862_7);

wire[31:0] addr_1863_7;

Selector_2 s1863_7(wires_465_6[3], addr_465_6, addr_positional[7455:7452], addr_1863_7);

wire[31:0] addr_1864_7;

Selector_2 s1864_7(wires_466_6[0], addr_466_6, addr_positional[7459:7456], addr_1864_7);

wire[31:0] addr_1865_7;

Selector_2 s1865_7(wires_466_6[1], addr_466_6, addr_positional[7463:7460], addr_1865_7);

wire[31:0] addr_1866_7;

Selector_2 s1866_7(wires_466_6[2], addr_466_6, addr_positional[7467:7464], addr_1866_7);

wire[31:0] addr_1867_7;

Selector_2 s1867_7(wires_466_6[3], addr_466_6, addr_positional[7471:7468], addr_1867_7);

wire[31:0] addr_1868_7;

Selector_2 s1868_7(wires_467_6[0], addr_467_6, addr_positional[7475:7472], addr_1868_7);

wire[31:0] addr_1869_7;

Selector_2 s1869_7(wires_467_6[1], addr_467_6, addr_positional[7479:7476], addr_1869_7);

wire[31:0] addr_1870_7;

Selector_2 s1870_7(wires_467_6[2], addr_467_6, addr_positional[7483:7480], addr_1870_7);

wire[31:0] addr_1871_7;

Selector_2 s1871_7(wires_467_6[3], addr_467_6, addr_positional[7487:7484], addr_1871_7);

wire[31:0] addr_1872_7;

Selector_2 s1872_7(wires_468_6[0], addr_468_6, addr_positional[7491:7488], addr_1872_7);

wire[31:0] addr_1873_7;

Selector_2 s1873_7(wires_468_6[1], addr_468_6, addr_positional[7495:7492], addr_1873_7);

wire[31:0] addr_1874_7;

Selector_2 s1874_7(wires_468_6[2], addr_468_6, addr_positional[7499:7496], addr_1874_7);

wire[31:0] addr_1875_7;

Selector_2 s1875_7(wires_468_6[3], addr_468_6, addr_positional[7503:7500], addr_1875_7);

wire[31:0] addr_1876_7;

Selector_2 s1876_7(wires_469_6[0], addr_469_6, addr_positional[7507:7504], addr_1876_7);

wire[31:0] addr_1877_7;

Selector_2 s1877_7(wires_469_6[1], addr_469_6, addr_positional[7511:7508], addr_1877_7);

wire[31:0] addr_1878_7;

Selector_2 s1878_7(wires_469_6[2], addr_469_6, addr_positional[7515:7512], addr_1878_7);

wire[31:0] addr_1879_7;

Selector_2 s1879_7(wires_469_6[3], addr_469_6, addr_positional[7519:7516], addr_1879_7);

wire[31:0] addr_1880_7;

Selector_2 s1880_7(wires_470_6[0], addr_470_6, addr_positional[7523:7520], addr_1880_7);

wire[31:0] addr_1881_7;

Selector_2 s1881_7(wires_470_6[1], addr_470_6, addr_positional[7527:7524], addr_1881_7);

wire[31:0] addr_1882_7;

Selector_2 s1882_7(wires_470_6[2], addr_470_6, addr_positional[7531:7528], addr_1882_7);

wire[31:0] addr_1883_7;

Selector_2 s1883_7(wires_470_6[3], addr_470_6, addr_positional[7535:7532], addr_1883_7);

wire[31:0] addr_1884_7;

Selector_2 s1884_7(wires_471_6[0], addr_471_6, addr_positional[7539:7536], addr_1884_7);

wire[31:0] addr_1885_7;

Selector_2 s1885_7(wires_471_6[1], addr_471_6, addr_positional[7543:7540], addr_1885_7);

wire[31:0] addr_1886_7;

Selector_2 s1886_7(wires_471_6[2], addr_471_6, addr_positional[7547:7544], addr_1886_7);

wire[31:0] addr_1887_7;

Selector_2 s1887_7(wires_471_6[3], addr_471_6, addr_positional[7551:7548], addr_1887_7);

wire[31:0] addr_1888_7;

Selector_2 s1888_7(wires_472_6[0], addr_472_6, addr_positional[7555:7552], addr_1888_7);

wire[31:0] addr_1889_7;

Selector_2 s1889_7(wires_472_6[1], addr_472_6, addr_positional[7559:7556], addr_1889_7);

wire[31:0] addr_1890_7;

Selector_2 s1890_7(wires_472_6[2], addr_472_6, addr_positional[7563:7560], addr_1890_7);

wire[31:0] addr_1891_7;

Selector_2 s1891_7(wires_472_6[3], addr_472_6, addr_positional[7567:7564], addr_1891_7);

wire[31:0] addr_1892_7;

Selector_2 s1892_7(wires_473_6[0], addr_473_6, addr_positional[7571:7568], addr_1892_7);

wire[31:0] addr_1893_7;

Selector_2 s1893_7(wires_473_6[1], addr_473_6, addr_positional[7575:7572], addr_1893_7);

wire[31:0] addr_1894_7;

Selector_2 s1894_7(wires_473_6[2], addr_473_6, addr_positional[7579:7576], addr_1894_7);

wire[31:0] addr_1895_7;

Selector_2 s1895_7(wires_473_6[3], addr_473_6, addr_positional[7583:7580], addr_1895_7);

wire[31:0] addr_1896_7;

Selector_2 s1896_7(wires_474_6[0], addr_474_6, addr_positional[7587:7584], addr_1896_7);

wire[31:0] addr_1897_7;

Selector_2 s1897_7(wires_474_6[1], addr_474_6, addr_positional[7591:7588], addr_1897_7);

wire[31:0] addr_1898_7;

Selector_2 s1898_7(wires_474_6[2], addr_474_6, addr_positional[7595:7592], addr_1898_7);

wire[31:0] addr_1899_7;

Selector_2 s1899_7(wires_474_6[3], addr_474_6, addr_positional[7599:7596], addr_1899_7);

wire[31:0] addr_1900_7;

Selector_2 s1900_7(wires_475_6[0], addr_475_6, addr_positional[7603:7600], addr_1900_7);

wire[31:0] addr_1901_7;

Selector_2 s1901_7(wires_475_6[1], addr_475_6, addr_positional[7607:7604], addr_1901_7);

wire[31:0] addr_1902_7;

Selector_2 s1902_7(wires_475_6[2], addr_475_6, addr_positional[7611:7608], addr_1902_7);

wire[31:0] addr_1903_7;

Selector_2 s1903_7(wires_475_6[3], addr_475_6, addr_positional[7615:7612], addr_1903_7);

wire[31:0] addr_1904_7;

Selector_2 s1904_7(wires_476_6[0], addr_476_6, addr_positional[7619:7616], addr_1904_7);

wire[31:0] addr_1905_7;

Selector_2 s1905_7(wires_476_6[1], addr_476_6, addr_positional[7623:7620], addr_1905_7);

wire[31:0] addr_1906_7;

Selector_2 s1906_7(wires_476_6[2], addr_476_6, addr_positional[7627:7624], addr_1906_7);

wire[31:0] addr_1907_7;

Selector_2 s1907_7(wires_476_6[3], addr_476_6, addr_positional[7631:7628], addr_1907_7);

wire[31:0] addr_1908_7;

Selector_2 s1908_7(wires_477_6[0], addr_477_6, addr_positional[7635:7632], addr_1908_7);

wire[31:0] addr_1909_7;

Selector_2 s1909_7(wires_477_6[1], addr_477_6, addr_positional[7639:7636], addr_1909_7);

wire[31:0] addr_1910_7;

Selector_2 s1910_7(wires_477_6[2], addr_477_6, addr_positional[7643:7640], addr_1910_7);

wire[31:0] addr_1911_7;

Selector_2 s1911_7(wires_477_6[3], addr_477_6, addr_positional[7647:7644], addr_1911_7);

wire[31:0] addr_1912_7;

Selector_2 s1912_7(wires_478_6[0], addr_478_6, addr_positional[7651:7648], addr_1912_7);

wire[31:0] addr_1913_7;

Selector_2 s1913_7(wires_478_6[1], addr_478_6, addr_positional[7655:7652], addr_1913_7);

wire[31:0] addr_1914_7;

Selector_2 s1914_7(wires_478_6[2], addr_478_6, addr_positional[7659:7656], addr_1914_7);

wire[31:0] addr_1915_7;

Selector_2 s1915_7(wires_478_6[3], addr_478_6, addr_positional[7663:7660], addr_1915_7);

wire[31:0] addr_1916_7;

Selector_2 s1916_7(wires_479_6[0], addr_479_6, addr_positional[7667:7664], addr_1916_7);

wire[31:0] addr_1917_7;

Selector_2 s1917_7(wires_479_6[1], addr_479_6, addr_positional[7671:7668], addr_1917_7);

wire[31:0] addr_1918_7;

Selector_2 s1918_7(wires_479_6[2], addr_479_6, addr_positional[7675:7672], addr_1918_7);

wire[31:0] addr_1919_7;

Selector_2 s1919_7(wires_479_6[3], addr_479_6, addr_positional[7679:7676], addr_1919_7);

wire[31:0] addr_1920_7;

Selector_2 s1920_7(wires_480_6[0], addr_480_6, addr_positional[7683:7680], addr_1920_7);

wire[31:0] addr_1921_7;

Selector_2 s1921_7(wires_480_6[1], addr_480_6, addr_positional[7687:7684], addr_1921_7);

wire[31:0] addr_1922_7;

Selector_2 s1922_7(wires_480_6[2], addr_480_6, addr_positional[7691:7688], addr_1922_7);

wire[31:0] addr_1923_7;

Selector_2 s1923_7(wires_480_6[3], addr_480_6, addr_positional[7695:7692], addr_1923_7);

wire[31:0] addr_1924_7;

Selector_2 s1924_7(wires_481_6[0], addr_481_6, addr_positional[7699:7696], addr_1924_7);

wire[31:0] addr_1925_7;

Selector_2 s1925_7(wires_481_6[1], addr_481_6, addr_positional[7703:7700], addr_1925_7);

wire[31:0] addr_1926_7;

Selector_2 s1926_7(wires_481_6[2], addr_481_6, addr_positional[7707:7704], addr_1926_7);

wire[31:0] addr_1927_7;

Selector_2 s1927_7(wires_481_6[3], addr_481_6, addr_positional[7711:7708], addr_1927_7);

wire[31:0] addr_1928_7;

Selector_2 s1928_7(wires_482_6[0], addr_482_6, addr_positional[7715:7712], addr_1928_7);

wire[31:0] addr_1929_7;

Selector_2 s1929_7(wires_482_6[1], addr_482_6, addr_positional[7719:7716], addr_1929_7);

wire[31:0] addr_1930_7;

Selector_2 s1930_7(wires_482_6[2], addr_482_6, addr_positional[7723:7720], addr_1930_7);

wire[31:0] addr_1931_7;

Selector_2 s1931_7(wires_482_6[3], addr_482_6, addr_positional[7727:7724], addr_1931_7);

wire[31:0] addr_1932_7;

Selector_2 s1932_7(wires_483_6[0], addr_483_6, addr_positional[7731:7728], addr_1932_7);

wire[31:0] addr_1933_7;

Selector_2 s1933_7(wires_483_6[1], addr_483_6, addr_positional[7735:7732], addr_1933_7);

wire[31:0] addr_1934_7;

Selector_2 s1934_7(wires_483_6[2], addr_483_6, addr_positional[7739:7736], addr_1934_7);

wire[31:0] addr_1935_7;

Selector_2 s1935_7(wires_483_6[3], addr_483_6, addr_positional[7743:7740], addr_1935_7);

wire[31:0] addr_1936_7;

Selector_2 s1936_7(wires_484_6[0], addr_484_6, addr_positional[7747:7744], addr_1936_7);

wire[31:0] addr_1937_7;

Selector_2 s1937_7(wires_484_6[1], addr_484_6, addr_positional[7751:7748], addr_1937_7);

wire[31:0] addr_1938_7;

Selector_2 s1938_7(wires_484_6[2], addr_484_6, addr_positional[7755:7752], addr_1938_7);

wire[31:0] addr_1939_7;

Selector_2 s1939_7(wires_484_6[3], addr_484_6, addr_positional[7759:7756], addr_1939_7);

wire[31:0] addr_1940_7;

Selector_2 s1940_7(wires_485_6[0], addr_485_6, addr_positional[7763:7760], addr_1940_7);

wire[31:0] addr_1941_7;

Selector_2 s1941_7(wires_485_6[1], addr_485_6, addr_positional[7767:7764], addr_1941_7);

wire[31:0] addr_1942_7;

Selector_2 s1942_7(wires_485_6[2], addr_485_6, addr_positional[7771:7768], addr_1942_7);

wire[31:0] addr_1943_7;

Selector_2 s1943_7(wires_485_6[3], addr_485_6, addr_positional[7775:7772], addr_1943_7);

wire[31:0] addr_1944_7;

Selector_2 s1944_7(wires_486_6[0], addr_486_6, addr_positional[7779:7776], addr_1944_7);

wire[31:0] addr_1945_7;

Selector_2 s1945_7(wires_486_6[1], addr_486_6, addr_positional[7783:7780], addr_1945_7);

wire[31:0] addr_1946_7;

Selector_2 s1946_7(wires_486_6[2], addr_486_6, addr_positional[7787:7784], addr_1946_7);

wire[31:0] addr_1947_7;

Selector_2 s1947_7(wires_486_6[3], addr_486_6, addr_positional[7791:7788], addr_1947_7);

wire[31:0] addr_1948_7;

Selector_2 s1948_7(wires_487_6[0], addr_487_6, addr_positional[7795:7792], addr_1948_7);

wire[31:0] addr_1949_7;

Selector_2 s1949_7(wires_487_6[1], addr_487_6, addr_positional[7799:7796], addr_1949_7);

wire[31:0] addr_1950_7;

Selector_2 s1950_7(wires_487_6[2], addr_487_6, addr_positional[7803:7800], addr_1950_7);

wire[31:0] addr_1951_7;

Selector_2 s1951_7(wires_487_6[3], addr_487_6, addr_positional[7807:7804], addr_1951_7);

wire[31:0] addr_1952_7;

Selector_2 s1952_7(wires_488_6[0], addr_488_6, addr_positional[7811:7808], addr_1952_7);

wire[31:0] addr_1953_7;

Selector_2 s1953_7(wires_488_6[1], addr_488_6, addr_positional[7815:7812], addr_1953_7);

wire[31:0] addr_1954_7;

Selector_2 s1954_7(wires_488_6[2], addr_488_6, addr_positional[7819:7816], addr_1954_7);

wire[31:0] addr_1955_7;

Selector_2 s1955_7(wires_488_6[3], addr_488_6, addr_positional[7823:7820], addr_1955_7);

wire[31:0] addr_1956_7;

Selector_2 s1956_7(wires_489_6[0], addr_489_6, addr_positional[7827:7824], addr_1956_7);

wire[31:0] addr_1957_7;

Selector_2 s1957_7(wires_489_6[1], addr_489_6, addr_positional[7831:7828], addr_1957_7);

wire[31:0] addr_1958_7;

Selector_2 s1958_7(wires_489_6[2], addr_489_6, addr_positional[7835:7832], addr_1958_7);

wire[31:0] addr_1959_7;

Selector_2 s1959_7(wires_489_6[3], addr_489_6, addr_positional[7839:7836], addr_1959_7);

wire[31:0] addr_1960_7;

Selector_2 s1960_7(wires_490_6[0], addr_490_6, addr_positional[7843:7840], addr_1960_7);

wire[31:0] addr_1961_7;

Selector_2 s1961_7(wires_490_6[1], addr_490_6, addr_positional[7847:7844], addr_1961_7);

wire[31:0] addr_1962_7;

Selector_2 s1962_7(wires_490_6[2], addr_490_6, addr_positional[7851:7848], addr_1962_7);

wire[31:0] addr_1963_7;

Selector_2 s1963_7(wires_490_6[3], addr_490_6, addr_positional[7855:7852], addr_1963_7);

wire[31:0] addr_1964_7;

Selector_2 s1964_7(wires_491_6[0], addr_491_6, addr_positional[7859:7856], addr_1964_7);

wire[31:0] addr_1965_7;

Selector_2 s1965_7(wires_491_6[1], addr_491_6, addr_positional[7863:7860], addr_1965_7);

wire[31:0] addr_1966_7;

Selector_2 s1966_7(wires_491_6[2], addr_491_6, addr_positional[7867:7864], addr_1966_7);

wire[31:0] addr_1967_7;

Selector_2 s1967_7(wires_491_6[3], addr_491_6, addr_positional[7871:7868], addr_1967_7);

wire[31:0] addr_1968_7;

Selector_2 s1968_7(wires_492_6[0], addr_492_6, addr_positional[7875:7872], addr_1968_7);

wire[31:0] addr_1969_7;

Selector_2 s1969_7(wires_492_6[1], addr_492_6, addr_positional[7879:7876], addr_1969_7);

wire[31:0] addr_1970_7;

Selector_2 s1970_7(wires_492_6[2], addr_492_6, addr_positional[7883:7880], addr_1970_7);

wire[31:0] addr_1971_7;

Selector_2 s1971_7(wires_492_6[3], addr_492_6, addr_positional[7887:7884], addr_1971_7);

wire[31:0] addr_1972_7;

Selector_2 s1972_7(wires_493_6[0], addr_493_6, addr_positional[7891:7888], addr_1972_7);

wire[31:0] addr_1973_7;

Selector_2 s1973_7(wires_493_6[1], addr_493_6, addr_positional[7895:7892], addr_1973_7);

wire[31:0] addr_1974_7;

Selector_2 s1974_7(wires_493_6[2], addr_493_6, addr_positional[7899:7896], addr_1974_7);

wire[31:0] addr_1975_7;

Selector_2 s1975_7(wires_493_6[3], addr_493_6, addr_positional[7903:7900], addr_1975_7);

wire[31:0] addr_1976_7;

Selector_2 s1976_7(wires_494_6[0], addr_494_6, addr_positional[7907:7904], addr_1976_7);

wire[31:0] addr_1977_7;

Selector_2 s1977_7(wires_494_6[1], addr_494_6, addr_positional[7911:7908], addr_1977_7);

wire[31:0] addr_1978_7;

Selector_2 s1978_7(wires_494_6[2], addr_494_6, addr_positional[7915:7912], addr_1978_7);

wire[31:0] addr_1979_7;

Selector_2 s1979_7(wires_494_6[3], addr_494_6, addr_positional[7919:7916], addr_1979_7);

wire[31:0] addr_1980_7;

Selector_2 s1980_7(wires_495_6[0], addr_495_6, addr_positional[7923:7920], addr_1980_7);

wire[31:0] addr_1981_7;

Selector_2 s1981_7(wires_495_6[1], addr_495_6, addr_positional[7927:7924], addr_1981_7);

wire[31:0] addr_1982_7;

Selector_2 s1982_7(wires_495_6[2], addr_495_6, addr_positional[7931:7928], addr_1982_7);

wire[31:0] addr_1983_7;

Selector_2 s1983_7(wires_495_6[3], addr_495_6, addr_positional[7935:7932], addr_1983_7);

wire[31:0] addr_1984_7;

Selector_2 s1984_7(wires_496_6[0], addr_496_6, addr_positional[7939:7936], addr_1984_7);

wire[31:0] addr_1985_7;

Selector_2 s1985_7(wires_496_6[1], addr_496_6, addr_positional[7943:7940], addr_1985_7);

wire[31:0] addr_1986_7;

Selector_2 s1986_7(wires_496_6[2], addr_496_6, addr_positional[7947:7944], addr_1986_7);

wire[31:0] addr_1987_7;

Selector_2 s1987_7(wires_496_6[3], addr_496_6, addr_positional[7951:7948], addr_1987_7);

wire[31:0] addr_1988_7;

Selector_2 s1988_7(wires_497_6[0], addr_497_6, addr_positional[7955:7952], addr_1988_7);

wire[31:0] addr_1989_7;

Selector_2 s1989_7(wires_497_6[1], addr_497_6, addr_positional[7959:7956], addr_1989_7);

wire[31:0] addr_1990_7;

Selector_2 s1990_7(wires_497_6[2], addr_497_6, addr_positional[7963:7960], addr_1990_7);

wire[31:0] addr_1991_7;

Selector_2 s1991_7(wires_497_6[3], addr_497_6, addr_positional[7967:7964], addr_1991_7);

wire[31:0] addr_1992_7;

Selector_2 s1992_7(wires_498_6[0], addr_498_6, addr_positional[7971:7968], addr_1992_7);

wire[31:0] addr_1993_7;

Selector_2 s1993_7(wires_498_6[1], addr_498_6, addr_positional[7975:7972], addr_1993_7);

wire[31:0] addr_1994_7;

Selector_2 s1994_7(wires_498_6[2], addr_498_6, addr_positional[7979:7976], addr_1994_7);

wire[31:0] addr_1995_7;

Selector_2 s1995_7(wires_498_6[3], addr_498_6, addr_positional[7983:7980], addr_1995_7);

wire[31:0] addr_1996_7;

Selector_2 s1996_7(wires_499_6[0], addr_499_6, addr_positional[7987:7984], addr_1996_7);

wire[31:0] addr_1997_7;

Selector_2 s1997_7(wires_499_6[1], addr_499_6, addr_positional[7991:7988], addr_1997_7);

wire[31:0] addr_1998_7;

Selector_2 s1998_7(wires_499_6[2], addr_499_6, addr_positional[7995:7992], addr_1998_7);

wire[31:0] addr_1999_7;

Selector_2 s1999_7(wires_499_6[3], addr_499_6, addr_positional[7999:7996], addr_1999_7);

wire[31:0] addr_2000_7;

Selector_2 s2000_7(wires_500_6[0], addr_500_6, addr_positional[8003:8000], addr_2000_7);

wire[31:0] addr_2001_7;

Selector_2 s2001_7(wires_500_6[1], addr_500_6, addr_positional[8007:8004], addr_2001_7);

wire[31:0] addr_2002_7;

Selector_2 s2002_7(wires_500_6[2], addr_500_6, addr_positional[8011:8008], addr_2002_7);

wire[31:0] addr_2003_7;

Selector_2 s2003_7(wires_500_6[3], addr_500_6, addr_positional[8015:8012], addr_2003_7);

wire[31:0] addr_2004_7;

Selector_2 s2004_7(wires_501_6[0], addr_501_6, addr_positional[8019:8016], addr_2004_7);

wire[31:0] addr_2005_7;

Selector_2 s2005_7(wires_501_6[1], addr_501_6, addr_positional[8023:8020], addr_2005_7);

wire[31:0] addr_2006_7;

Selector_2 s2006_7(wires_501_6[2], addr_501_6, addr_positional[8027:8024], addr_2006_7);

wire[31:0] addr_2007_7;

Selector_2 s2007_7(wires_501_6[3], addr_501_6, addr_positional[8031:8028], addr_2007_7);

wire[31:0] addr_2008_7;

Selector_2 s2008_7(wires_502_6[0], addr_502_6, addr_positional[8035:8032], addr_2008_7);

wire[31:0] addr_2009_7;

Selector_2 s2009_7(wires_502_6[1], addr_502_6, addr_positional[8039:8036], addr_2009_7);

wire[31:0] addr_2010_7;

Selector_2 s2010_7(wires_502_6[2], addr_502_6, addr_positional[8043:8040], addr_2010_7);

wire[31:0] addr_2011_7;

Selector_2 s2011_7(wires_502_6[3], addr_502_6, addr_positional[8047:8044], addr_2011_7);

wire[31:0] addr_2012_7;

Selector_2 s2012_7(wires_503_6[0], addr_503_6, addr_positional[8051:8048], addr_2012_7);

wire[31:0] addr_2013_7;

Selector_2 s2013_7(wires_503_6[1], addr_503_6, addr_positional[8055:8052], addr_2013_7);

wire[31:0] addr_2014_7;

Selector_2 s2014_7(wires_503_6[2], addr_503_6, addr_positional[8059:8056], addr_2014_7);

wire[31:0] addr_2015_7;

Selector_2 s2015_7(wires_503_6[3], addr_503_6, addr_positional[8063:8060], addr_2015_7);

wire[31:0] addr_2016_7;

Selector_2 s2016_7(wires_504_6[0], addr_504_6, addr_positional[8067:8064], addr_2016_7);

wire[31:0] addr_2017_7;

Selector_2 s2017_7(wires_504_6[1], addr_504_6, addr_positional[8071:8068], addr_2017_7);

wire[31:0] addr_2018_7;

Selector_2 s2018_7(wires_504_6[2], addr_504_6, addr_positional[8075:8072], addr_2018_7);

wire[31:0] addr_2019_7;

Selector_2 s2019_7(wires_504_6[3], addr_504_6, addr_positional[8079:8076], addr_2019_7);

wire[31:0] addr_2020_7;

Selector_2 s2020_7(wires_505_6[0], addr_505_6, addr_positional[8083:8080], addr_2020_7);

wire[31:0] addr_2021_7;

Selector_2 s2021_7(wires_505_6[1], addr_505_6, addr_positional[8087:8084], addr_2021_7);

wire[31:0] addr_2022_7;

Selector_2 s2022_7(wires_505_6[2], addr_505_6, addr_positional[8091:8088], addr_2022_7);

wire[31:0] addr_2023_7;

Selector_2 s2023_7(wires_505_6[3], addr_505_6, addr_positional[8095:8092], addr_2023_7);

wire[31:0] addr_2024_7;

Selector_2 s2024_7(wires_506_6[0], addr_506_6, addr_positional[8099:8096], addr_2024_7);

wire[31:0] addr_2025_7;

Selector_2 s2025_7(wires_506_6[1], addr_506_6, addr_positional[8103:8100], addr_2025_7);

wire[31:0] addr_2026_7;

Selector_2 s2026_7(wires_506_6[2], addr_506_6, addr_positional[8107:8104], addr_2026_7);

wire[31:0] addr_2027_7;

Selector_2 s2027_7(wires_506_6[3], addr_506_6, addr_positional[8111:8108], addr_2027_7);

wire[31:0] addr_2028_7;

Selector_2 s2028_7(wires_507_6[0], addr_507_6, addr_positional[8115:8112], addr_2028_7);

wire[31:0] addr_2029_7;

Selector_2 s2029_7(wires_507_6[1], addr_507_6, addr_positional[8119:8116], addr_2029_7);

wire[31:0] addr_2030_7;

Selector_2 s2030_7(wires_507_6[2], addr_507_6, addr_positional[8123:8120], addr_2030_7);

wire[31:0] addr_2031_7;

Selector_2 s2031_7(wires_507_6[3], addr_507_6, addr_positional[8127:8124], addr_2031_7);

wire[31:0] addr_2032_7;

Selector_2 s2032_7(wires_508_6[0], addr_508_6, addr_positional[8131:8128], addr_2032_7);

wire[31:0] addr_2033_7;

Selector_2 s2033_7(wires_508_6[1], addr_508_6, addr_positional[8135:8132], addr_2033_7);

wire[31:0] addr_2034_7;

Selector_2 s2034_7(wires_508_6[2], addr_508_6, addr_positional[8139:8136], addr_2034_7);

wire[31:0] addr_2035_7;

Selector_2 s2035_7(wires_508_6[3], addr_508_6, addr_positional[8143:8140], addr_2035_7);

wire[31:0] addr_2036_7;

Selector_2 s2036_7(wires_509_6[0], addr_509_6, addr_positional[8147:8144], addr_2036_7);

wire[31:0] addr_2037_7;

Selector_2 s2037_7(wires_509_6[1], addr_509_6, addr_positional[8151:8148], addr_2037_7);

wire[31:0] addr_2038_7;

Selector_2 s2038_7(wires_509_6[2], addr_509_6, addr_positional[8155:8152], addr_2038_7);

wire[31:0] addr_2039_7;

Selector_2 s2039_7(wires_509_6[3], addr_509_6, addr_positional[8159:8156], addr_2039_7);

wire[31:0] addr_2040_7;

Selector_2 s2040_7(wires_510_6[0], addr_510_6, addr_positional[8163:8160], addr_2040_7);

wire[31:0] addr_2041_7;

Selector_2 s2041_7(wires_510_6[1], addr_510_6, addr_positional[8167:8164], addr_2041_7);

wire[31:0] addr_2042_7;

Selector_2 s2042_7(wires_510_6[2], addr_510_6, addr_positional[8171:8168], addr_2042_7);

wire[31:0] addr_2043_7;

Selector_2 s2043_7(wires_510_6[3], addr_510_6, addr_positional[8175:8172], addr_2043_7);

wire[31:0] addr_2044_7;

Selector_2 s2044_7(wires_511_6[0], addr_511_6, addr_positional[8179:8176], addr_2044_7);

wire[31:0] addr_2045_7;

Selector_2 s2045_7(wires_511_6[1], addr_511_6, addr_positional[8183:8180], addr_2045_7);

wire[31:0] addr_2046_7;

Selector_2 s2046_7(wires_511_6[2], addr_511_6, addr_positional[8187:8184], addr_2046_7);

wire[31:0] addr_2047_7;

Selector_2 s2047_7(wires_511_6[3], addr_511_6, addr_positional[8191:8188], addr_2047_7);

wire[31:0] addr_2048_7;

Selector_2 s2048_7(wires_512_6[0], addr_512_6, addr_positional[8195:8192], addr_2048_7);

wire[31:0] addr_2049_7;

Selector_2 s2049_7(wires_512_6[1], addr_512_6, addr_positional[8199:8196], addr_2049_7);

wire[31:0] addr_2050_7;

Selector_2 s2050_7(wires_512_6[2], addr_512_6, addr_positional[8203:8200], addr_2050_7);

wire[31:0] addr_2051_7;

Selector_2 s2051_7(wires_512_6[3], addr_512_6, addr_positional[8207:8204], addr_2051_7);

wire[31:0] addr_2052_7;

Selector_2 s2052_7(wires_513_6[0], addr_513_6, addr_positional[8211:8208], addr_2052_7);

wire[31:0] addr_2053_7;

Selector_2 s2053_7(wires_513_6[1], addr_513_6, addr_positional[8215:8212], addr_2053_7);

wire[31:0] addr_2054_7;

Selector_2 s2054_7(wires_513_6[2], addr_513_6, addr_positional[8219:8216], addr_2054_7);

wire[31:0] addr_2055_7;

Selector_2 s2055_7(wires_513_6[3], addr_513_6, addr_positional[8223:8220], addr_2055_7);

wire[31:0] addr_2056_7;

Selector_2 s2056_7(wires_514_6[0], addr_514_6, addr_positional[8227:8224], addr_2056_7);

wire[31:0] addr_2057_7;

Selector_2 s2057_7(wires_514_6[1], addr_514_6, addr_positional[8231:8228], addr_2057_7);

wire[31:0] addr_2058_7;

Selector_2 s2058_7(wires_514_6[2], addr_514_6, addr_positional[8235:8232], addr_2058_7);

wire[31:0] addr_2059_7;

Selector_2 s2059_7(wires_514_6[3], addr_514_6, addr_positional[8239:8236], addr_2059_7);

wire[31:0] addr_2060_7;

Selector_2 s2060_7(wires_515_6[0], addr_515_6, addr_positional[8243:8240], addr_2060_7);

wire[31:0] addr_2061_7;

Selector_2 s2061_7(wires_515_6[1], addr_515_6, addr_positional[8247:8244], addr_2061_7);

wire[31:0] addr_2062_7;

Selector_2 s2062_7(wires_515_6[2], addr_515_6, addr_positional[8251:8248], addr_2062_7);

wire[31:0] addr_2063_7;

Selector_2 s2063_7(wires_515_6[3], addr_515_6, addr_positional[8255:8252], addr_2063_7);

wire[31:0] addr_2064_7;

Selector_2 s2064_7(wires_516_6[0], addr_516_6, addr_positional[8259:8256], addr_2064_7);

wire[31:0] addr_2065_7;

Selector_2 s2065_7(wires_516_6[1], addr_516_6, addr_positional[8263:8260], addr_2065_7);

wire[31:0] addr_2066_7;

Selector_2 s2066_7(wires_516_6[2], addr_516_6, addr_positional[8267:8264], addr_2066_7);

wire[31:0] addr_2067_7;

Selector_2 s2067_7(wires_516_6[3], addr_516_6, addr_positional[8271:8268], addr_2067_7);

wire[31:0] addr_2068_7;

Selector_2 s2068_7(wires_517_6[0], addr_517_6, addr_positional[8275:8272], addr_2068_7);

wire[31:0] addr_2069_7;

Selector_2 s2069_7(wires_517_6[1], addr_517_6, addr_positional[8279:8276], addr_2069_7);

wire[31:0] addr_2070_7;

Selector_2 s2070_7(wires_517_6[2], addr_517_6, addr_positional[8283:8280], addr_2070_7);

wire[31:0] addr_2071_7;

Selector_2 s2071_7(wires_517_6[3], addr_517_6, addr_positional[8287:8284], addr_2071_7);

wire[31:0] addr_2072_7;

Selector_2 s2072_7(wires_518_6[0], addr_518_6, addr_positional[8291:8288], addr_2072_7);

wire[31:0] addr_2073_7;

Selector_2 s2073_7(wires_518_6[1], addr_518_6, addr_positional[8295:8292], addr_2073_7);

wire[31:0] addr_2074_7;

Selector_2 s2074_7(wires_518_6[2], addr_518_6, addr_positional[8299:8296], addr_2074_7);

wire[31:0] addr_2075_7;

Selector_2 s2075_7(wires_518_6[3], addr_518_6, addr_positional[8303:8300], addr_2075_7);

wire[31:0] addr_2076_7;

Selector_2 s2076_7(wires_519_6[0], addr_519_6, addr_positional[8307:8304], addr_2076_7);

wire[31:0] addr_2077_7;

Selector_2 s2077_7(wires_519_6[1], addr_519_6, addr_positional[8311:8308], addr_2077_7);

wire[31:0] addr_2078_7;

Selector_2 s2078_7(wires_519_6[2], addr_519_6, addr_positional[8315:8312], addr_2078_7);

wire[31:0] addr_2079_7;

Selector_2 s2079_7(wires_519_6[3], addr_519_6, addr_positional[8319:8316], addr_2079_7);

wire[31:0] addr_2080_7;

Selector_2 s2080_7(wires_520_6[0], addr_520_6, addr_positional[8323:8320], addr_2080_7);

wire[31:0] addr_2081_7;

Selector_2 s2081_7(wires_520_6[1], addr_520_6, addr_positional[8327:8324], addr_2081_7);

wire[31:0] addr_2082_7;

Selector_2 s2082_7(wires_520_6[2], addr_520_6, addr_positional[8331:8328], addr_2082_7);

wire[31:0] addr_2083_7;

Selector_2 s2083_7(wires_520_6[3], addr_520_6, addr_positional[8335:8332], addr_2083_7);

wire[31:0] addr_2084_7;

Selector_2 s2084_7(wires_521_6[0], addr_521_6, addr_positional[8339:8336], addr_2084_7);

wire[31:0] addr_2085_7;

Selector_2 s2085_7(wires_521_6[1], addr_521_6, addr_positional[8343:8340], addr_2085_7);

wire[31:0] addr_2086_7;

Selector_2 s2086_7(wires_521_6[2], addr_521_6, addr_positional[8347:8344], addr_2086_7);

wire[31:0] addr_2087_7;

Selector_2 s2087_7(wires_521_6[3], addr_521_6, addr_positional[8351:8348], addr_2087_7);

wire[31:0] addr_2088_7;

Selector_2 s2088_7(wires_522_6[0], addr_522_6, addr_positional[8355:8352], addr_2088_7);

wire[31:0] addr_2089_7;

Selector_2 s2089_7(wires_522_6[1], addr_522_6, addr_positional[8359:8356], addr_2089_7);

wire[31:0] addr_2090_7;

Selector_2 s2090_7(wires_522_6[2], addr_522_6, addr_positional[8363:8360], addr_2090_7);

wire[31:0] addr_2091_7;

Selector_2 s2091_7(wires_522_6[3], addr_522_6, addr_positional[8367:8364], addr_2091_7);

wire[31:0] addr_2092_7;

Selector_2 s2092_7(wires_523_6[0], addr_523_6, addr_positional[8371:8368], addr_2092_7);

wire[31:0] addr_2093_7;

Selector_2 s2093_7(wires_523_6[1], addr_523_6, addr_positional[8375:8372], addr_2093_7);

wire[31:0] addr_2094_7;

Selector_2 s2094_7(wires_523_6[2], addr_523_6, addr_positional[8379:8376], addr_2094_7);

wire[31:0] addr_2095_7;

Selector_2 s2095_7(wires_523_6[3], addr_523_6, addr_positional[8383:8380], addr_2095_7);

wire[31:0] addr_2096_7;

Selector_2 s2096_7(wires_524_6[0], addr_524_6, addr_positional[8387:8384], addr_2096_7);

wire[31:0] addr_2097_7;

Selector_2 s2097_7(wires_524_6[1], addr_524_6, addr_positional[8391:8388], addr_2097_7);

wire[31:0] addr_2098_7;

Selector_2 s2098_7(wires_524_6[2], addr_524_6, addr_positional[8395:8392], addr_2098_7);

wire[31:0] addr_2099_7;

Selector_2 s2099_7(wires_524_6[3], addr_524_6, addr_positional[8399:8396], addr_2099_7);

wire[31:0] addr_2100_7;

Selector_2 s2100_7(wires_525_6[0], addr_525_6, addr_positional[8403:8400], addr_2100_7);

wire[31:0] addr_2101_7;

Selector_2 s2101_7(wires_525_6[1], addr_525_6, addr_positional[8407:8404], addr_2101_7);

wire[31:0] addr_2102_7;

Selector_2 s2102_7(wires_525_6[2], addr_525_6, addr_positional[8411:8408], addr_2102_7);

wire[31:0] addr_2103_7;

Selector_2 s2103_7(wires_525_6[3], addr_525_6, addr_positional[8415:8412], addr_2103_7);

wire[31:0] addr_2104_7;

Selector_2 s2104_7(wires_526_6[0], addr_526_6, addr_positional[8419:8416], addr_2104_7);

wire[31:0] addr_2105_7;

Selector_2 s2105_7(wires_526_6[1], addr_526_6, addr_positional[8423:8420], addr_2105_7);

wire[31:0] addr_2106_7;

Selector_2 s2106_7(wires_526_6[2], addr_526_6, addr_positional[8427:8424], addr_2106_7);

wire[31:0] addr_2107_7;

Selector_2 s2107_7(wires_526_6[3], addr_526_6, addr_positional[8431:8428], addr_2107_7);

wire[31:0] addr_2108_7;

Selector_2 s2108_7(wires_527_6[0], addr_527_6, addr_positional[8435:8432], addr_2108_7);

wire[31:0] addr_2109_7;

Selector_2 s2109_7(wires_527_6[1], addr_527_6, addr_positional[8439:8436], addr_2109_7);

wire[31:0] addr_2110_7;

Selector_2 s2110_7(wires_527_6[2], addr_527_6, addr_positional[8443:8440], addr_2110_7);

wire[31:0] addr_2111_7;

Selector_2 s2111_7(wires_527_6[3], addr_527_6, addr_positional[8447:8444], addr_2111_7);

wire[31:0] addr_2112_7;

Selector_2 s2112_7(wires_528_6[0], addr_528_6, addr_positional[8451:8448], addr_2112_7);

wire[31:0] addr_2113_7;

Selector_2 s2113_7(wires_528_6[1], addr_528_6, addr_positional[8455:8452], addr_2113_7);

wire[31:0] addr_2114_7;

Selector_2 s2114_7(wires_528_6[2], addr_528_6, addr_positional[8459:8456], addr_2114_7);

wire[31:0] addr_2115_7;

Selector_2 s2115_7(wires_528_6[3], addr_528_6, addr_positional[8463:8460], addr_2115_7);

wire[31:0] addr_2116_7;

Selector_2 s2116_7(wires_529_6[0], addr_529_6, addr_positional[8467:8464], addr_2116_7);

wire[31:0] addr_2117_7;

Selector_2 s2117_7(wires_529_6[1], addr_529_6, addr_positional[8471:8468], addr_2117_7);

wire[31:0] addr_2118_7;

Selector_2 s2118_7(wires_529_6[2], addr_529_6, addr_positional[8475:8472], addr_2118_7);

wire[31:0] addr_2119_7;

Selector_2 s2119_7(wires_529_6[3], addr_529_6, addr_positional[8479:8476], addr_2119_7);

wire[31:0] addr_2120_7;

Selector_2 s2120_7(wires_530_6[0], addr_530_6, addr_positional[8483:8480], addr_2120_7);

wire[31:0] addr_2121_7;

Selector_2 s2121_7(wires_530_6[1], addr_530_6, addr_positional[8487:8484], addr_2121_7);

wire[31:0] addr_2122_7;

Selector_2 s2122_7(wires_530_6[2], addr_530_6, addr_positional[8491:8488], addr_2122_7);

wire[31:0] addr_2123_7;

Selector_2 s2123_7(wires_530_6[3], addr_530_6, addr_positional[8495:8492], addr_2123_7);

wire[31:0] addr_2124_7;

Selector_2 s2124_7(wires_531_6[0], addr_531_6, addr_positional[8499:8496], addr_2124_7);

wire[31:0] addr_2125_7;

Selector_2 s2125_7(wires_531_6[1], addr_531_6, addr_positional[8503:8500], addr_2125_7);

wire[31:0] addr_2126_7;

Selector_2 s2126_7(wires_531_6[2], addr_531_6, addr_positional[8507:8504], addr_2126_7);

wire[31:0] addr_2127_7;

Selector_2 s2127_7(wires_531_6[3], addr_531_6, addr_positional[8511:8508], addr_2127_7);

wire[31:0] addr_2128_7;

Selector_2 s2128_7(wires_532_6[0], addr_532_6, addr_positional[8515:8512], addr_2128_7);

wire[31:0] addr_2129_7;

Selector_2 s2129_7(wires_532_6[1], addr_532_6, addr_positional[8519:8516], addr_2129_7);

wire[31:0] addr_2130_7;

Selector_2 s2130_7(wires_532_6[2], addr_532_6, addr_positional[8523:8520], addr_2130_7);

wire[31:0] addr_2131_7;

Selector_2 s2131_7(wires_532_6[3], addr_532_6, addr_positional[8527:8524], addr_2131_7);

wire[31:0] addr_2132_7;

Selector_2 s2132_7(wires_533_6[0], addr_533_6, addr_positional[8531:8528], addr_2132_7);

wire[31:0] addr_2133_7;

Selector_2 s2133_7(wires_533_6[1], addr_533_6, addr_positional[8535:8532], addr_2133_7);

wire[31:0] addr_2134_7;

Selector_2 s2134_7(wires_533_6[2], addr_533_6, addr_positional[8539:8536], addr_2134_7);

wire[31:0] addr_2135_7;

Selector_2 s2135_7(wires_533_6[3], addr_533_6, addr_positional[8543:8540], addr_2135_7);

wire[31:0] addr_2136_7;

Selector_2 s2136_7(wires_534_6[0], addr_534_6, addr_positional[8547:8544], addr_2136_7);

wire[31:0] addr_2137_7;

Selector_2 s2137_7(wires_534_6[1], addr_534_6, addr_positional[8551:8548], addr_2137_7);

wire[31:0] addr_2138_7;

Selector_2 s2138_7(wires_534_6[2], addr_534_6, addr_positional[8555:8552], addr_2138_7);

wire[31:0] addr_2139_7;

Selector_2 s2139_7(wires_534_6[3], addr_534_6, addr_positional[8559:8556], addr_2139_7);

wire[31:0] addr_2140_7;

Selector_2 s2140_7(wires_535_6[0], addr_535_6, addr_positional[8563:8560], addr_2140_7);

wire[31:0] addr_2141_7;

Selector_2 s2141_7(wires_535_6[1], addr_535_6, addr_positional[8567:8564], addr_2141_7);

wire[31:0] addr_2142_7;

Selector_2 s2142_7(wires_535_6[2], addr_535_6, addr_positional[8571:8568], addr_2142_7);

wire[31:0] addr_2143_7;

Selector_2 s2143_7(wires_535_6[3], addr_535_6, addr_positional[8575:8572], addr_2143_7);

wire[31:0] addr_2144_7;

Selector_2 s2144_7(wires_536_6[0], addr_536_6, addr_positional[8579:8576], addr_2144_7);

wire[31:0] addr_2145_7;

Selector_2 s2145_7(wires_536_6[1], addr_536_6, addr_positional[8583:8580], addr_2145_7);

wire[31:0] addr_2146_7;

Selector_2 s2146_7(wires_536_6[2], addr_536_6, addr_positional[8587:8584], addr_2146_7);

wire[31:0] addr_2147_7;

Selector_2 s2147_7(wires_536_6[3], addr_536_6, addr_positional[8591:8588], addr_2147_7);

wire[31:0] addr_2148_7;

Selector_2 s2148_7(wires_537_6[0], addr_537_6, addr_positional[8595:8592], addr_2148_7);

wire[31:0] addr_2149_7;

Selector_2 s2149_7(wires_537_6[1], addr_537_6, addr_positional[8599:8596], addr_2149_7);

wire[31:0] addr_2150_7;

Selector_2 s2150_7(wires_537_6[2], addr_537_6, addr_positional[8603:8600], addr_2150_7);

wire[31:0] addr_2151_7;

Selector_2 s2151_7(wires_537_6[3], addr_537_6, addr_positional[8607:8604], addr_2151_7);

wire[31:0] addr_2152_7;

Selector_2 s2152_7(wires_538_6[0], addr_538_6, addr_positional[8611:8608], addr_2152_7);

wire[31:0] addr_2153_7;

Selector_2 s2153_7(wires_538_6[1], addr_538_6, addr_positional[8615:8612], addr_2153_7);

wire[31:0] addr_2154_7;

Selector_2 s2154_7(wires_538_6[2], addr_538_6, addr_positional[8619:8616], addr_2154_7);

wire[31:0] addr_2155_7;

Selector_2 s2155_7(wires_538_6[3], addr_538_6, addr_positional[8623:8620], addr_2155_7);

wire[31:0] addr_2156_7;

Selector_2 s2156_7(wires_539_6[0], addr_539_6, addr_positional[8627:8624], addr_2156_7);

wire[31:0] addr_2157_7;

Selector_2 s2157_7(wires_539_6[1], addr_539_6, addr_positional[8631:8628], addr_2157_7);

wire[31:0] addr_2158_7;

Selector_2 s2158_7(wires_539_6[2], addr_539_6, addr_positional[8635:8632], addr_2158_7);

wire[31:0] addr_2159_7;

Selector_2 s2159_7(wires_539_6[3], addr_539_6, addr_positional[8639:8636], addr_2159_7);

wire[31:0] addr_2160_7;

Selector_2 s2160_7(wires_540_6[0], addr_540_6, addr_positional[8643:8640], addr_2160_7);

wire[31:0] addr_2161_7;

Selector_2 s2161_7(wires_540_6[1], addr_540_6, addr_positional[8647:8644], addr_2161_7);

wire[31:0] addr_2162_7;

Selector_2 s2162_7(wires_540_6[2], addr_540_6, addr_positional[8651:8648], addr_2162_7);

wire[31:0] addr_2163_7;

Selector_2 s2163_7(wires_540_6[3], addr_540_6, addr_positional[8655:8652], addr_2163_7);

wire[31:0] addr_2164_7;

Selector_2 s2164_7(wires_541_6[0], addr_541_6, addr_positional[8659:8656], addr_2164_7);

wire[31:0] addr_2165_7;

Selector_2 s2165_7(wires_541_6[1], addr_541_6, addr_positional[8663:8660], addr_2165_7);

wire[31:0] addr_2166_7;

Selector_2 s2166_7(wires_541_6[2], addr_541_6, addr_positional[8667:8664], addr_2166_7);

wire[31:0] addr_2167_7;

Selector_2 s2167_7(wires_541_6[3], addr_541_6, addr_positional[8671:8668], addr_2167_7);

wire[31:0] addr_2168_7;

Selector_2 s2168_7(wires_542_6[0], addr_542_6, addr_positional[8675:8672], addr_2168_7);

wire[31:0] addr_2169_7;

Selector_2 s2169_7(wires_542_6[1], addr_542_6, addr_positional[8679:8676], addr_2169_7);

wire[31:0] addr_2170_7;

Selector_2 s2170_7(wires_542_6[2], addr_542_6, addr_positional[8683:8680], addr_2170_7);

wire[31:0] addr_2171_7;

Selector_2 s2171_7(wires_542_6[3], addr_542_6, addr_positional[8687:8684], addr_2171_7);

wire[31:0] addr_2172_7;

Selector_2 s2172_7(wires_543_6[0], addr_543_6, addr_positional[8691:8688], addr_2172_7);

wire[31:0] addr_2173_7;

Selector_2 s2173_7(wires_543_6[1], addr_543_6, addr_positional[8695:8692], addr_2173_7);

wire[31:0] addr_2174_7;

Selector_2 s2174_7(wires_543_6[2], addr_543_6, addr_positional[8699:8696], addr_2174_7);

wire[31:0] addr_2175_7;

Selector_2 s2175_7(wires_543_6[3], addr_543_6, addr_positional[8703:8700], addr_2175_7);

wire[31:0] addr_2176_7;

Selector_2 s2176_7(wires_544_6[0], addr_544_6, addr_positional[8707:8704], addr_2176_7);

wire[31:0] addr_2177_7;

Selector_2 s2177_7(wires_544_6[1], addr_544_6, addr_positional[8711:8708], addr_2177_7);

wire[31:0] addr_2178_7;

Selector_2 s2178_7(wires_544_6[2], addr_544_6, addr_positional[8715:8712], addr_2178_7);

wire[31:0] addr_2179_7;

Selector_2 s2179_7(wires_544_6[3], addr_544_6, addr_positional[8719:8716], addr_2179_7);

wire[31:0] addr_2180_7;

Selector_2 s2180_7(wires_545_6[0], addr_545_6, addr_positional[8723:8720], addr_2180_7);

wire[31:0] addr_2181_7;

Selector_2 s2181_7(wires_545_6[1], addr_545_6, addr_positional[8727:8724], addr_2181_7);

wire[31:0] addr_2182_7;

Selector_2 s2182_7(wires_545_6[2], addr_545_6, addr_positional[8731:8728], addr_2182_7);

wire[31:0] addr_2183_7;

Selector_2 s2183_7(wires_545_6[3], addr_545_6, addr_positional[8735:8732], addr_2183_7);

wire[31:0] addr_2184_7;

Selector_2 s2184_7(wires_546_6[0], addr_546_6, addr_positional[8739:8736], addr_2184_7);

wire[31:0] addr_2185_7;

Selector_2 s2185_7(wires_546_6[1], addr_546_6, addr_positional[8743:8740], addr_2185_7);

wire[31:0] addr_2186_7;

Selector_2 s2186_7(wires_546_6[2], addr_546_6, addr_positional[8747:8744], addr_2186_7);

wire[31:0] addr_2187_7;

Selector_2 s2187_7(wires_546_6[3], addr_546_6, addr_positional[8751:8748], addr_2187_7);

wire[31:0] addr_2188_7;

Selector_2 s2188_7(wires_547_6[0], addr_547_6, addr_positional[8755:8752], addr_2188_7);

wire[31:0] addr_2189_7;

Selector_2 s2189_7(wires_547_6[1], addr_547_6, addr_positional[8759:8756], addr_2189_7);

wire[31:0] addr_2190_7;

Selector_2 s2190_7(wires_547_6[2], addr_547_6, addr_positional[8763:8760], addr_2190_7);

wire[31:0] addr_2191_7;

Selector_2 s2191_7(wires_547_6[3], addr_547_6, addr_positional[8767:8764], addr_2191_7);

wire[31:0] addr_2192_7;

Selector_2 s2192_7(wires_548_6[0], addr_548_6, addr_positional[8771:8768], addr_2192_7);

wire[31:0] addr_2193_7;

Selector_2 s2193_7(wires_548_6[1], addr_548_6, addr_positional[8775:8772], addr_2193_7);

wire[31:0] addr_2194_7;

Selector_2 s2194_7(wires_548_6[2], addr_548_6, addr_positional[8779:8776], addr_2194_7);

wire[31:0] addr_2195_7;

Selector_2 s2195_7(wires_548_6[3], addr_548_6, addr_positional[8783:8780], addr_2195_7);

wire[31:0] addr_2196_7;

Selector_2 s2196_7(wires_549_6[0], addr_549_6, addr_positional[8787:8784], addr_2196_7);

wire[31:0] addr_2197_7;

Selector_2 s2197_7(wires_549_6[1], addr_549_6, addr_positional[8791:8788], addr_2197_7);

wire[31:0] addr_2198_7;

Selector_2 s2198_7(wires_549_6[2], addr_549_6, addr_positional[8795:8792], addr_2198_7);

wire[31:0] addr_2199_7;

Selector_2 s2199_7(wires_549_6[3], addr_549_6, addr_positional[8799:8796], addr_2199_7);

wire[31:0] addr_2200_7;

Selector_2 s2200_7(wires_550_6[0], addr_550_6, addr_positional[8803:8800], addr_2200_7);

wire[31:0] addr_2201_7;

Selector_2 s2201_7(wires_550_6[1], addr_550_6, addr_positional[8807:8804], addr_2201_7);

wire[31:0] addr_2202_7;

Selector_2 s2202_7(wires_550_6[2], addr_550_6, addr_positional[8811:8808], addr_2202_7);

wire[31:0] addr_2203_7;

Selector_2 s2203_7(wires_550_6[3], addr_550_6, addr_positional[8815:8812], addr_2203_7);

wire[31:0] addr_2204_7;

Selector_2 s2204_7(wires_551_6[0], addr_551_6, addr_positional[8819:8816], addr_2204_7);

wire[31:0] addr_2205_7;

Selector_2 s2205_7(wires_551_6[1], addr_551_6, addr_positional[8823:8820], addr_2205_7);

wire[31:0] addr_2206_7;

Selector_2 s2206_7(wires_551_6[2], addr_551_6, addr_positional[8827:8824], addr_2206_7);

wire[31:0] addr_2207_7;

Selector_2 s2207_7(wires_551_6[3], addr_551_6, addr_positional[8831:8828], addr_2207_7);

wire[31:0] addr_2208_7;

Selector_2 s2208_7(wires_552_6[0], addr_552_6, addr_positional[8835:8832], addr_2208_7);

wire[31:0] addr_2209_7;

Selector_2 s2209_7(wires_552_6[1], addr_552_6, addr_positional[8839:8836], addr_2209_7);

wire[31:0] addr_2210_7;

Selector_2 s2210_7(wires_552_6[2], addr_552_6, addr_positional[8843:8840], addr_2210_7);

wire[31:0] addr_2211_7;

Selector_2 s2211_7(wires_552_6[3], addr_552_6, addr_positional[8847:8844], addr_2211_7);

wire[31:0] addr_2212_7;

Selector_2 s2212_7(wires_553_6[0], addr_553_6, addr_positional[8851:8848], addr_2212_7);

wire[31:0] addr_2213_7;

Selector_2 s2213_7(wires_553_6[1], addr_553_6, addr_positional[8855:8852], addr_2213_7);

wire[31:0] addr_2214_7;

Selector_2 s2214_7(wires_553_6[2], addr_553_6, addr_positional[8859:8856], addr_2214_7);

wire[31:0] addr_2215_7;

Selector_2 s2215_7(wires_553_6[3], addr_553_6, addr_positional[8863:8860], addr_2215_7);

wire[31:0] addr_2216_7;

Selector_2 s2216_7(wires_554_6[0], addr_554_6, addr_positional[8867:8864], addr_2216_7);

wire[31:0] addr_2217_7;

Selector_2 s2217_7(wires_554_6[1], addr_554_6, addr_positional[8871:8868], addr_2217_7);

wire[31:0] addr_2218_7;

Selector_2 s2218_7(wires_554_6[2], addr_554_6, addr_positional[8875:8872], addr_2218_7);

wire[31:0] addr_2219_7;

Selector_2 s2219_7(wires_554_6[3], addr_554_6, addr_positional[8879:8876], addr_2219_7);

wire[31:0] addr_2220_7;

Selector_2 s2220_7(wires_555_6[0], addr_555_6, addr_positional[8883:8880], addr_2220_7);

wire[31:0] addr_2221_7;

Selector_2 s2221_7(wires_555_6[1], addr_555_6, addr_positional[8887:8884], addr_2221_7);

wire[31:0] addr_2222_7;

Selector_2 s2222_7(wires_555_6[2], addr_555_6, addr_positional[8891:8888], addr_2222_7);

wire[31:0] addr_2223_7;

Selector_2 s2223_7(wires_555_6[3], addr_555_6, addr_positional[8895:8892], addr_2223_7);

wire[31:0] addr_2224_7;

Selector_2 s2224_7(wires_556_6[0], addr_556_6, addr_positional[8899:8896], addr_2224_7);

wire[31:0] addr_2225_7;

Selector_2 s2225_7(wires_556_6[1], addr_556_6, addr_positional[8903:8900], addr_2225_7);

wire[31:0] addr_2226_7;

Selector_2 s2226_7(wires_556_6[2], addr_556_6, addr_positional[8907:8904], addr_2226_7);

wire[31:0] addr_2227_7;

Selector_2 s2227_7(wires_556_6[3], addr_556_6, addr_positional[8911:8908], addr_2227_7);

wire[31:0] addr_2228_7;

Selector_2 s2228_7(wires_557_6[0], addr_557_6, addr_positional[8915:8912], addr_2228_7);

wire[31:0] addr_2229_7;

Selector_2 s2229_7(wires_557_6[1], addr_557_6, addr_positional[8919:8916], addr_2229_7);

wire[31:0] addr_2230_7;

Selector_2 s2230_7(wires_557_6[2], addr_557_6, addr_positional[8923:8920], addr_2230_7);

wire[31:0] addr_2231_7;

Selector_2 s2231_7(wires_557_6[3], addr_557_6, addr_positional[8927:8924], addr_2231_7);

wire[31:0] addr_2232_7;

Selector_2 s2232_7(wires_558_6[0], addr_558_6, addr_positional[8931:8928], addr_2232_7);

wire[31:0] addr_2233_7;

Selector_2 s2233_7(wires_558_6[1], addr_558_6, addr_positional[8935:8932], addr_2233_7);

wire[31:0] addr_2234_7;

Selector_2 s2234_7(wires_558_6[2], addr_558_6, addr_positional[8939:8936], addr_2234_7);

wire[31:0] addr_2235_7;

Selector_2 s2235_7(wires_558_6[3], addr_558_6, addr_positional[8943:8940], addr_2235_7);

wire[31:0] addr_2236_7;

Selector_2 s2236_7(wires_559_6[0], addr_559_6, addr_positional[8947:8944], addr_2236_7);

wire[31:0] addr_2237_7;

Selector_2 s2237_7(wires_559_6[1], addr_559_6, addr_positional[8951:8948], addr_2237_7);

wire[31:0] addr_2238_7;

Selector_2 s2238_7(wires_559_6[2], addr_559_6, addr_positional[8955:8952], addr_2238_7);

wire[31:0] addr_2239_7;

Selector_2 s2239_7(wires_559_6[3], addr_559_6, addr_positional[8959:8956], addr_2239_7);

wire[31:0] addr_2240_7;

Selector_2 s2240_7(wires_560_6[0], addr_560_6, addr_positional[8963:8960], addr_2240_7);

wire[31:0] addr_2241_7;

Selector_2 s2241_7(wires_560_6[1], addr_560_6, addr_positional[8967:8964], addr_2241_7);

wire[31:0] addr_2242_7;

Selector_2 s2242_7(wires_560_6[2], addr_560_6, addr_positional[8971:8968], addr_2242_7);

wire[31:0] addr_2243_7;

Selector_2 s2243_7(wires_560_6[3], addr_560_6, addr_positional[8975:8972], addr_2243_7);

wire[31:0] addr_2244_7;

Selector_2 s2244_7(wires_561_6[0], addr_561_6, addr_positional[8979:8976], addr_2244_7);

wire[31:0] addr_2245_7;

Selector_2 s2245_7(wires_561_6[1], addr_561_6, addr_positional[8983:8980], addr_2245_7);

wire[31:0] addr_2246_7;

Selector_2 s2246_7(wires_561_6[2], addr_561_6, addr_positional[8987:8984], addr_2246_7);

wire[31:0] addr_2247_7;

Selector_2 s2247_7(wires_561_6[3], addr_561_6, addr_positional[8991:8988], addr_2247_7);

wire[31:0] addr_2248_7;

Selector_2 s2248_7(wires_562_6[0], addr_562_6, addr_positional[8995:8992], addr_2248_7);

wire[31:0] addr_2249_7;

Selector_2 s2249_7(wires_562_6[1], addr_562_6, addr_positional[8999:8996], addr_2249_7);

wire[31:0] addr_2250_7;

Selector_2 s2250_7(wires_562_6[2], addr_562_6, addr_positional[9003:9000], addr_2250_7);

wire[31:0] addr_2251_7;

Selector_2 s2251_7(wires_562_6[3], addr_562_6, addr_positional[9007:9004], addr_2251_7);

wire[31:0] addr_2252_7;

Selector_2 s2252_7(wires_563_6[0], addr_563_6, addr_positional[9011:9008], addr_2252_7);

wire[31:0] addr_2253_7;

Selector_2 s2253_7(wires_563_6[1], addr_563_6, addr_positional[9015:9012], addr_2253_7);

wire[31:0] addr_2254_7;

Selector_2 s2254_7(wires_563_6[2], addr_563_6, addr_positional[9019:9016], addr_2254_7);

wire[31:0] addr_2255_7;

Selector_2 s2255_7(wires_563_6[3], addr_563_6, addr_positional[9023:9020], addr_2255_7);

wire[31:0] addr_2256_7;

Selector_2 s2256_7(wires_564_6[0], addr_564_6, addr_positional[9027:9024], addr_2256_7);

wire[31:0] addr_2257_7;

Selector_2 s2257_7(wires_564_6[1], addr_564_6, addr_positional[9031:9028], addr_2257_7);

wire[31:0] addr_2258_7;

Selector_2 s2258_7(wires_564_6[2], addr_564_6, addr_positional[9035:9032], addr_2258_7);

wire[31:0] addr_2259_7;

Selector_2 s2259_7(wires_564_6[3], addr_564_6, addr_positional[9039:9036], addr_2259_7);

wire[31:0] addr_2260_7;

Selector_2 s2260_7(wires_565_6[0], addr_565_6, addr_positional[9043:9040], addr_2260_7);

wire[31:0] addr_2261_7;

Selector_2 s2261_7(wires_565_6[1], addr_565_6, addr_positional[9047:9044], addr_2261_7);

wire[31:0] addr_2262_7;

Selector_2 s2262_7(wires_565_6[2], addr_565_6, addr_positional[9051:9048], addr_2262_7);

wire[31:0] addr_2263_7;

Selector_2 s2263_7(wires_565_6[3], addr_565_6, addr_positional[9055:9052], addr_2263_7);

wire[31:0] addr_2264_7;

Selector_2 s2264_7(wires_566_6[0], addr_566_6, addr_positional[9059:9056], addr_2264_7);

wire[31:0] addr_2265_7;

Selector_2 s2265_7(wires_566_6[1], addr_566_6, addr_positional[9063:9060], addr_2265_7);

wire[31:0] addr_2266_7;

Selector_2 s2266_7(wires_566_6[2], addr_566_6, addr_positional[9067:9064], addr_2266_7);

wire[31:0] addr_2267_7;

Selector_2 s2267_7(wires_566_6[3], addr_566_6, addr_positional[9071:9068], addr_2267_7);

wire[31:0] addr_2268_7;

Selector_2 s2268_7(wires_567_6[0], addr_567_6, addr_positional[9075:9072], addr_2268_7);

wire[31:0] addr_2269_7;

Selector_2 s2269_7(wires_567_6[1], addr_567_6, addr_positional[9079:9076], addr_2269_7);

wire[31:0] addr_2270_7;

Selector_2 s2270_7(wires_567_6[2], addr_567_6, addr_positional[9083:9080], addr_2270_7);

wire[31:0] addr_2271_7;

Selector_2 s2271_7(wires_567_6[3], addr_567_6, addr_positional[9087:9084], addr_2271_7);

wire[31:0] addr_2272_7;

Selector_2 s2272_7(wires_568_6[0], addr_568_6, addr_positional[9091:9088], addr_2272_7);

wire[31:0] addr_2273_7;

Selector_2 s2273_7(wires_568_6[1], addr_568_6, addr_positional[9095:9092], addr_2273_7);

wire[31:0] addr_2274_7;

Selector_2 s2274_7(wires_568_6[2], addr_568_6, addr_positional[9099:9096], addr_2274_7);

wire[31:0] addr_2275_7;

Selector_2 s2275_7(wires_568_6[3], addr_568_6, addr_positional[9103:9100], addr_2275_7);

wire[31:0] addr_2276_7;

Selector_2 s2276_7(wires_569_6[0], addr_569_6, addr_positional[9107:9104], addr_2276_7);

wire[31:0] addr_2277_7;

Selector_2 s2277_7(wires_569_6[1], addr_569_6, addr_positional[9111:9108], addr_2277_7);

wire[31:0] addr_2278_7;

Selector_2 s2278_7(wires_569_6[2], addr_569_6, addr_positional[9115:9112], addr_2278_7);

wire[31:0] addr_2279_7;

Selector_2 s2279_7(wires_569_6[3], addr_569_6, addr_positional[9119:9116], addr_2279_7);

wire[31:0] addr_2280_7;

Selector_2 s2280_7(wires_570_6[0], addr_570_6, addr_positional[9123:9120], addr_2280_7);

wire[31:0] addr_2281_7;

Selector_2 s2281_7(wires_570_6[1], addr_570_6, addr_positional[9127:9124], addr_2281_7);

wire[31:0] addr_2282_7;

Selector_2 s2282_7(wires_570_6[2], addr_570_6, addr_positional[9131:9128], addr_2282_7);

wire[31:0] addr_2283_7;

Selector_2 s2283_7(wires_570_6[3], addr_570_6, addr_positional[9135:9132], addr_2283_7);

wire[31:0] addr_2284_7;

Selector_2 s2284_7(wires_571_6[0], addr_571_6, addr_positional[9139:9136], addr_2284_7);

wire[31:0] addr_2285_7;

Selector_2 s2285_7(wires_571_6[1], addr_571_6, addr_positional[9143:9140], addr_2285_7);

wire[31:0] addr_2286_7;

Selector_2 s2286_7(wires_571_6[2], addr_571_6, addr_positional[9147:9144], addr_2286_7);

wire[31:0] addr_2287_7;

Selector_2 s2287_7(wires_571_6[3], addr_571_6, addr_positional[9151:9148], addr_2287_7);

wire[31:0] addr_2288_7;

Selector_2 s2288_7(wires_572_6[0], addr_572_6, addr_positional[9155:9152], addr_2288_7);

wire[31:0] addr_2289_7;

Selector_2 s2289_7(wires_572_6[1], addr_572_6, addr_positional[9159:9156], addr_2289_7);

wire[31:0] addr_2290_7;

Selector_2 s2290_7(wires_572_6[2], addr_572_6, addr_positional[9163:9160], addr_2290_7);

wire[31:0] addr_2291_7;

Selector_2 s2291_7(wires_572_6[3], addr_572_6, addr_positional[9167:9164], addr_2291_7);

wire[31:0] addr_2292_7;

Selector_2 s2292_7(wires_573_6[0], addr_573_6, addr_positional[9171:9168], addr_2292_7);

wire[31:0] addr_2293_7;

Selector_2 s2293_7(wires_573_6[1], addr_573_6, addr_positional[9175:9172], addr_2293_7);

wire[31:0] addr_2294_7;

Selector_2 s2294_7(wires_573_6[2], addr_573_6, addr_positional[9179:9176], addr_2294_7);

wire[31:0] addr_2295_7;

Selector_2 s2295_7(wires_573_6[3], addr_573_6, addr_positional[9183:9180], addr_2295_7);

wire[31:0] addr_2296_7;

Selector_2 s2296_7(wires_574_6[0], addr_574_6, addr_positional[9187:9184], addr_2296_7);

wire[31:0] addr_2297_7;

Selector_2 s2297_7(wires_574_6[1], addr_574_6, addr_positional[9191:9188], addr_2297_7);

wire[31:0] addr_2298_7;

Selector_2 s2298_7(wires_574_6[2], addr_574_6, addr_positional[9195:9192], addr_2298_7);

wire[31:0] addr_2299_7;

Selector_2 s2299_7(wires_574_6[3], addr_574_6, addr_positional[9199:9196], addr_2299_7);

wire[31:0] addr_2300_7;

Selector_2 s2300_7(wires_575_6[0], addr_575_6, addr_positional[9203:9200], addr_2300_7);

wire[31:0] addr_2301_7;

Selector_2 s2301_7(wires_575_6[1], addr_575_6, addr_positional[9207:9204], addr_2301_7);

wire[31:0] addr_2302_7;

Selector_2 s2302_7(wires_575_6[2], addr_575_6, addr_positional[9211:9208], addr_2302_7);

wire[31:0] addr_2303_7;

Selector_2 s2303_7(wires_575_6[3], addr_575_6, addr_positional[9215:9212], addr_2303_7);

wire[31:0] addr_2304_7;

Selector_2 s2304_7(wires_576_6[0], addr_576_6, addr_positional[9219:9216], addr_2304_7);

wire[31:0] addr_2305_7;

Selector_2 s2305_7(wires_576_6[1], addr_576_6, addr_positional[9223:9220], addr_2305_7);

wire[31:0] addr_2306_7;

Selector_2 s2306_7(wires_576_6[2], addr_576_6, addr_positional[9227:9224], addr_2306_7);

wire[31:0] addr_2307_7;

Selector_2 s2307_7(wires_576_6[3], addr_576_6, addr_positional[9231:9228], addr_2307_7);

wire[31:0] addr_2308_7;

Selector_2 s2308_7(wires_577_6[0], addr_577_6, addr_positional[9235:9232], addr_2308_7);

wire[31:0] addr_2309_7;

Selector_2 s2309_7(wires_577_6[1], addr_577_6, addr_positional[9239:9236], addr_2309_7);

wire[31:0] addr_2310_7;

Selector_2 s2310_7(wires_577_6[2], addr_577_6, addr_positional[9243:9240], addr_2310_7);

wire[31:0] addr_2311_7;

Selector_2 s2311_7(wires_577_6[3], addr_577_6, addr_positional[9247:9244], addr_2311_7);

wire[31:0] addr_2312_7;

Selector_2 s2312_7(wires_578_6[0], addr_578_6, addr_positional[9251:9248], addr_2312_7);

wire[31:0] addr_2313_7;

Selector_2 s2313_7(wires_578_6[1], addr_578_6, addr_positional[9255:9252], addr_2313_7);

wire[31:0] addr_2314_7;

Selector_2 s2314_7(wires_578_6[2], addr_578_6, addr_positional[9259:9256], addr_2314_7);

wire[31:0] addr_2315_7;

Selector_2 s2315_7(wires_578_6[3], addr_578_6, addr_positional[9263:9260], addr_2315_7);

wire[31:0] addr_2316_7;

Selector_2 s2316_7(wires_579_6[0], addr_579_6, addr_positional[9267:9264], addr_2316_7);

wire[31:0] addr_2317_7;

Selector_2 s2317_7(wires_579_6[1], addr_579_6, addr_positional[9271:9268], addr_2317_7);

wire[31:0] addr_2318_7;

Selector_2 s2318_7(wires_579_6[2], addr_579_6, addr_positional[9275:9272], addr_2318_7);

wire[31:0] addr_2319_7;

Selector_2 s2319_7(wires_579_6[3], addr_579_6, addr_positional[9279:9276], addr_2319_7);

wire[31:0] addr_2320_7;

Selector_2 s2320_7(wires_580_6[0], addr_580_6, addr_positional[9283:9280], addr_2320_7);

wire[31:0] addr_2321_7;

Selector_2 s2321_7(wires_580_6[1], addr_580_6, addr_positional[9287:9284], addr_2321_7);

wire[31:0] addr_2322_7;

Selector_2 s2322_7(wires_580_6[2], addr_580_6, addr_positional[9291:9288], addr_2322_7);

wire[31:0] addr_2323_7;

Selector_2 s2323_7(wires_580_6[3], addr_580_6, addr_positional[9295:9292], addr_2323_7);

wire[31:0] addr_2324_7;

Selector_2 s2324_7(wires_581_6[0], addr_581_6, addr_positional[9299:9296], addr_2324_7);

wire[31:0] addr_2325_7;

Selector_2 s2325_7(wires_581_6[1], addr_581_6, addr_positional[9303:9300], addr_2325_7);

wire[31:0] addr_2326_7;

Selector_2 s2326_7(wires_581_6[2], addr_581_6, addr_positional[9307:9304], addr_2326_7);

wire[31:0] addr_2327_7;

Selector_2 s2327_7(wires_581_6[3], addr_581_6, addr_positional[9311:9308], addr_2327_7);

wire[31:0] addr_2328_7;

Selector_2 s2328_7(wires_582_6[0], addr_582_6, addr_positional[9315:9312], addr_2328_7);

wire[31:0] addr_2329_7;

Selector_2 s2329_7(wires_582_6[1], addr_582_6, addr_positional[9319:9316], addr_2329_7);

wire[31:0] addr_2330_7;

Selector_2 s2330_7(wires_582_6[2], addr_582_6, addr_positional[9323:9320], addr_2330_7);

wire[31:0] addr_2331_7;

Selector_2 s2331_7(wires_582_6[3], addr_582_6, addr_positional[9327:9324], addr_2331_7);

wire[31:0] addr_2332_7;

Selector_2 s2332_7(wires_583_6[0], addr_583_6, addr_positional[9331:9328], addr_2332_7);

wire[31:0] addr_2333_7;

Selector_2 s2333_7(wires_583_6[1], addr_583_6, addr_positional[9335:9332], addr_2333_7);

wire[31:0] addr_2334_7;

Selector_2 s2334_7(wires_583_6[2], addr_583_6, addr_positional[9339:9336], addr_2334_7);

wire[31:0] addr_2335_7;

Selector_2 s2335_7(wires_583_6[3], addr_583_6, addr_positional[9343:9340], addr_2335_7);

wire[31:0] addr_2336_7;

Selector_2 s2336_7(wires_584_6[0], addr_584_6, addr_positional[9347:9344], addr_2336_7);

wire[31:0] addr_2337_7;

Selector_2 s2337_7(wires_584_6[1], addr_584_6, addr_positional[9351:9348], addr_2337_7);

wire[31:0] addr_2338_7;

Selector_2 s2338_7(wires_584_6[2], addr_584_6, addr_positional[9355:9352], addr_2338_7);

wire[31:0] addr_2339_7;

Selector_2 s2339_7(wires_584_6[3], addr_584_6, addr_positional[9359:9356], addr_2339_7);

wire[31:0] addr_2340_7;

Selector_2 s2340_7(wires_585_6[0], addr_585_6, addr_positional[9363:9360], addr_2340_7);

wire[31:0] addr_2341_7;

Selector_2 s2341_7(wires_585_6[1], addr_585_6, addr_positional[9367:9364], addr_2341_7);

wire[31:0] addr_2342_7;

Selector_2 s2342_7(wires_585_6[2], addr_585_6, addr_positional[9371:9368], addr_2342_7);

wire[31:0] addr_2343_7;

Selector_2 s2343_7(wires_585_6[3], addr_585_6, addr_positional[9375:9372], addr_2343_7);

wire[31:0] addr_2344_7;

Selector_2 s2344_7(wires_586_6[0], addr_586_6, addr_positional[9379:9376], addr_2344_7);

wire[31:0] addr_2345_7;

Selector_2 s2345_7(wires_586_6[1], addr_586_6, addr_positional[9383:9380], addr_2345_7);

wire[31:0] addr_2346_7;

Selector_2 s2346_7(wires_586_6[2], addr_586_6, addr_positional[9387:9384], addr_2346_7);

wire[31:0] addr_2347_7;

Selector_2 s2347_7(wires_586_6[3], addr_586_6, addr_positional[9391:9388], addr_2347_7);

wire[31:0] addr_2348_7;

Selector_2 s2348_7(wires_587_6[0], addr_587_6, addr_positional[9395:9392], addr_2348_7);

wire[31:0] addr_2349_7;

Selector_2 s2349_7(wires_587_6[1], addr_587_6, addr_positional[9399:9396], addr_2349_7);

wire[31:0] addr_2350_7;

Selector_2 s2350_7(wires_587_6[2], addr_587_6, addr_positional[9403:9400], addr_2350_7);

wire[31:0] addr_2351_7;

Selector_2 s2351_7(wires_587_6[3], addr_587_6, addr_positional[9407:9404], addr_2351_7);

wire[31:0] addr_2352_7;

Selector_2 s2352_7(wires_588_6[0], addr_588_6, addr_positional[9411:9408], addr_2352_7);

wire[31:0] addr_2353_7;

Selector_2 s2353_7(wires_588_6[1], addr_588_6, addr_positional[9415:9412], addr_2353_7);

wire[31:0] addr_2354_7;

Selector_2 s2354_7(wires_588_6[2], addr_588_6, addr_positional[9419:9416], addr_2354_7);

wire[31:0] addr_2355_7;

Selector_2 s2355_7(wires_588_6[3], addr_588_6, addr_positional[9423:9420], addr_2355_7);

wire[31:0] addr_2356_7;

Selector_2 s2356_7(wires_589_6[0], addr_589_6, addr_positional[9427:9424], addr_2356_7);

wire[31:0] addr_2357_7;

Selector_2 s2357_7(wires_589_6[1], addr_589_6, addr_positional[9431:9428], addr_2357_7);

wire[31:0] addr_2358_7;

Selector_2 s2358_7(wires_589_6[2], addr_589_6, addr_positional[9435:9432], addr_2358_7);

wire[31:0] addr_2359_7;

Selector_2 s2359_7(wires_589_6[3], addr_589_6, addr_positional[9439:9436], addr_2359_7);

wire[31:0] addr_2360_7;

Selector_2 s2360_7(wires_590_6[0], addr_590_6, addr_positional[9443:9440], addr_2360_7);

wire[31:0] addr_2361_7;

Selector_2 s2361_7(wires_590_6[1], addr_590_6, addr_positional[9447:9444], addr_2361_7);

wire[31:0] addr_2362_7;

Selector_2 s2362_7(wires_590_6[2], addr_590_6, addr_positional[9451:9448], addr_2362_7);

wire[31:0] addr_2363_7;

Selector_2 s2363_7(wires_590_6[3], addr_590_6, addr_positional[9455:9452], addr_2363_7);

wire[31:0] addr_2364_7;

Selector_2 s2364_7(wires_591_6[0], addr_591_6, addr_positional[9459:9456], addr_2364_7);

wire[31:0] addr_2365_7;

Selector_2 s2365_7(wires_591_6[1], addr_591_6, addr_positional[9463:9460], addr_2365_7);

wire[31:0] addr_2366_7;

Selector_2 s2366_7(wires_591_6[2], addr_591_6, addr_positional[9467:9464], addr_2366_7);

wire[31:0] addr_2367_7;

Selector_2 s2367_7(wires_591_6[3], addr_591_6, addr_positional[9471:9468], addr_2367_7);

wire[31:0] addr_2368_7;

Selector_2 s2368_7(wires_592_6[0], addr_592_6, addr_positional[9475:9472], addr_2368_7);

wire[31:0] addr_2369_7;

Selector_2 s2369_7(wires_592_6[1], addr_592_6, addr_positional[9479:9476], addr_2369_7);

wire[31:0] addr_2370_7;

Selector_2 s2370_7(wires_592_6[2], addr_592_6, addr_positional[9483:9480], addr_2370_7);

wire[31:0] addr_2371_7;

Selector_2 s2371_7(wires_592_6[3], addr_592_6, addr_positional[9487:9484], addr_2371_7);

wire[31:0] addr_2372_7;

Selector_2 s2372_7(wires_593_6[0], addr_593_6, addr_positional[9491:9488], addr_2372_7);

wire[31:0] addr_2373_7;

Selector_2 s2373_7(wires_593_6[1], addr_593_6, addr_positional[9495:9492], addr_2373_7);

wire[31:0] addr_2374_7;

Selector_2 s2374_7(wires_593_6[2], addr_593_6, addr_positional[9499:9496], addr_2374_7);

wire[31:0] addr_2375_7;

Selector_2 s2375_7(wires_593_6[3], addr_593_6, addr_positional[9503:9500], addr_2375_7);

wire[31:0] addr_2376_7;

Selector_2 s2376_7(wires_594_6[0], addr_594_6, addr_positional[9507:9504], addr_2376_7);

wire[31:0] addr_2377_7;

Selector_2 s2377_7(wires_594_6[1], addr_594_6, addr_positional[9511:9508], addr_2377_7);

wire[31:0] addr_2378_7;

Selector_2 s2378_7(wires_594_6[2], addr_594_6, addr_positional[9515:9512], addr_2378_7);

wire[31:0] addr_2379_7;

Selector_2 s2379_7(wires_594_6[3], addr_594_6, addr_positional[9519:9516], addr_2379_7);

wire[31:0] addr_2380_7;

Selector_2 s2380_7(wires_595_6[0], addr_595_6, addr_positional[9523:9520], addr_2380_7);

wire[31:0] addr_2381_7;

Selector_2 s2381_7(wires_595_6[1], addr_595_6, addr_positional[9527:9524], addr_2381_7);

wire[31:0] addr_2382_7;

Selector_2 s2382_7(wires_595_6[2], addr_595_6, addr_positional[9531:9528], addr_2382_7);

wire[31:0] addr_2383_7;

Selector_2 s2383_7(wires_595_6[3], addr_595_6, addr_positional[9535:9532], addr_2383_7);

wire[31:0] addr_2384_7;

Selector_2 s2384_7(wires_596_6[0], addr_596_6, addr_positional[9539:9536], addr_2384_7);

wire[31:0] addr_2385_7;

Selector_2 s2385_7(wires_596_6[1], addr_596_6, addr_positional[9543:9540], addr_2385_7);

wire[31:0] addr_2386_7;

Selector_2 s2386_7(wires_596_6[2], addr_596_6, addr_positional[9547:9544], addr_2386_7);

wire[31:0] addr_2387_7;

Selector_2 s2387_7(wires_596_6[3], addr_596_6, addr_positional[9551:9548], addr_2387_7);

wire[31:0] addr_2388_7;

Selector_2 s2388_7(wires_597_6[0], addr_597_6, addr_positional[9555:9552], addr_2388_7);

wire[31:0] addr_2389_7;

Selector_2 s2389_7(wires_597_6[1], addr_597_6, addr_positional[9559:9556], addr_2389_7);

wire[31:0] addr_2390_7;

Selector_2 s2390_7(wires_597_6[2], addr_597_6, addr_positional[9563:9560], addr_2390_7);

wire[31:0] addr_2391_7;

Selector_2 s2391_7(wires_597_6[3], addr_597_6, addr_positional[9567:9564], addr_2391_7);

wire[31:0] addr_2392_7;

Selector_2 s2392_7(wires_598_6[0], addr_598_6, addr_positional[9571:9568], addr_2392_7);

wire[31:0] addr_2393_7;

Selector_2 s2393_7(wires_598_6[1], addr_598_6, addr_positional[9575:9572], addr_2393_7);

wire[31:0] addr_2394_7;

Selector_2 s2394_7(wires_598_6[2], addr_598_6, addr_positional[9579:9576], addr_2394_7);

wire[31:0] addr_2395_7;

Selector_2 s2395_7(wires_598_6[3], addr_598_6, addr_positional[9583:9580], addr_2395_7);

wire[31:0] addr_2396_7;

Selector_2 s2396_7(wires_599_6[0], addr_599_6, addr_positional[9587:9584], addr_2396_7);

wire[31:0] addr_2397_7;

Selector_2 s2397_7(wires_599_6[1], addr_599_6, addr_positional[9591:9588], addr_2397_7);

wire[31:0] addr_2398_7;

Selector_2 s2398_7(wires_599_6[2], addr_599_6, addr_positional[9595:9592], addr_2398_7);

wire[31:0] addr_2399_7;

Selector_2 s2399_7(wires_599_6[3], addr_599_6, addr_positional[9599:9596], addr_2399_7);

wire[31:0] addr_2400_7;

Selector_2 s2400_7(wires_600_6[0], addr_600_6, addr_positional[9603:9600], addr_2400_7);

wire[31:0] addr_2401_7;

Selector_2 s2401_7(wires_600_6[1], addr_600_6, addr_positional[9607:9604], addr_2401_7);

wire[31:0] addr_2402_7;

Selector_2 s2402_7(wires_600_6[2], addr_600_6, addr_positional[9611:9608], addr_2402_7);

wire[31:0] addr_2403_7;

Selector_2 s2403_7(wires_600_6[3], addr_600_6, addr_positional[9615:9612], addr_2403_7);

wire[31:0] addr_2404_7;

Selector_2 s2404_7(wires_601_6[0], addr_601_6, addr_positional[9619:9616], addr_2404_7);

wire[31:0] addr_2405_7;

Selector_2 s2405_7(wires_601_6[1], addr_601_6, addr_positional[9623:9620], addr_2405_7);

wire[31:0] addr_2406_7;

Selector_2 s2406_7(wires_601_6[2], addr_601_6, addr_positional[9627:9624], addr_2406_7);

wire[31:0] addr_2407_7;

Selector_2 s2407_7(wires_601_6[3], addr_601_6, addr_positional[9631:9628], addr_2407_7);

wire[31:0] addr_2408_7;

Selector_2 s2408_7(wires_602_6[0], addr_602_6, addr_positional[9635:9632], addr_2408_7);

wire[31:0] addr_2409_7;

Selector_2 s2409_7(wires_602_6[1], addr_602_6, addr_positional[9639:9636], addr_2409_7);

wire[31:0] addr_2410_7;

Selector_2 s2410_7(wires_602_6[2], addr_602_6, addr_positional[9643:9640], addr_2410_7);

wire[31:0] addr_2411_7;

Selector_2 s2411_7(wires_602_6[3], addr_602_6, addr_positional[9647:9644], addr_2411_7);

wire[31:0] addr_2412_7;

Selector_2 s2412_7(wires_603_6[0], addr_603_6, addr_positional[9651:9648], addr_2412_7);

wire[31:0] addr_2413_7;

Selector_2 s2413_7(wires_603_6[1], addr_603_6, addr_positional[9655:9652], addr_2413_7);

wire[31:0] addr_2414_7;

Selector_2 s2414_7(wires_603_6[2], addr_603_6, addr_positional[9659:9656], addr_2414_7);

wire[31:0] addr_2415_7;

Selector_2 s2415_7(wires_603_6[3], addr_603_6, addr_positional[9663:9660], addr_2415_7);

wire[31:0] addr_2416_7;

Selector_2 s2416_7(wires_604_6[0], addr_604_6, addr_positional[9667:9664], addr_2416_7);

wire[31:0] addr_2417_7;

Selector_2 s2417_7(wires_604_6[1], addr_604_6, addr_positional[9671:9668], addr_2417_7);

wire[31:0] addr_2418_7;

Selector_2 s2418_7(wires_604_6[2], addr_604_6, addr_positional[9675:9672], addr_2418_7);

wire[31:0] addr_2419_7;

Selector_2 s2419_7(wires_604_6[3], addr_604_6, addr_positional[9679:9676], addr_2419_7);

wire[31:0] addr_2420_7;

Selector_2 s2420_7(wires_605_6[0], addr_605_6, addr_positional[9683:9680], addr_2420_7);

wire[31:0] addr_2421_7;

Selector_2 s2421_7(wires_605_6[1], addr_605_6, addr_positional[9687:9684], addr_2421_7);

wire[31:0] addr_2422_7;

Selector_2 s2422_7(wires_605_6[2], addr_605_6, addr_positional[9691:9688], addr_2422_7);

wire[31:0] addr_2423_7;

Selector_2 s2423_7(wires_605_6[3], addr_605_6, addr_positional[9695:9692], addr_2423_7);

wire[31:0] addr_2424_7;

Selector_2 s2424_7(wires_606_6[0], addr_606_6, addr_positional[9699:9696], addr_2424_7);

wire[31:0] addr_2425_7;

Selector_2 s2425_7(wires_606_6[1], addr_606_6, addr_positional[9703:9700], addr_2425_7);

wire[31:0] addr_2426_7;

Selector_2 s2426_7(wires_606_6[2], addr_606_6, addr_positional[9707:9704], addr_2426_7);

wire[31:0] addr_2427_7;

Selector_2 s2427_7(wires_606_6[3], addr_606_6, addr_positional[9711:9708], addr_2427_7);

wire[31:0] addr_2428_7;

Selector_2 s2428_7(wires_607_6[0], addr_607_6, addr_positional[9715:9712], addr_2428_7);

wire[31:0] addr_2429_7;

Selector_2 s2429_7(wires_607_6[1], addr_607_6, addr_positional[9719:9716], addr_2429_7);

wire[31:0] addr_2430_7;

Selector_2 s2430_7(wires_607_6[2], addr_607_6, addr_positional[9723:9720], addr_2430_7);

wire[31:0] addr_2431_7;

Selector_2 s2431_7(wires_607_6[3], addr_607_6, addr_positional[9727:9724], addr_2431_7);

wire[31:0] addr_2432_7;

Selector_2 s2432_7(wires_608_6[0], addr_608_6, addr_positional[9731:9728], addr_2432_7);

wire[31:0] addr_2433_7;

Selector_2 s2433_7(wires_608_6[1], addr_608_6, addr_positional[9735:9732], addr_2433_7);

wire[31:0] addr_2434_7;

Selector_2 s2434_7(wires_608_6[2], addr_608_6, addr_positional[9739:9736], addr_2434_7);

wire[31:0] addr_2435_7;

Selector_2 s2435_7(wires_608_6[3], addr_608_6, addr_positional[9743:9740], addr_2435_7);

wire[31:0] addr_2436_7;

Selector_2 s2436_7(wires_609_6[0], addr_609_6, addr_positional[9747:9744], addr_2436_7);

wire[31:0] addr_2437_7;

Selector_2 s2437_7(wires_609_6[1], addr_609_6, addr_positional[9751:9748], addr_2437_7);

wire[31:0] addr_2438_7;

Selector_2 s2438_7(wires_609_6[2], addr_609_6, addr_positional[9755:9752], addr_2438_7);

wire[31:0] addr_2439_7;

Selector_2 s2439_7(wires_609_6[3], addr_609_6, addr_positional[9759:9756], addr_2439_7);

wire[31:0] addr_2440_7;

Selector_2 s2440_7(wires_610_6[0], addr_610_6, addr_positional[9763:9760], addr_2440_7);

wire[31:0] addr_2441_7;

Selector_2 s2441_7(wires_610_6[1], addr_610_6, addr_positional[9767:9764], addr_2441_7);

wire[31:0] addr_2442_7;

Selector_2 s2442_7(wires_610_6[2], addr_610_6, addr_positional[9771:9768], addr_2442_7);

wire[31:0] addr_2443_7;

Selector_2 s2443_7(wires_610_6[3], addr_610_6, addr_positional[9775:9772], addr_2443_7);

wire[31:0] addr_2444_7;

Selector_2 s2444_7(wires_611_6[0], addr_611_6, addr_positional[9779:9776], addr_2444_7);

wire[31:0] addr_2445_7;

Selector_2 s2445_7(wires_611_6[1], addr_611_6, addr_positional[9783:9780], addr_2445_7);

wire[31:0] addr_2446_7;

Selector_2 s2446_7(wires_611_6[2], addr_611_6, addr_positional[9787:9784], addr_2446_7);

wire[31:0] addr_2447_7;

Selector_2 s2447_7(wires_611_6[3], addr_611_6, addr_positional[9791:9788], addr_2447_7);

wire[31:0] addr_2448_7;

Selector_2 s2448_7(wires_612_6[0], addr_612_6, addr_positional[9795:9792], addr_2448_7);

wire[31:0] addr_2449_7;

Selector_2 s2449_7(wires_612_6[1], addr_612_6, addr_positional[9799:9796], addr_2449_7);

wire[31:0] addr_2450_7;

Selector_2 s2450_7(wires_612_6[2], addr_612_6, addr_positional[9803:9800], addr_2450_7);

wire[31:0] addr_2451_7;

Selector_2 s2451_7(wires_612_6[3], addr_612_6, addr_positional[9807:9804], addr_2451_7);

wire[31:0] addr_2452_7;

Selector_2 s2452_7(wires_613_6[0], addr_613_6, addr_positional[9811:9808], addr_2452_7);

wire[31:0] addr_2453_7;

Selector_2 s2453_7(wires_613_6[1], addr_613_6, addr_positional[9815:9812], addr_2453_7);

wire[31:0] addr_2454_7;

Selector_2 s2454_7(wires_613_6[2], addr_613_6, addr_positional[9819:9816], addr_2454_7);

wire[31:0] addr_2455_7;

Selector_2 s2455_7(wires_613_6[3], addr_613_6, addr_positional[9823:9820], addr_2455_7);

wire[31:0] addr_2456_7;

Selector_2 s2456_7(wires_614_6[0], addr_614_6, addr_positional[9827:9824], addr_2456_7);

wire[31:0] addr_2457_7;

Selector_2 s2457_7(wires_614_6[1], addr_614_6, addr_positional[9831:9828], addr_2457_7);

wire[31:0] addr_2458_7;

Selector_2 s2458_7(wires_614_6[2], addr_614_6, addr_positional[9835:9832], addr_2458_7);

wire[31:0] addr_2459_7;

Selector_2 s2459_7(wires_614_6[3], addr_614_6, addr_positional[9839:9836], addr_2459_7);

wire[31:0] addr_2460_7;

Selector_2 s2460_7(wires_615_6[0], addr_615_6, addr_positional[9843:9840], addr_2460_7);

wire[31:0] addr_2461_7;

Selector_2 s2461_7(wires_615_6[1], addr_615_6, addr_positional[9847:9844], addr_2461_7);

wire[31:0] addr_2462_7;

Selector_2 s2462_7(wires_615_6[2], addr_615_6, addr_positional[9851:9848], addr_2462_7);

wire[31:0] addr_2463_7;

Selector_2 s2463_7(wires_615_6[3], addr_615_6, addr_positional[9855:9852], addr_2463_7);

wire[31:0] addr_2464_7;

Selector_2 s2464_7(wires_616_6[0], addr_616_6, addr_positional[9859:9856], addr_2464_7);

wire[31:0] addr_2465_7;

Selector_2 s2465_7(wires_616_6[1], addr_616_6, addr_positional[9863:9860], addr_2465_7);

wire[31:0] addr_2466_7;

Selector_2 s2466_7(wires_616_6[2], addr_616_6, addr_positional[9867:9864], addr_2466_7);

wire[31:0] addr_2467_7;

Selector_2 s2467_7(wires_616_6[3], addr_616_6, addr_positional[9871:9868], addr_2467_7);

wire[31:0] addr_2468_7;

Selector_2 s2468_7(wires_617_6[0], addr_617_6, addr_positional[9875:9872], addr_2468_7);

wire[31:0] addr_2469_7;

Selector_2 s2469_7(wires_617_6[1], addr_617_6, addr_positional[9879:9876], addr_2469_7);

wire[31:0] addr_2470_7;

Selector_2 s2470_7(wires_617_6[2], addr_617_6, addr_positional[9883:9880], addr_2470_7);

wire[31:0] addr_2471_7;

Selector_2 s2471_7(wires_617_6[3], addr_617_6, addr_positional[9887:9884], addr_2471_7);

wire[31:0] addr_2472_7;

Selector_2 s2472_7(wires_618_6[0], addr_618_6, addr_positional[9891:9888], addr_2472_7);

wire[31:0] addr_2473_7;

Selector_2 s2473_7(wires_618_6[1], addr_618_6, addr_positional[9895:9892], addr_2473_7);

wire[31:0] addr_2474_7;

Selector_2 s2474_7(wires_618_6[2], addr_618_6, addr_positional[9899:9896], addr_2474_7);

wire[31:0] addr_2475_7;

Selector_2 s2475_7(wires_618_6[3], addr_618_6, addr_positional[9903:9900], addr_2475_7);

wire[31:0] addr_2476_7;

Selector_2 s2476_7(wires_619_6[0], addr_619_6, addr_positional[9907:9904], addr_2476_7);

wire[31:0] addr_2477_7;

Selector_2 s2477_7(wires_619_6[1], addr_619_6, addr_positional[9911:9908], addr_2477_7);

wire[31:0] addr_2478_7;

Selector_2 s2478_7(wires_619_6[2], addr_619_6, addr_positional[9915:9912], addr_2478_7);

wire[31:0] addr_2479_7;

Selector_2 s2479_7(wires_619_6[3], addr_619_6, addr_positional[9919:9916], addr_2479_7);

wire[31:0] addr_2480_7;

Selector_2 s2480_7(wires_620_6[0], addr_620_6, addr_positional[9923:9920], addr_2480_7);

wire[31:0] addr_2481_7;

Selector_2 s2481_7(wires_620_6[1], addr_620_6, addr_positional[9927:9924], addr_2481_7);

wire[31:0] addr_2482_7;

Selector_2 s2482_7(wires_620_6[2], addr_620_6, addr_positional[9931:9928], addr_2482_7);

wire[31:0] addr_2483_7;

Selector_2 s2483_7(wires_620_6[3], addr_620_6, addr_positional[9935:9932], addr_2483_7);

wire[31:0] addr_2484_7;

Selector_2 s2484_7(wires_621_6[0], addr_621_6, addr_positional[9939:9936], addr_2484_7);

wire[31:0] addr_2485_7;

Selector_2 s2485_7(wires_621_6[1], addr_621_6, addr_positional[9943:9940], addr_2485_7);

wire[31:0] addr_2486_7;

Selector_2 s2486_7(wires_621_6[2], addr_621_6, addr_positional[9947:9944], addr_2486_7);

wire[31:0] addr_2487_7;

Selector_2 s2487_7(wires_621_6[3], addr_621_6, addr_positional[9951:9948], addr_2487_7);

wire[31:0] addr_2488_7;

Selector_2 s2488_7(wires_622_6[0], addr_622_6, addr_positional[9955:9952], addr_2488_7);

wire[31:0] addr_2489_7;

Selector_2 s2489_7(wires_622_6[1], addr_622_6, addr_positional[9959:9956], addr_2489_7);

wire[31:0] addr_2490_7;

Selector_2 s2490_7(wires_622_6[2], addr_622_6, addr_positional[9963:9960], addr_2490_7);

wire[31:0] addr_2491_7;

Selector_2 s2491_7(wires_622_6[3], addr_622_6, addr_positional[9967:9964], addr_2491_7);

wire[31:0] addr_2492_7;

Selector_2 s2492_7(wires_623_6[0], addr_623_6, addr_positional[9971:9968], addr_2492_7);

wire[31:0] addr_2493_7;

Selector_2 s2493_7(wires_623_6[1], addr_623_6, addr_positional[9975:9972], addr_2493_7);

wire[31:0] addr_2494_7;

Selector_2 s2494_7(wires_623_6[2], addr_623_6, addr_positional[9979:9976], addr_2494_7);

wire[31:0] addr_2495_7;

Selector_2 s2495_7(wires_623_6[3], addr_623_6, addr_positional[9983:9980], addr_2495_7);

wire[31:0] addr_2496_7;

Selector_2 s2496_7(wires_624_6[0], addr_624_6, addr_positional[9987:9984], addr_2496_7);

wire[31:0] addr_2497_7;

Selector_2 s2497_7(wires_624_6[1], addr_624_6, addr_positional[9991:9988], addr_2497_7);

wire[31:0] addr_2498_7;

Selector_2 s2498_7(wires_624_6[2], addr_624_6, addr_positional[9995:9992], addr_2498_7);

wire[31:0] addr_2499_7;

Selector_2 s2499_7(wires_624_6[3], addr_624_6, addr_positional[9999:9996], addr_2499_7);

wire[31:0] addr_2500_7;

Selector_2 s2500_7(wires_625_6[0], addr_625_6, addr_positional[10003:10000], addr_2500_7);

wire[31:0] addr_2501_7;

Selector_2 s2501_7(wires_625_6[1], addr_625_6, addr_positional[10007:10004], addr_2501_7);

wire[31:0] addr_2502_7;

Selector_2 s2502_7(wires_625_6[2], addr_625_6, addr_positional[10011:10008], addr_2502_7);

wire[31:0] addr_2503_7;

Selector_2 s2503_7(wires_625_6[3], addr_625_6, addr_positional[10015:10012], addr_2503_7);

wire[31:0] addr_2504_7;

Selector_2 s2504_7(wires_626_6[0], addr_626_6, addr_positional[10019:10016], addr_2504_7);

wire[31:0] addr_2505_7;

Selector_2 s2505_7(wires_626_6[1], addr_626_6, addr_positional[10023:10020], addr_2505_7);

wire[31:0] addr_2506_7;

Selector_2 s2506_7(wires_626_6[2], addr_626_6, addr_positional[10027:10024], addr_2506_7);

wire[31:0] addr_2507_7;

Selector_2 s2507_7(wires_626_6[3], addr_626_6, addr_positional[10031:10028], addr_2507_7);

wire[31:0] addr_2508_7;

Selector_2 s2508_7(wires_627_6[0], addr_627_6, addr_positional[10035:10032], addr_2508_7);

wire[31:0] addr_2509_7;

Selector_2 s2509_7(wires_627_6[1], addr_627_6, addr_positional[10039:10036], addr_2509_7);

wire[31:0] addr_2510_7;

Selector_2 s2510_7(wires_627_6[2], addr_627_6, addr_positional[10043:10040], addr_2510_7);

wire[31:0] addr_2511_7;

Selector_2 s2511_7(wires_627_6[3], addr_627_6, addr_positional[10047:10044], addr_2511_7);

wire[31:0] addr_2512_7;

Selector_2 s2512_7(wires_628_6[0], addr_628_6, addr_positional[10051:10048], addr_2512_7);

wire[31:0] addr_2513_7;

Selector_2 s2513_7(wires_628_6[1], addr_628_6, addr_positional[10055:10052], addr_2513_7);

wire[31:0] addr_2514_7;

Selector_2 s2514_7(wires_628_6[2], addr_628_6, addr_positional[10059:10056], addr_2514_7);

wire[31:0] addr_2515_7;

Selector_2 s2515_7(wires_628_6[3], addr_628_6, addr_positional[10063:10060], addr_2515_7);

wire[31:0] addr_2516_7;

Selector_2 s2516_7(wires_629_6[0], addr_629_6, addr_positional[10067:10064], addr_2516_7);

wire[31:0] addr_2517_7;

Selector_2 s2517_7(wires_629_6[1], addr_629_6, addr_positional[10071:10068], addr_2517_7);

wire[31:0] addr_2518_7;

Selector_2 s2518_7(wires_629_6[2], addr_629_6, addr_positional[10075:10072], addr_2518_7);

wire[31:0] addr_2519_7;

Selector_2 s2519_7(wires_629_6[3], addr_629_6, addr_positional[10079:10076], addr_2519_7);

wire[31:0] addr_2520_7;

Selector_2 s2520_7(wires_630_6[0], addr_630_6, addr_positional[10083:10080], addr_2520_7);

wire[31:0] addr_2521_7;

Selector_2 s2521_7(wires_630_6[1], addr_630_6, addr_positional[10087:10084], addr_2521_7);

wire[31:0] addr_2522_7;

Selector_2 s2522_7(wires_630_6[2], addr_630_6, addr_positional[10091:10088], addr_2522_7);

wire[31:0] addr_2523_7;

Selector_2 s2523_7(wires_630_6[3], addr_630_6, addr_positional[10095:10092], addr_2523_7);

wire[31:0] addr_2524_7;

Selector_2 s2524_7(wires_631_6[0], addr_631_6, addr_positional[10099:10096], addr_2524_7);

wire[31:0] addr_2525_7;

Selector_2 s2525_7(wires_631_6[1], addr_631_6, addr_positional[10103:10100], addr_2525_7);

wire[31:0] addr_2526_7;

Selector_2 s2526_7(wires_631_6[2], addr_631_6, addr_positional[10107:10104], addr_2526_7);

wire[31:0] addr_2527_7;

Selector_2 s2527_7(wires_631_6[3], addr_631_6, addr_positional[10111:10108], addr_2527_7);

wire[31:0] addr_2528_7;

Selector_2 s2528_7(wires_632_6[0], addr_632_6, addr_positional[10115:10112], addr_2528_7);

wire[31:0] addr_2529_7;

Selector_2 s2529_7(wires_632_6[1], addr_632_6, addr_positional[10119:10116], addr_2529_7);

wire[31:0] addr_2530_7;

Selector_2 s2530_7(wires_632_6[2], addr_632_6, addr_positional[10123:10120], addr_2530_7);

wire[31:0] addr_2531_7;

Selector_2 s2531_7(wires_632_6[3], addr_632_6, addr_positional[10127:10124], addr_2531_7);

wire[31:0] addr_2532_7;

Selector_2 s2532_7(wires_633_6[0], addr_633_6, addr_positional[10131:10128], addr_2532_7);

wire[31:0] addr_2533_7;

Selector_2 s2533_7(wires_633_6[1], addr_633_6, addr_positional[10135:10132], addr_2533_7);

wire[31:0] addr_2534_7;

Selector_2 s2534_7(wires_633_6[2], addr_633_6, addr_positional[10139:10136], addr_2534_7);

wire[31:0] addr_2535_7;

Selector_2 s2535_7(wires_633_6[3], addr_633_6, addr_positional[10143:10140], addr_2535_7);

wire[31:0] addr_2536_7;

Selector_2 s2536_7(wires_634_6[0], addr_634_6, addr_positional[10147:10144], addr_2536_7);

wire[31:0] addr_2537_7;

Selector_2 s2537_7(wires_634_6[1], addr_634_6, addr_positional[10151:10148], addr_2537_7);

wire[31:0] addr_2538_7;

Selector_2 s2538_7(wires_634_6[2], addr_634_6, addr_positional[10155:10152], addr_2538_7);

wire[31:0] addr_2539_7;

Selector_2 s2539_7(wires_634_6[3], addr_634_6, addr_positional[10159:10156], addr_2539_7);

wire[31:0] addr_2540_7;

Selector_2 s2540_7(wires_635_6[0], addr_635_6, addr_positional[10163:10160], addr_2540_7);

wire[31:0] addr_2541_7;

Selector_2 s2541_7(wires_635_6[1], addr_635_6, addr_positional[10167:10164], addr_2541_7);

wire[31:0] addr_2542_7;

Selector_2 s2542_7(wires_635_6[2], addr_635_6, addr_positional[10171:10168], addr_2542_7);

wire[31:0] addr_2543_7;

Selector_2 s2543_7(wires_635_6[3], addr_635_6, addr_positional[10175:10172], addr_2543_7);

wire[31:0] addr_2544_7;

Selector_2 s2544_7(wires_636_6[0], addr_636_6, addr_positional[10179:10176], addr_2544_7);

wire[31:0] addr_2545_7;

Selector_2 s2545_7(wires_636_6[1], addr_636_6, addr_positional[10183:10180], addr_2545_7);

wire[31:0] addr_2546_7;

Selector_2 s2546_7(wires_636_6[2], addr_636_6, addr_positional[10187:10184], addr_2546_7);

wire[31:0] addr_2547_7;

Selector_2 s2547_7(wires_636_6[3], addr_636_6, addr_positional[10191:10188], addr_2547_7);

wire[31:0] addr_2548_7;

Selector_2 s2548_7(wires_637_6[0], addr_637_6, addr_positional[10195:10192], addr_2548_7);

wire[31:0] addr_2549_7;

Selector_2 s2549_7(wires_637_6[1], addr_637_6, addr_positional[10199:10196], addr_2549_7);

wire[31:0] addr_2550_7;

Selector_2 s2550_7(wires_637_6[2], addr_637_6, addr_positional[10203:10200], addr_2550_7);

wire[31:0] addr_2551_7;

Selector_2 s2551_7(wires_637_6[3], addr_637_6, addr_positional[10207:10204], addr_2551_7);

wire[31:0] addr_2552_7;

Selector_2 s2552_7(wires_638_6[0], addr_638_6, addr_positional[10211:10208], addr_2552_7);

wire[31:0] addr_2553_7;

Selector_2 s2553_7(wires_638_6[1], addr_638_6, addr_positional[10215:10212], addr_2553_7);

wire[31:0] addr_2554_7;

Selector_2 s2554_7(wires_638_6[2], addr_638_6, addr_positional[10219:10216], addr_2554_7);

wire[31:0] addr_2555_7;

Selector_2 s2555_7(wires_638_6[3], addr_638_6, addr_positional[10223:10220], addr_2555_7);

wire[31:0] addr_2556_7;

Selector_2 s2556_7(wires_639_6[0], addr_639_6, addr_positional[10227:10224], addr_2556_7);

wire[31:0] addr_2557_7;

Selector_2 s2557_7(wires_639_6[1], addr_639_6, addr_positional[10231:10228], addr_2557_7);

wire[31:0] addr_2558_7;

Selector_2 s2558_7(wires_639_6[2], addr_639_6, addr_positional[10235:10232], addr_2558_7);

wire[31:0] addr_2559_7;

Selector_2 s2559_7(wires_639_6[3], addr_639_6, addr_positional[10239:10236], addr_2559_7);

wire[31:0] addr_2560_7;

Selector_2 s2560_7(wires_640_6[0], addr_640_6, addr_positional[10243:10240], addr_2560_7);

wire[31:0] addr_2561_7;

Selector_2 s2561_7(wires_640_6[1], addr_640_6, addr_positional[10247:10244], addr_2561_7);

wire[31:0] addr_2562_7;

Selector_2 s2562_7(wires_640_6[2], addr_640_6, addr_positional[10251:10248], addr_2562_7);

wire[31:0] addr_2563_7;

Selector_2 s2563_7(wires_640_6[3], addr_640_6, addr_positional[10255:10252], addr_2563_7);

wire[31:0] addr_2564_7;

Selector_2 s2564_7(wires_641_6[0], addr_641_6, addr_positional[10259:10256], addr_2564_7);

wire[31:0] addr_2565_7;

Selector_2 s2565_7(wires_641_6[1], addr_641_6, addr_positional[10263:10260], addr_2565_7);

wire[31:0] addr_2566_7;

Selector_2 s2566_7(wires_641_6[2], addr_641_6, addr_positional[10267:10264], addr_2566_7);

wire[31:0] addr_2567_7;

Selector_2 s2567_7(wires_641_6[3], addr_641_6, addr_positional[10271:10268], addr_2567_7);

wire[31:0] addr_2568_7;

Selector_2 s2568_7(wires_642_6[0], addr_642_6, addr_positional[10275:10272], addr_2568_7);

wire[31:0] addr_2569_7;

Selector_2 s2569_7(wires_642_6[1], addr_642_6, addr_positional[10279:10276], addr_2569_7);

wire[31:0] addr_2570_7;

Selector_2 s2570_7(wires_642_6[2], addr_642_6, addr_positional[10283:10280], addr_2570_7);

wire[31:0] addr_2571_7;

Selector_2 s2571_7(wires_642_6[3], addr_642_6, addr_positional[10287:10284], addr_2571_7);

wire[31:0] addr_2572_7;

Selector_2 s2572_7(wires_643_6[0], addr_643_6, addr_positional[10291:10288], addr_2572_7);

wire[31:0] addr_2573_7;

Selector_2 s2573_7(wires_643_6[1], addr_643_6, addr_positional[10295:10292], addr_2573_7);

wire[31:0] addr_2574_7;

Selector_2 s2574_7(wires_643_6[2], addr_643_6, addr_positional[10299:10296], addr_2574_7);

wire[31:0] addr_2575_7;

Selector_2 s2575_7(wires_643_6[3], addr_643_6, addr_positional[10303:10300], addr_2575_7);

wire[31:0] addr_2576_7;

Selector_2 s2576_7(wires_644_6[0], addr_644_6, addr_positional[10307:10304], addr_2576_7);

wire[31:0] addr_2577_7;

Selector_2 s2577_7(wires_644_6[1], addr_644_6, addr_positional[10311:10308], addr_2577_7);

wire[31:0] addr_2578_7;

Selector_2 s2578_7(wires_644_6[2], addr_644_6, addr_positional[10315:10312], addr_2578_7);

wire[31:0] addr_2579_7;

Selector_2 s2579_7(wires_644_6[3], addr_644_6, addr_positional[10319:10316], addr_2579_7);

wire[31:0] addr_2580_7;

Selector_2 s2580_7(wires_645_6[0], addr_645_6, addr_positional[10323:10320], addr_2580_7);

wire[31:0] addr_2581_7;

Selector_2 s2581_7(wires_645_6[1], addr_645_6, addr_positional[10327:10324], addr_2581_7);

wire[31:0] addr_2582_7;

Selector_2 s2582_7(wires_645_6[2], addr_645_6, addr_positional[10331:10328], addr_2582_7);

wire[31:0] addr_2583_7;

Selector_2 s2583_7(wires_645_6[3], addr_645_6, addr_positional[10335:10332], addr_2583_7);

wire[31:0] addr_2584_7;

Selector_2 s2584_7(wires_646_6[0], addr_646_6, addr_positional[10339:10336], addr_2584_7);

wire[31:0] addr_2585_7;

Selector_2 s2585_7(wires_646_6[1], addr_646_6, addr_positional[10343:10340], addr_2585_7);

wire[31:0] addr_2586_7;

Selector_2 s2586_7(wires_646_6[2], addr_646_6, addr_positional[10347:10344], addr_2586_7);

wire[31:0] addr_2587_7;

Selector_2 s2587_7(wires_646_6[3], addr_646_6, addr_positional[10351:10348], addr_2587_7);

wire[31:0] addr_2588_7;

Selector_2 s2588_7(wires_647_6[0], addr_647_6, addr_positional[10355:10352], addr_2588_7);

wire[31:0] addr_2589_7;

Selector_2 s2589_7(wires_647_6[1], addr_647_6, addr_positional[10359:10356], addr_2589_7);

wire[31:0] addr_2590_7;

Selector_2 s2590_7(wires_647_6[2], addr_647_6, addr_positional[10363:10360], addr_2590_7);

wire[31:0] addr_2591_7;

Selector_2 s2591_7(wires_647_6[3], addr_647_6, addr_positional[10367:10364], addr_2591_7);

wire[31:0] addr_2592_7;

Selector_2 s2592_7(wires_648_6[0], addr_648_6, addr_positional[10371:10368], addr_2592_7);

wire[31:0] addr_2593_7;

Selector_2 s2593_7(wires_648_6[1], addr_648_6, addr_positional[10375:10372], addr_2593_7);

wire[31:0] addr_2594_7;

Selector_2 s2594_7(wires_648_6[2], addr_648_6, addr_positional[10379:10376], addr_2594_7);

wire[31:0] addr_2595_7;

Selector_2 s2595_7(wires_648_6[3], addr_648_6, addr_positional[10383:10380], addr_2595_7);

wire[31:0] addr_2596_7;

Selector_2 s2596_7(wires_649_6[0], addr_649_6, addr_positional[10387:10384], addr_2596_7);

wire[31:0] addr_2597_7;

Selector_2 s2597_7(wires_649_6[1], addr_649_6, addr_positional[10391:10388], addr_2597_7);

wire[31:0] addr_2598_7;

Selector_2 s2598_7(wires_649_6[2], addr_649_6, addr_positional[10395:10392], addr_2598_7);

wire[31:0] addr_2599_7;

Selector_2 s2599_7(wires_649_6[3], addr_649_6, addr_positional[10399:10396], addr_2599_7);

wire[31:0] addr_2600_7;

Selector_2 s2600_7(wires_650_6[0], addr_650_6, addr_positional[10403:10400], addr_2600_7);

wire[31:0] addr_2601_7;

Selector_2 s2601_7(wires_650_6[1], addr_650_6, addr_positional[10407:10404], addr_2601_7);

wire[31:0] addr_2602_7;

Selector_2 s2602_7(wires_650_6[2], addr_650_6, addr_positional[10411:10408], addr_2602_7);

wire[31:0] addr_2603_7;

Selector_2 s2603_7(wires_650_6[3], addr_650_6, addr_positional[10415:10412], addr_2603_7);

wire[31:0] addr_2604_7;

Selector_2 s2604_7(wires_651_6[0], addr_651_6, addr_positional[10419:10416], addr_2604_7);

wire[31:0] addr_2605_7;

Selector_2 s2605_7(wires_651_6[1], addr_651_6, addr_positional[10423:10420], addr_2605_7);

wire[31:0] addr_2606_7;

Selector_2 s2606_7(wires_651_6[2], addr_651_6, addr_positional[10427:10424], addr_2606_7);

wire[31:0] addr_2607_7;

Selector_2 s2607_7(wires_651_6[3], addr_651_6, addr_positional[10431:10428], addr_2607_7);

wire[31:0] addr_2608_7;

Selector_2 s2608_7(wires_652_6[0], addr_652_6, addr_positional[10435:10432], addr_2608_7);

wire[31:0] addr_2609_7;

Selector_2 s2609_7(wires_652_6[1], addr_652_6, addr_positional[10439:10436], addr_2609_7);

wire[31:0] addr_2610_7;

Selector_2 s2610_7(wires_652_6[2], addr_652_6, addr_positional[10443:10440], addr_2610_7);

wire[31:0] addr_2611_7;

Selector_2 s2611_7(wires_652_6[3], addr_652_6, addr_positional[10447:10444], addr_2611_7);

wire[31:0] addr_2612_7;

Selector_2 s2612_7(wires_653_6[0], addr_653_6, addr_positional[10451:10448], addr_2612_7);

wire[31:0] addr_2613_7;

Selector_2 s2613_7(wires_653_6[1], addr_653_6, addr_positional[10455:10452], addr_2613_7);

wire[31:0] addr_2614_7;

Selector_2 s2614_7(wires_653_6[2], addr_653_6, addr_positional[10459:10456], addr_2614_7);

wire[31:0] addr_2615_7;

Selector_2 s2615_7(wires_653_6[3], addr_653_6, addr_positional[10463:10460], addr_2615_7);

wire[31:0] addr_2616_7;

Selector_2 s2616_7(wires_654_6[0], addr_654_6, addr_positional[10467:10464], addr_2616_7);

wire[31:0] addr_2617_7;

Selector_2 s2617_7(wires_654_6[1], addr_654_6, addr_positional[10471:10468], addr_2617_7);

wire[31:0] addr_2618_7;

Selector_2 s2618_7(wires_654_6[2], addr_654_6, addr_positional[10475:10472], addr_2618_7);

wire[31:0] addr_2619_7;

Selector_2 s2619_7(wires_654_6[3], addr_654_6, addr_positional[10479:10476], addr_2619_7);

wire[31:0] addr_2620_7;

Selector_2 s2620_7(wires_655_6[0], addr_655_6, addr_positional[10483:10480], addr_2620_7);

wire[31:0] addr_2621_7;

Selector_2 s2621_7(wires_655_6[1], addr_655_6, addr_positional[10487:10484], addr_2621_7);

wire[31:0] addr_2622_7;

Selector_2 s2622_7(wires_655_6[2], addr_655_6, addr_positional[10491:10488], addr_2622_7);

wire[31:0] addr_2623_7;

Selector_2 s2623_7(wires_655_6[3], addr_655_6, addr_positional[10495:10492], addr_2623_7);

wire[31:0] addr_2624_7;

Selector_2 s2624_7(wires_656_6[0], addr_656_6, addr_positional[10499:10496], addr_2624_7);

wire[31:0] addr_2625_7;

Selector_2 s2625_7(wires_656_6[1], addr_656_6, addr_positional[10503:10500], addr_2625_7);

wire[31:0] addr_2626_7;

Selector_2 s2626_7(wires_656_6[2], addr_656_6, addr_positional[10507:10504], addr_2626_7);

wire[31:0] addr_2627_7;

Selector_2 s2627_7(wires_656_6[3], addr_656_6, addr_positional[10511:10508], addr_2627_7);

wire[31:0] addr_2628_7;

Selector_2 s2628_7(wires_657_6[0], addr_657_6, addr_positional[10515:10512], addr_2628_7);

wire[31:0] addr_2629_7;

Selector_2 s2629_7(wires_657_6[1], addr_657_6, addr_positional[10519:10516], addr_2629_7);

wire[31:0] addr_2630_7;

Selector_2 s2630_7(wires_657_6[2], addr_657_6, addr_positional[10523:10520], addr_2630_7);

wire[31:0] addr_2631_7;

Selector_2 s2631_7(wires_657_6[3], addr_657_6, addr_positional[10527:10524], addr_2631_7);

wire[31:0] addr_2632_7;

Selector_2 s2632_7(wires_658_6[0], addr_658_6, addr_positional[10531:10528], addr_2632_7);

wire[31:0] addr_2633_7;

Selector_2 s2633_7(wires_658_6[1], addr_658_6, addr_positional[10535:10532], addr_2633_7);

wire[31:0] addr_2634_7;

Selector_2 s2634_7(wires_658_6[2], addr_658_6, addr_positional[10539:10536], addr_2634_7);

wire[31:0] addr_2635_7;

Selector_2 s2635_7(wires_658_6[3], addr_658_6, addr_positional[10543:10540], addr_2635_7);

wire[31:0] addr_2636_7;

Selector_2 s2636_7(wires_659_6[0], addr_659_6, addr_positional[10547:10544], addr_2636_7);

wire[31:0] addr_2637_7;

Selector_2 s2637_7(wires_659_6[1], addr_659_6, addr_positional[10551:10548], addr_2637_7);

wire[31:0] addr_2638_7;

Selector_2 s2638_7(wires_659_6[2], addr_659_6, addr_positional[10555:10552], addr_2638_7);

wire[31:0] addr_2639_7;

Selector_2 s2639_7(wires_659_6[3], addr_659_6, addr_positional[10559:10556], addr_2639_7);

wire[31:0] addr_2640_7;

Selector_2 s2640_7(wires_660_6[0], addr_660_6, addr_positional[10563:10560], addr_2640_7);

wire[31:0] addr_2641_7;

Selector_2 s2641_7(wires_660_6[1], addr_660_6, addr_positional[10567:10564], addr_2641_7);

wire[31:0] addr_2642_7;

Selector_2 s2642_7(wires_660_6[2], addr_660_6, addr_positional[10571:10568], addr_2642_7);

wire[31:0] addr_2643_7;

Selector_2 s2643_7(wires_660_6[3], addr_660_6, addr_positional[10575:10572], addr_2643_7);

wire[31:0] addr_2644_7;

Selector_2 s2644_7(wires_661_6[0], addr_661_6, addr_positional[10579:10576], addr_2644_7);

wire[31:0] addr_2645_7;

Selector_2 s2645_7(wires_661_6[1], addr_661_6, addr_positional[10583:10580], addr_2645_7);

wire[31:0] addr_2646_7;

Selector_2 s2646_7(wires_661_6[2], addr_661_6, addr_positional[10587:10584], addr_2646_7);

wire[31:0] addr_2647_7;

Selector_2 s2647_7(wires_661_6[3], addr_661_6, addr_positional[10591:10588], addr_2647_7);

wire[31:0] addr_2648_7;

Selector_2 s2648_7(wires_662_6[0], addr_662_6, addr_positional[10595:10592], addr_2648_7);

wire[31:0] addr_2649_7;

Selector_2 s2649_7(wires_662_6[1], addr_662_6, addr_positional[10599:10596], addr_2649_7);

wire[31:0] addr_2650_7;

Selector_2 s2650_7(wires_662_6[2], addr_662_6, addr_positional[10603:10600], addr_2650_7);

wire[31:0] addr_2651_7;

Selector_2 s2651_7(wires_662_6[3], addr_662_6, addr_positional[10607:10604], addr_2651_7);

wire[31:0] addr_2652_7;

Selector_2 s2652_7(wires_663_6[0], addr_663_6, addr_positional[10611:10608], addr_2652_7);

wire[31:0] addr_2653_7;

Selector_2 s2653_7(wires_663_6[1], addr_663_6, addr_positional[10615:10612], addr_2653_7);

wire[31:0] addr_2654_7;

Selector_2 s2654_7(wires_663_6[2], addr_663_6, addr_positional[10619:10616], addr_2654_7);

wire[31:0] addr_2655_7;

Selector_2 s2655_7(wires_663_6[3], addr_663_6, addr_positional[10623:10620], addr_2655_7);

wire[31:0] addr_2656_7;

Selector_2 s2656_7(wires_664_6[0], addr_664_6, addr_positional[10627:10624], addr_2656_7);

wire[31:0] addr_2657_7;

Selector_2 s2657_7(wires_664_6[1], addr_664_6, addr_positional[10631:10628], addr_2657_7);

wire[31:0] addr_2658_7;

Selector_2 s2658_7(wires_664_6[2], addr_664_6, addr_positional[10635:10632], addr_2658_7);

wire[31:0] addr_2659_7;

Selector_2 s2659_7(wires_664_6[3], addr_664_6, addr_positional[10639:10636], addr_2659_7);

wire[31:0] addr_2660_7;

Selector_2 s2660_7(wires_665_6[0], addr_665_6, addr_positional[10643:10640], addr_2660_7);

wire[31:0] addr_2661_7;

Selector_2 s2661_7(wires_665_6[1], addr_665_6, addr_positional[10647:10644], addr_2661_7);

wire[31:0] addr_2662_7;

Selector_2 s2662_7(wires_665_6[2], addr_665_6, addr_positional[10651:10648], addr_2662_7);

wire[31:0] addr_2663_7;

Selector_2 s2663_7(wires_665_6[3], addr_665_6, addr_positional[10655:10652], addr_2663_7);

wire[31:0] addr_2664_7;

Selector_2 s2664_7(wires_666_6[0], addr_666_6, addr_positional[10659:10656], addr_2664_7);

wire[31:0] addr_2665_7;

Selector_2 s2665_7(wires_666_6[1], addr_666_6, addr_positional[10663:10660], addr_2665_7);

wire[31:0] addr_2666_7;

Selector_2 s2666_7(wires_666_6[2], addr_666_6, addr_positional[10667:10664], addr_2666_7);

wire[31:0] addr_2667_7;

Selector_2 s2667_7(wires_666_6[3], addr_666_6, addr_positional[10671:10668], addr_2667_7);

wire[31:0] addr_2668_7;

Selector_2 s2668_7(wires_667_6[0], addr_667_6, addr_positional[10675:10672], addr_2668_7);

wire[31:0] addr_2669_7;

Selector_2 s2669_7(wires_667_6[1], addr_667_6, addr_positional[10679:10676], addr_2669_7);

wire[31:0] addr_2670_7;

Selector_2 s2670_7(wires_667_6[2], addr_667_6, addr_positional[10683:10680], addr_2670_7);

wire[31:0] addr_2671_7;

Selector_2 s2671_7(wires_667_6[3], addr_667_6, addr_positional[10687:10684], addr_2671_7);

wire[31:0] addr_2672_7;

Selector_2 s2672_7(wires_668_6[0], addr_668_6, addr_positional[10691:10688], addr_2672_7);

wire[31:0] addr_2673_7;

Selector_2 s2673_7(wires_668_6[1], addr_668_6, addr_positional[10695:10692], addr_2673_7);

wire[31:0] addr_2674_7;

Selector_2 s2674_7(wires_668_6[2], addr_668_6, addr_positional[10699:10696], addr_2674_7);

wire[31:0] addr_2675_7;

Selector_2 s2675_7(wires_668_6[3], addr_668_6, addr_positional[10703:10700], addr_2675_7);

wire[31:0] addr_2676_7;

Selector_2 s2676_7(wires_669_6[0], addr_669_6, addr_positional[10707:10704], addr_2676_7);

wire[31:0] addr_2677_7;

Selector_2 s2677_7(wires_669_6[1], addr_669_6, addr_positional[10711:10708], addr_2677_7);

wire[31:0] addr_2678_7;

Selector_2 s2678_7(wires_669_6[2], addr_669_6, addr_positional[10715:10712], addr_2678_7);

wire[31:0] addr_2679_7;

Selector_2 s2679_7(wires_669_6[3], addr_669_6, addr_positional[10719:10716], addr_2679_7);

wire[31:0] addr_2680_7;

Selector_2 s2680_7(wires_670_6[0], addr_670_6, addr_positional[10723:10720], addr_2680_7);

wire[31:0] addr_2681_7;

Selector_2 s2681_7(wires_670_6[1], addr_670_6, addr_positional[10727:10724], addr_2681_7);

wire[31:0] addr_2682_7;

Selector_2 s2682_7(wires_670_6[2], addr_670_6, addr_positional[10731:10728], addr_2682_7);

wire[31:0] addr_2683_7;

Selector_2 s2683_7(wires_670_6[3], addr_670_6, addr_positional[10735:10732], addr_2683_7);

wire[31:0] addr_2684_7;

Selector_2 s2684_7(wires_671_6[0], addr_671_6, addr_positional[10739:10736], addr_2684_7);

wire[31:0] addr_2685_7;

Selector_2 s2685_7(wires_671_6[1], addr_671_6, addr_positional[10743:10740], addr_2685_7);

wire[31:0] addr_2686_7;

Selector_2 s2686_7(wires_671_6[2], addr_671_6, addr_positional[10747:10744], addr_2686_7);

wire[31:0] addr_2687_7;

Selector_2 s2687_7(wires_671_6[3], addr_671_6, addr_positional[10751:10748], addr_2687_7);

wire[31:0] addr_2688_7;

Selector_2 s2688_7(wires_672_6[0], addr_672_6, addr_positional[10755:10752], addr_2688_7);

wire[31:0] addr_2689_7;

Selector_2 s2689_7(wires_672_6[1], addr_672_6, addr_positional[10759:10756], addr_2689_7);

wire[31:0] addr_2690_7;

Selector_2 s2690_7(wires_672_6[2], addr_672_6, addr_positional[10763:10760], addr_2690_7);

wire[31:0] addr_2691_7;

Selector_2 s2691_7(wires_672_6[3], addr_672_6, addr_positional[10767:10764], addr_2691_7);

wire[31:0] addr_2692_7;

Selector_2 s2692_7(wires_673_6[0], addr_673_6, addr_positional[10771:10768], addr_2692_7);

wire[31:0] addr_2693_7;

Selector_2 s2693_7(wires_673_6[1], addr_673_6, addr_positional[10775:10772], addr_2693_7);

wire[31:0] addr_2694_7;

Selector_2 s2694_7(wires_673_6[2], addr_673_6, addr_positional[10779:10776], addr_2694_7);

wire[31:0] addr_2695_7;

Selector_2 s2695_7(wires_673_6[3], addr_673_6, addr_positional[10783:10780], addr_2695_7);

wire[31:0] addr_2696_7;

Selector_2 s2696_7(wires_674_6[0], addr_674_6, addr_positional[10787:10784], addr_2696_7);

wire[31:0] addr_2697_7;

Selector_2 s2697_7(wires_674_6[1], addr_674_6, addr_positional[10791:10788], addr_2697_7);

wire[31:0] addr_2698_7;

Selector_2 s2698_7(wires_674_6[2], addr_674_6, addr_positional[10795:10792], addr_2698_7);

wire[31:0] addr_2699_7;

Selector_2 s2699_7(wires_674_6[3], addr_674_6, addr_positional[10799:10796], addr_2699_7);

wire[31:0] addr_2700_7;

Selector_2 s2700_7(wires_675_6[0], addr_675_6, addr_positional[10803:10800], addr_2700_7);

wire[31:0] addr_2701_7;

Selector_2 s2701_7(wires_675_6[1], addr_675_6, addr_positional[10807:10804], addr_2701_7);

wire[31:0] addr_2702_7;

Selector_2 s2702_7(wires_675_6[2], addr_675_6, addr_positional[10811:10808], addr_2702_7);

wire[31:0] addr_2703_7;

Selector_2 s2703_7(wires_675_6[3], addr_675_6, addr_positional[10815:10812], addr_2703_7);

wire[31:0] addr_2704_7;

Selector_2 s2704_7(wires_676_6[0], addr_676_6, addr_positional[10819:10816], addr_2704_7);

wire[31:0] addr_2705_7;

Selector_2 s2705_7(wires_676_6[1], addr_676_6, addr_positional[10823:10820], addr_2705_7);

wire[31:0] addr_2706_7;

Selector_2 s2706_7(wires_676_6[2], addr_676_6, addr_positional[10827:10824], addr_2706_7);

wire[31:0] addr_2707_7;

Selector_2 s2707_7(wires_676_6[3], addr_676_6, addr_positional[10831:10828], addr_2707_7);

wire[31:0] addr_2708_7;

Selector_2 s2708_7(wires_677_6[0], addr_677_6, addr_positional[10835:10832], addr_2708_7);

wire[31:0] addr_2709_7;

Selector_2 s2709_7(wires_677_6[1], addr_677_6, addr_positional[10839:10836], addr_2709_7);

wire[31:0] addr_2710_7;

Selector_2 s2710_7(wires_677_6[2], addr_677_6, addr_positional[10843:10840], addr_2710_7);

wire[31:0] addr_2711_7;

Selector_2 s2711_7(wires_677_6[3], addr_677_6, addr_positional[10847:10844], addr_2711_7);

wire[31:0] addr_2712_7;

Selector_2 s2712_7(wires_678_6[0], addr_678_6, addr_positional[10851:10848], addr_2712_7);

wire[31:0] addr_2713_7;

Selector_2 s2713_7(wires_678_6[1], addr_678_6, addr_positional[10855:10852], addr_2713_7);

wire[31:0] addr_2714_7;

Selector_2 s2714_7(wires_678_6[2], addr_678_6, addr_positional[10859:10856], addr_2714_7);

wire[31:0] addr_2715_7;

Selector_2 s2715_7(wires_678_6[3], addr_678_6, addr_positional[10863:10860], addr_2715_7);

wire[31:0] addr_2716_7;

Selector_2 s2716_7(wires_679_6[0], addr_679_6, addr_positional[10867:10864], addr_2716_7);

wire[31:0] addr_2717_7;

Selector_2 s2717_7(wires_679_6[1], addr_679_6, addr_positional[10871:10868], addr_2717_7);

wire[31:0] addr_2718_7;

Selector_2 s2718_7(wires_679_6[2], addr_679_6, addr_positional[10875:10872], addr_2718_7);

wire[31:0] addr_2719_7;

Selector_2 s2719_7(wires_679_6[3], addr_679_6, addr_positional[10879:10876], addr_2719_7);

wire[31:0] addr_2720_7;

Selector_2 s2720_7(wires_680_6[0], addr_680_6, addr_positional[10883:10880], addr_2720_7);

wire[31:0] addr_2721_7;

Selector_2 s2721_7(wires_680_6[1], addr_680_6, addr_positional[10887:10884], addr_2721_7);

wire[31:0] addr_2722_7;

Selector_2 s2722_7(wires_680_6[2], addr_680_6, addr_positional[10891:10888], addr_2722_7);

wire[31:0] addr_2723_7;

Selector_2 s2723_7(wires_680_6[3], addr_680_6, addr_positional[10895:10892], addr_2723_7);

wire[31:0] addr_2724_7;

Selector_2 s2724_7(wires_681_6[0], addr_681_6, addr_positional[10899:10896], addr_2724_7);

wire[31:0] addr_2725_7;

Selector_2 s2725_7(wires_681_6[1], addr_681_6, addr_positional[10903:10900], addr_2725_7);

wire[31:0] addr_2726_7;

Selector_2 s2726_7(wires_681_6[2], addr_681_6, addr_positional[10907:10904], addr_2726_7);

wire[31:0] addr_2727_7;

Selector_2 s2727_7(wires_681_6[3], addr_681_6, addr_positional[10911:10908], addr_2727_7);

wire[31:0] addr_2728_7;

Selector_2 s2728_7(wires_682_6[0], addr_682_6, addr_positional[10915:10912], addr_2728_7);

wire[31:0] addr_2729_7;

Selector_2 s2729_7(wires_682_6[1], addr_682_6, addr_positional[10919:10916], addr_2729_7);

wire[31:0] addr_2730_7;

Selector_2 s2730_7(wires_682_6[2], addr_682_6, addr_positional[10923:10920], addr_2730_7);

wire[31:0] addr_2731_7;

Selector_2 s2731_7(wires_682_6[3], addr_682_6, addr_positional[10927:10924], addr_2731_7);

wire[31:0] addr_2732_7;

Selector_2 s2732_7(wires_683_6[0], addr_683_6, addr_positional[10931:10928], addr_2732_7);

wire[31:0] addr_2733_7;

Selector_2 s2733_7(wires_683_6[1], addr_683_6, addr_positional[10935:10932], addr_2733_7);

wire[31:0] addr_2734_7;

Selector_2 s2734_7(wires_683_6[2], addr_683_6, addr_positional[10939:10936], addr_2734_7);

wire[31:0] addr_2735_7;

Selector_2 s2735_7(wires_683_6[3], addr_683_6, addr_positional[10943:10940], addr_2735_7);

wire[31:0] addr_2736_7;

Selector_2 s2736_7(wires_684_6[0], addr_684_6, addr_positional[10947:10944], addr_2736_7);

wire[31:0] addr_2737_7;

Selector_2 s2737_7(wires_684_6[1], addr_684_6, addr_positional[10951:10948], addr_2737_7);

wire[31:0] addr_2738_7;

Selector_2 s2738_7(wires_684_6[2], addr_684_6, addr_positional[10955:10952], addr_2738_7);

wire[31:0] addr_2739_7;

Selector_2 s2739_7(wires_684_6[3], addr_684_6, addr_positional[10959:10956], addr_2739_7);

wire[31:0] addr_2740_7;

Selector_2 s2740_7(wires_685_6[0], addr_685_6, addr_positional[10963:10960], addr_2740_7);

wire[31:0] addr_2741_7;

Selector_2 s2741_7(wires_685_6[1], addr_685_6, addr_positional[10967:10964], addr_2741_7);

wire[31:0] addr_2742_7;

Selector_2 s2742_7(wires_685_6[2], addr_685_6, addr_positional[10971:10968], addr_2742_7);

wire[31:0] addr_2743_7;

Selector_2 s2743_7(wires_685_6[3], addr_685_6, addr_positional[10975:10972], addr_2743_7);

wire[31:0] addr_2744_7;

Selector_2 s2744_7(wires_686_6[0], addr_686_6, addr_positional[10979:10976], addr_2744_7);

wire[31:0] addr_2745_7;

Selector_2 s2745_7(wires_686_6[1], addr_686_6, addr_positional[10983:10980], addr_2745_7);

wire[31:0] addr_2746_7;

Selector_2 s2746_7(wires_686_6[2], addr_686_6, addr_positional[10987:10984], addr_2746_7);

wire[31:0] addr_2747_7;

Selector_2 s2747_7(wires_686_6[3], addr_686_6, addr_positional[10991:10988], addr_2747_7);

wire[31:0] addr_2748_7;

Selector_2 s2748_7(wires_687_6[0], addr_687_6, addr_positional[10995:10992], addr_2748_7);

wire[31:0] addr_2749_7;

Selector_2 s2749_7(wires_687_6[1], addr_687_6, addr_positional[10999:10996], addr_2749_7);

wire[31:0] addr_2750_7;

Selector_2 s2750_7(wires_687_6[2], addr_687_6, addr_positional[11003:11000], addr_2750_7);

wire[31:0] addr_2751_7;

Selector_2 s2751_7(wires_687_6[3], addr_687_6, addr_positional[11007:11004], addr_2751_7);

wire[31:0] addr_2752_7;

Selector_2 s2752_7(wires_688_6[0], addr_688_6, addr_positional[11011:11008], addr_2752_7);

wire[31:0] addr_2753_7;

Selector_2 s2753_7(wires_688_6[1], addr_688_6, addr_positional[11015:11012], addr_2753_7);

wire[31:0] addr_2754_7;

Selector_2 s2754_7(wires_688_6[2], addr_688_6, addr_positional[11019:11016], addr_2754_7);

wire[31:0] addr_2755_7;

Selector_2 s2755_7(wires_688_6[3], addr_688_6, addr_positional[11023:11020], addr_2755_7);

wire[31:0] addr_2756_7;

Selector_2 s2756_7(wires_689_6[0], addr_689_6, addr_positional[11027:11024], addr_2756_7);

wire[31:0] addr_2757_7;

Selector_2 s2757_7(wires_689_6[1], addr_689_6, addr_positional[11031:11028], addr_2757_7);

wire[31:0] addr_2758_7;

Selector_2 s2758_7(wires_689_6[2], addr_689_6, addr_positional[11035:11032], addr_2758_7);

wire[31:0] addr_2759_7;

Selector_2 s2759_7(wires_689_6[3], addr_689_6, addr_positional[11039:11036], addr_2759_7);

wire[31:0] addr_2760_7;

Selector_2 s2760_7(wires_690_6[0], addr_690_6, addr_positional[11043:11040], addr_2760_7);

wire[31:0] addr_2761_7;

Selector_2 s2761_7(wires_690_6[1], addr_690_6, addr_positional[11047:11044], addr_2761_7);

wire[31:0] addr_2762_7;

Selector_2 s2762_7(wires_690_6[2], addr_690_6, addr_positional[11051:11048], addr_2762_7);

wire[31:0] addr_2763_7;

Selector_2 s2763_7(wires_690_6[3], addr_690_6, addr_positional[11055:11052], addr_2763_7);

wire[31:0] addr_2764_7;

Selector_2 s2764_7(wires_691_6[0], addr_691_6, addr_positional[11059:11056], addr_2764_7);

wire[31:0] addr_2765_7;

Selector_2 s2765_7(wires_691_6[1], addr_691_6, addr_positional[11063:11060], addr_2765_7);

wire[31:0] addr_2766_7;

Selector_2 s2766_7(wires_691_6[2], addr_691_6, addr_positional[11067:11064], addr_2766_7);

wire[31:0] addr_2767_7;

Selector_2 s2767_7(wires_691_6[3], addr_691_6, addr_positional[11071:11068], addr_2767_7);

wire[31:0] addr_2768_7;

Selector_2 s2768_7(wires_692_6[0], addr_692_6, addr_positional[11075:11072], addr_2768_7);

wire[31:0] addr_2769_7;

Selector_2 s2769_7(wires_692_6[1], addr_692_6, addr_positional[11079:11076], addr_2769_7);

wire[31:0] addr_2770_7;

Selector_2 s2770_7(wires_692_6[2], addr_692_6, addr_positional[11083:11080], addr_2770_7);

wire[31:0] addr_2771_7;

Selector_2 s2771_7(wires_692_6[3], addr_692_6, addr_positional[11087:11084], addr_2771_7);

wire[31:0] addr_2772_7;

Selector_2 s2772_7(wires_693_6[0], addr_693_6, addr_positional[11091:11088], addr_2772_7);

wire[31:0] addr_2773_7;

Selector_2 s2773_7(wires_693_6[1], addr_693_6, addr_positional[11095:11092], addr_2773_7);

wire[31:0] addr_2774_7;

Selector_2 s2774_7(wires_693_6[2], addr_693_6, addr_positional[11099:11096], addr_2774_7);

wire[31:0] addr_2775_7;

Selector_2 s2775_7(wires_693_6[3], addr_693_6, addr_positional[11103:11100], addr_2775_7);

wire[31:0] addr_2776_7;

Selector_2 s2776_7(wires_694_6[0], addr_694_6, addr_positional[11107:11104], addr_2776_7);

wire[31:0] addr_2777_7;

Selector_2 s2777_7(wires_694_6[1], addr_694_6, addr_positional[11111:11108], addr_2777_7);

wire[31:0] addr_2778_7;

Selector_2 s2778_7(wires_694_6[2], addr_694_6, addr_positional[11115:11112], addr_2778_7);

wire[31:0] addr_2779_7;

Selector_2 s2779_7(wires_694_6[3], addr_694_6, addr_positional[11119:11116], addr_2779_7);

wire[31:0] addr_2780_7;

Selector_2 s2780_7(wires_695_6[0], addr_695_6, addr_positional[11123:11120], addr_2780_7);

wire[31:0] addr_2781_7;

Selector_2 s2781_7(wires_695_6[1], addr_695_6, addr_positional[11127:11124], addr_2781_7);

wire[31:0] addr_2782_7;

Selector_2 s2782_7(wires_695_6[2], addr_695_6, addr_positional[11131:11128], addr_2782_7);

wire[31:0] addr_2783_7;

Selector_2 s2783_7(wires_695_6[3], addr_695_6, addr_positional[11135:11132], addr_2783_7);

wire[31:0] addr_2784_7;

Selector_2 s2784_7(wires_696_6[0], addr_696_6, addr_positional[11139:11136], addr_2784_7);

wire[31:0] addr_2785_7;

Selector_2 s2785_7(wires_696_6[1], addr_696_6, addr_positional[11143:11140], addr_2785_7);

wire[31:0] addr_2786_7;

Selector_2 s2786_7(wires_696_6[2], addr_696_6, addr_positional[11147:11144], addr_2786_7);

wire[31:0] addr_2787_7;

Selector_2 s2787_7(wires_696_6[3], addr_696_6, addr_positional[11151:11148], addr_2787_7);

wire[31:0] addr_2788_7;

Selector_2 s2788_7(wires_697_6[0], addr_697_6, addr_positional[11155:11152], addr_2788_7);

wire[31:0] addr_2789_7;

Selector_2 s2789_7(wires_697_6[1], addr_697_6, addr_positional[11159:11156], addr_2789_7);

wire[31:0] addr_2790_7;

Selector_2 s2790_7(wires_697_6[2], addr_697_6, addr_positional[11163:11160], addr_2790_7);

wire[31:0] addr_2791_7;

Selector_2 s2791_7(wires_697_6[3], addr_697_6, addr_positional[11167:11164], addr_2791_7);

wire[31:0] addr_2792_7;

Selector_2 s2792_7(wires_698_6[0], addr_698_6, addr_positional[11171:11168], addr_2792_7);

wire[31:0] addr_2793_7;

Selector_2 s2793_7(wires_698_6[1], addr_698_6, addr_positional[11175:11172], addr_2793_7);

wire[31:0] addr_2794_7;

Selector_2 s2794_7(wires_698_6[2], addr_698_6, addr_positional[11179:11176], addr_2794_7);

wire[31:0] addr_2795_7;

Selector_2 s2795_7(wires_698_6[3], addr_698_6, addr_positional[11183:11180], addr_2795_7);

wire[31:0] addr_2796_7;

Selector_2 s2796_7(wires_699_6[0], addr_699_6, addr_positional[11187:11184], addr_2796_7);

wire[31:0] addr_2797_7;

Selector_2 s2797_7(wires_699_6[1], addr_699_6, addr_positional[11191:11188], addr_2797_7);

wire[31:0] addr_2798_7;

Selector_2 s2798_7(wires_699_6[2], addr_699_6, addr_positional[11195:11192], addr_2798_7);

wire[31:0] addr_2799_7;

Selector_2 s2799_7(wires_699_6[3], addr_699_6, addr_positional[11199:11196], addr_2799_7);

wire[31:0] addr_2800_7;

Selector_2 s2800_7(wires_700_6[0], addr_700_6, addr_positional[11203:11200], addr_2800_7);

wire[31:0] addr_2801_7;

Selector_2 s2801_7(wires_700_6[1], addr_700_6, addr_positional[11207:11204], addr_2801_7);

wire[31:0] addr_2802_7;

Selector_2 s2802_7(wires_700_6[2], addr_700_6, addr_positional[11211:11208], addr_2802_7);

wire[31:0] addr_2803_7;

Selector_2 s2803_7(wires_700_6[3], addr_700_6, addr_positional[11215:11212], addr_2803_7);

wire[31:0] addr_2804_7;

Selector_2 s2804_7(wires_701_6[0], addr_701_6, addr_positional[11219:11216], addr_2804_7);

wire[31:0] addr_2805_7;

Selector_2 s2805_7(wires_701_6[1], addr_701_6, addr_positional[11223:11220], addr_2805_7);

wire[31:0] addr_2806_7;

Selector_2 s2806_7(wires_701_6[2], addr_701_6, addr_positional[11227:11224], addr_2806_7);

wire[31:0] addr_2807_7;

Selector_2 s2807_7(wires_701_6[3], addr_701_6, addr_positional[11231:11228], addr_2807_7);

wire[31:0] addr_2808_7;

Selector_2 s2808_7(wires_702_6[0], addr_702_6, addr_positional[11235:11232], addr_2808_7);

wire[31:0] addr_2809_7;

Selector_2 s2809_7(wires_702_6[1], addr_702_6, addr_positional[11239:11236], addr_2809_7);

wire[31:0] addr_2810_7;

Selector_2 s2810_7(wires_702_6[2], addr_702_6, addr_positional[11243:11240], addr_2810_7);

wire[31:0] addr_2811_7;

Selector_2 s2811_7(wires_702_6[3], addr_702_6, addr_positional[11247:11244], addr_2811_7);

wire[31:0] addr_2812_7;

Selector_2 s2812_7(wires_703_6[0], addr_703_6, addr_positional[11251:11248], addr_2812_7);

wire[31:0] addr_2813_7;

Selector_2 s2813_7(wires_703_6[1], addr_703_6, addr_positional[11255:11252], addr_2813_7);

wire[31:0] addr_2814_7;

Selector_2 s2814_7(wires_703_6[2], addr_703_6, addr_positional[11259:11256], addr_2814_7);

wire[31:0] addr_2815_7;

Selector_2 s2815_7(wires_703_6[3], addr_703_6, addr_positional[11263:11260], addr_2815_7);

wire[31:0] addr_2816_7;

Selector_2 s2816_7(wires_704_6[0], addr_704_6, addr_positional[11267:11264], addr_2816_7);

wire[31:0] addr_2817_7;

Selector_2 s2817_7(wires_704_6[1], addr_704_6, addr_positional[11271:11268], addr_2817_7);

wire[31:0] addr_2818_7;

Selector_2 s2818_7(wires_704_6[2], addr_704_6, addr_positional[11275:11272], addr_2818_7);

wire[31:0] addr_2819_7;

Selector_2 s2819_7(wires_704_6[3], addr_704_6, addr_positional[11279:11276], addr_2819_7);

wire[31:0] addr_2820_7;

Selector_2 s2820_7(wires_705_6[0], addr_705_6, addr_positional[11283:11280], addr_2820_7);

wire[31:0] addr_2821_7;

Selector_2 s2821_7(wires_705_6[1], addr_705_6, addr_positional[11287:11284], addr_2821_7);

wire[31:0] addr_2822_7;

Selector_2 s2822_7(wires_705_6[2], addr_705_6, addr_positional[11291:11288], addr_2822_7);

wire[31:0] addr_2823_7;

Selector_2 s2823_7(wires_705_6[3], addr_705_6, addr_positional[11295:11292], addr_2823_7);

wire[31:0] addr_2824_7;

Selector_2 s2824_7(wires_706_6[0], addr_706_6, addr_positional[11299:11296], addr_2824_7);

wire[31:0] addr_2825_7;

Selector_2 s2825_7(wires_706_6[1], addr_706_6, addr_positional[11303:11300], addr_2825_7);

wire[31:0] addr_2826_7;

Selector_2 s2826_7(wires_706_6[2], addr_706_6, addr_positional[11307:11304], addr_2826_7);

wire[31:0] addr_2827_7;

Selector_2 s2827_7(wires_706_6[3], addr_706_6, addr_positional[11311:11308], addr_2827_7);

wire[31:0] addr_2828_7;

Selector_2 s2828_7(wires_707_6[0], addr_707_6, addr_positional[11315:11312], addr_2828_7);

wire[31:0] addr_2829_7;

Selector_2 s2829_7(wires_707_6[1], addr_707_6, addr_positional[11319:11316], addr_2829_7);

wire[31:0] addr_2830_7;

Selector_2 s2830_7(wires_707_6[2], addr_707_6, addr_positional[11323:11320], addr_2830_7);

wire[31:0] addr_2831_7;

Selector_2 s2831_7(wires_707_6[3], addr_707_6, addr_positional[11327:11324], addr_2831_7);

wire[31:0] addr_2832_7;

Selector_2 s2832_7(wires_708_6[0], addr_708_6, addr_positional[11331:11328], addr_2832_7);

wire[31:0] addr_2833_7;

Selector_2 s2833_7(wires_708_6[1], addr_708_6, addr_positional[11335:11332], addr_2833_7);

wire[31:0] addr_2834_7;

Selector_2 s2834_7(wires_708_6[2], addr_708_6, addr_positional[11339:11336], addr_2834_7);

wire[31:0] addr_2835_7;

Selector_2 s2835_7(wires_708_6[3], addr_708_6, addr_positional[11343:11340], addr_2835_7);

wire[31:0] addr_2836_7;

Selector_2 s2836_7(wires_709_6[0], addr_709_6, addr_positional[11347:11344], addr_2836_7);

wire[31:0] addr_2837_7;

Selector_2 s2837_7(wires_709_6[1], addr_709_6, addr_positional[11351:11348], addr_2837_7);

wire[31:0] addr_2838_7;

Selector_2 s2838_7(wires_709_6[2], addr_709_6, addr_positional[11355:11352], addr_2838_7);

wire[31:0] addr_2839_7;

Selector_2 s2839_7(wires_709_6[3], addr_709_6, addr_positional[11359:11356], addr_2839_7);

wire[31:0] addr_2840_7;

Selector_2 s2840_7(wires_710_6[0], addr_710_6, addr_positional[11363:11360], addr_2840_7);

wire[31:0] addr_2841_7;

Selector_2 s2841_7(wires_710_6[1], addr_710_6, addr_positional[11367:11364], addr_2841_7);

wire[31:0] addr_2842_7;

Selector_2 s2842_7(wires_710_6[2], addr_710_6, addr_positional[11371:11368], addr_2842_7);

wire[31:0] addr_2843_7;

Selector_2 s2843_7(wires_710_6[3], addr_710_6, addr_positional[11375:11372], addr_2843_7);

wire[31:0] addr_2844_7;

Selector_2 s2844_7(wires_711_6[0], addr_711_6, addr_positional[11379:11376], addr_2844_7);

wire[31:0] addr_2845_7;

Selector_2 s2845_7(wires_711_6[1], addr_711_6, addr_positional[11383:11380], addr_2845_7);

wire[31:0] addr_2846_7;

Selector_2 s2846_7(wires_711_6[2], addr_711_6, addr_positional[11387:11384], addr_2846_7);

wire[31:0] addr_2847_7;

Selector_2 s2847_7(wires_711_6[3], addr_711_6, addr_positional[11391:11388], addr_2847_7);

wire[31:0] addr_2848_7;

Selector_2 s2848_7(wires_712_6[0], addr_712_6, addr_positional[11395:11392], addr_2848_7);

wire[31:0] addr_2849_7;

Selector_2 s2849_7(wires_712_6[1], addr_712_6, addr_positional[11399:11396], addr_2849_7);

wire[31:0] addr_2850_7;

Selector_2 s2850_7(wires_712_6[2], addr_712_6, addr_positional[11403:11400], addr_2850_7);

wire[31:0] addr_2851_7;

Selector_2 s2851_7(wires_712_6[3], addr_712_6, addr_positional[11407:11404], addr_2851_7);

wire[31:0] addr_2852_7;

Selector_2 s2852_7(wires_713_6[0], addr_713_6, addr_positional[11411:11408], addr_2852_7);

wire[31:0] addr_2853_7;

Selector_2 s2853_7(wires_713_6[1], addr_713_6, addr_positional[11415:11412], addr_2853_7);

wire[31:0] addr_2854_7;

Selector_2 s2854_7(wires_713_6[2], addr_713_6, addr_positional[11419:11416], addr_2854_7);

wire[31:0] addr_2855_7;

Selector_2 s2855_7(wires_713_6[3], addr_713_6, addr_positional[11423:11420], addr_2855_7);

wire[31:0] addr_2856_7;

Selector_2 s2856_7(wires_714_6[0], addr_714_6, addr_positional[11427:11424], addr_2856_7);

wire[31:0] addr_2857_7;

Selector_2 s2857_7(wires_714_6[1], addr_714_6, addr_positional[11431:11428], addr_2857_7);

wire[31:0] addr_2858_7;

Selector_2 s2858_7(wires_714_6[2], addr_714_6, addr_positional[11435:11432], addr_2858_7);

wire[31:0] addr_2859_7;

Selector_2 s2859_7(wires_714_6[3], addr_714_6, addr_positional[11439:11436], addr_2859_7);

wire[31:0] addr_2860_7;

Selector_2 s2860_7(wires_715_6[0], addr_715_6, addr_positional[11443:11440], addr_2860_7);

wire[31:0] addr_2861_7;

Selector_2 s2861_7(wires_715_6[1], addr_715_6, addr_positional[11447:11444], addr_2861_7);

wire[31:0] addr_2862_7;

Selector_2 s2862_7(wires_715_6[2], addr_715_6, addr_positional[11451:11448], addr_2862_7);

wire[31:0] addr_2863_7;

Selector_2 s2863_7(wires_715_6[3], addr_715_6, addr_positional[11455:11452], addr_2863_7);

wire[31:0] addr_2864_7;

Selector_2 s2864_7(wires_716_6[0], addr_716_6, addr_positional[11459:11456], addr_2864_7);

wire[31:0] addr_2865_7;

Selector_2 s2865_7(wires_716_6[1], addr_716_6, addr_positional[11463:11460], addr_2865_7);

wire[31:0] addr_2866_7;

Selector_2 s2866_7(wires_716_6[2], addr_716_6, addr_positional[11467:11464], addr_2866_7);

wire[31:0] addr_2867_7;

Selector_2 s2867_7(wires_716_6[3], addr_716_6, addr_positional[11471:11468], addr_2867_7);

wire[31:0] addr_2868_7;

Selector_2 s2868_7(wires_717_6[0], addr_717_6, addr_positional[11475:11472], addr_2868_7);

wire[31:0] addr_2869_7;

Selector_2 s2869_7(wires_717_6[1], addr_717_6, addr_positional[11479:11476], addr_2869_7);

wire[31:0] addr_2870_7;

Selector_2 s2870_7(wires_717_6[2], addr_717_6, addr_positional[11483:11480], addr_2870_7);

wire[31:0] addr_2871_7;

Selector_2 s2871_7(wires_717_6[3], addr_717_6, addr_positional[11487:11484], addr_2871_7);

wire[31:0] addr_2872_7;

Selector_2 s2872_7(wires_718_6[0], addr_718_6, addr_positional[11491:11488], addr_2872_7);

wire[31:0] addr_2873_7;

Selector_2 s2873_7(wires_718_6[1], addr_718_6, addr_positional[11495:11492], addr_2873_7);

wire[31:0] addr_2874_7;

Selector_2 s2874_7(wires_718_6[2], addr_718_6, addr_positional[11499:11496], addr_2874_7);

wire[31:0] addr_2875_7;

Selector_2 s2875_7(wires_718_6[3], addr_718_6, addr_positional[11503:11500], addr_2875_7);

wire[31:0] addr_2876_7;

Selector_2 s2876_7(wires_719_6[0], addr_719_6, addr_positional[11507:11504], addr_2876_7);

wire[31:0] addr_2877_7;

Selector_2 s2877_7(wires_719_6[1], addr_719_6, addr_positional[11511:11508], addr_2877_7);

wire[31:0] addr_2878_7;

Selector_2 s2878_7(wires_719_6[2], addr_719_6, addr_positional[11515:11512], addr_2878_7);

wire[31:0] addr_2879_7;

Selector_2 s2879_7(wires_719_6[3], addr_719_6, addr_positional[11519:11516], addr_2879_7);

wire[31:0] addr_2880_7;

Selector_2 s2880_7(wires_720_6[0], addr_720_6, addr_positional[11523:11520], addr_2880_7);

wire[31:0] addr_2881_7;

Selector_2 s2881_7(wires_720_6[1], addr_720_6, addr_positional[11527:11524], addr_2881_7);

wire[31:0] addr_2882_7;

Selector_2 s2882_7(wires_720_6[2], addr_720_6, addr_positional[11531:11528], addr_2882_7);

wire[31:0] addr_2883_7;

Selector_2 s2883_7(wires_720_6[3], addr_720_6, addr_positional[11535:11532], addr_2883_7);

wire[31:0] addr_2884_7;

Selector_2 s2884_7(wires_721_6[0], addr_721_6, addr_positional[11539:11536], addr_2884_7);

wire[31:0] addr_2885_7;

Selector_2 s2885_7(wires_721_6[1], addr_721_6, addr_positional[11543:11540], addr_2885_7);

wire[31:0] addr_2886_7;

Selector_2 s2886_7(wires_721_6[2], addr_721_6, addr_positional[11547:11544], addr_2886_7);

wire[31:0] addr_2887_7;

Selector_2 s2887_7(wires_721_6[3], addr_721_6, addr_positional[11551:11548], addr_2887_7);

wire[31:0] addr_2888_7;

Selector_2 s2888_7(wires_722_6[0], addr_722_6, addr_positional[11555:11552], addr_2888_7);

wire[31:0] addr_2889_7;

Selector_2 s2889_7(wires_722_6[1], addr_722_6, addr_positional[11559:11556], addr_2889_7);

wire[31:0] addr_2890_7;

Selector_2 s2890_7(wires_722_6[2], addr_722_6, addr_positional[11563:11560], addr_2890_7);

wire[31:0] addr_2891_7;

Selector_2 s2891_7(wires_722_6[3], addr_722_6, addr_positional[11567:11564], addr_2891_7);

wire[31:0] addr_2892_7;

Selector_2 s2892_7(wires_723_6[0], addr_723_6, addr_positional[11571:11568], addr_2892_7);

wire[31:0] addr_2893_7;

Selector_2 s2893_7(wires_723_6[1], addr_723_6, addr_positional[11575:11572], addr_2893_7);

wire[31:0] addr_2894_7;

Selector_2 s2894_7(wires_723_6[2], addr_723_6, addr_positional[11579:11576], addr_2894_7);

wire[31:0] addr_2895_7;

Selector_2 s2895_7(wires_723_6[3], addr_723_6, addr_positional[11583:11580], addr_2895_7);

wire[31:0] addr_2896_7;

Selector_2 s2896_7(wires_724_6[0], addr_724_6, addr_positional[11587:11584], addr_2896_7);

wire[31:0] addr_2897_7;

Selector_2 s2897_7(wires_724_6[1], addr_724_6, addr_positional[11591:11588], addr_2897_7);

wire[31:0] addr_2898_7;

Selector_2 s2898_7(wires_724_6[2], addr_724_6, addr_positional[11595:11592], addr_2898_7);

wire[31:0] addr_2899_7;

Selector_2 s2899_7(wires_724_6[3], addr_724_6, addr_positional[11599:11596], addr_2899_7);

wire[31:0] addr_2900_7;

Selector_2 s2900_7(wires_725_6[0], addr_725_6, addr_positional[11603:11600], addr_2900_7);

wire[31:0] addr_2901_7;

Selector_2 s2901_7(wires_725_6[1], addr_725_6, addr_positional[11607:11604], addr_2901_7);

wire[31:0] addr_2902_7;

Selector_2 s2902_7(wires_725_6[2], addr_725_6, addr_positional[11611:11608], addr_2902_7);

wire[31:0] addr_2903_7;

Selector_2 s2903_7(wires_725_6[3], addr_725_6, addr_positional[11615:11612], addr_2903_7);

wire[31:0] addr_2904_7;

Selector_2 s2904_7(wires_726_6[0], addr_726_6, addr_positional[11619:11616], addr_2904_7);

wire[31:0] addr_2905_7;

Selector_2 s2905_7(wires_726_6[1], addr_726_6, addr_positional[11623:11620], addr_2905_7);

wire[31:0] addr_2906_7;

Selector_2 s2906_7(wires_726_6[2], addr_726_6, addr_positional[11627:11624], addr_2906_7);

wire[31:0] addr_2907_7;

Selector_2 s2907_7(wires_726_6[3], addr_726_6, addr_positional[11631:11628], addr_2907_7);

wire[31:0] addr_2908_7;

Selector_2 s2908_7(wires_727_6[0], addr_727_6, addr_positional[11635:11632], addr_2908_7);

wire[31:0] addr_2909_7;

Selector_2 s2909_7(wires_727_6[1], addr_727_6, addr_positional[11639:11636], addr_2909_7);

wire[31:0] addr_2910_7;

Selector_2 s2910_7(wires_727_6[2], addr_727_6, addr_positional[11643:11640], addr_2910_7);

wire[31:0] addr_2911_7;

Selector_2 s2911_7(wires_727_6[3], addr_727_6, addr_positional[11647:11644], addr_2911_7);

wire[31:0] addr_2912_7;

Selector_2 s2912_7(wires_728_6[0], addr_728_6, addr_positional[11651:11648], addr_2912_7);

wire[31:0] addr_2913_7;

Selector_2 s2913_7(wires_728_6[1], addr_728_6, addr_positional[11655:11652], addr_2913_7);

wire[31:0] addr_2914_7;

Selector_2 s2914_7(wires_728_6[2], addr_728_6, addr_positional[11659:11656], addr_2914_7);

wire[31:0] addr_2915_7;

Selector_2 s2915_7(wires_728_6[3], addr_728_6, addr_positional[11663:11660], addr_2915_7);

wire[31:0] addr_2916_7;

Selector_2 s2916_7(wires_729_6[0], addr_729_6, addr_positional[11667:11664], addr_2916_7);

wire[31:0] addr_2917_7;

Selector_2 s2917_7(wires_729_6[1], addr_729_6, addr_positional[11671:11668], addr_2917_7);

wire[31:0] addr_2918_7;

Selector_2 s2918_7(wires_729_6[2], addr_729_6, addr_positional[11675:11672], addr_2918_7);

wire[31:0] addr_2919_7;

Selector_2 s2919_7(wires_729_6[3], addr_729_6, addr_positional[11679:11676], addr_2919_7);

wire[31:0] addr_2920_7;

Selector_2 s2920_7(wires_730_6[0], addr_730_6, addr_positional[11683:11680], addr_2920_7);

wire[31:0] addr_2921_7;

Selector_2 s2921_7(wires_730_6[1], addr_730_6, addr_positional[11687:11684], addr_2921_7);

wire[31:0] addr_2922_7;

Selector_2 s2922_7(wires_730_6[2], addr_730_6, addr_positional[11691:11688], addr_2922_7);

wire[31:0] addr_2923_7;

Selector_2 s2923_7(wires_730_6[3], addr_730_6, addr_positional[11695:11692], addr_2923_7);

wire[31:0] addr_2924_7;

Selector_2 s2924_7(wires_731_6[0], addr_731_6, addr_positional[11699:11696], addr_2924_7);

wire[31:0] addr_2925_7;

Selector_2 s2925_7(wires_731_6[1], addr_731_6, addr_positional[11703:11700], addr_2925_7);

wire[31:0] addr_2926_7;

Selector_2 s2926_7(wires_731_6[2], addr_731_6, addr_positional[11707:11704], addr_2926_7);

wire[31:0] addr_2927_7;

Selector_2 s2927_7(wires_731_6[3], addr_731_6, addr_positional[11711:11708], addr_2927_7);

wire[31:0] addr_2928_7;

Selector_2 s2928_7(wires_732_6[0], addr_732_6, addr_positional[11715:11712], addr_2928_7);

wire[31:0] addr_2929_7;

Selector_2 s2929_7(wires_732_6[1], addr_732_6, addr_positional[11719:11716], addr_2929_7);

wire[31:0] addr_2930_7;

Selector_2 s2930_7(wires_732_6[2], addr_732_6, addr_positional[11723:11720], addr_2930_7);

wire[31:0] addr_2931_7;

Selector_2 s2931_7(wires_732_6[3], addr_732_6, addr_positional[11727:11724], addr_2931_7);

wire[31:0] addr_2932_7;

Selector_2 s2932_7(wires_733_6[0], addr_733_6, addr_positional[11731:11728], addr_2932_7);

wire[31:0] addr_2933_7;

Selector_2 s2933_7(wires_733_6[1], addr_733_6, addr_positional[11735:11732], addr_2933_7);

wire[31:0] addr_2934_7;

Selector_2 s2934_7(wires_733_6[2], addr_733_6, addr_positional[11739:11736], addr_2934_7);

wire[31:0] addr_2935_7;

Selector_2 s2935_7(wires_733_6[3], addr_733_6, addr_positional[11743:11740], addr_2935_7);

wire[31:0] addr_2936_7;

Selector_2 s2936_7(wires_734_6[0], addr_734_6, addr_positional[11747:11744], addr_2936_7);

wire[31:0] addr_2937_7;

Selector_2 s2937_7(wires_734_6[1], addr_734_6, addr_positional[11751:11748], addr_2937_7);

wire[31:0] addr_2938_7;

Selector_2 s2938_7(wires_734_6[2], addr_734_6, addr_positional[11755:11752], addr_2938_7);

wire[31:0] addr_2939_7;

Selector_2 s2939_7(wires_734_6[3], addr_734_6, addr_positional[11759:11756], addr_2939_7);

wire[31:0] addr_2940_7;

Selector_2 s2940_7(wires_735_6[0], addr_735_6, addr_positional[11763:11760], addr_2940_7);

wire[31:0] addr_2941_7;

Selector_2 s2941_7(wires_735_6[1], addr_735_6, addr_positional[11767:11764], addr_2941_7);

wire[31:0] addr_2942_7;

Selector_2 s2942_7(wires_735_6[2], addr_735_6, addr_positional[11771:11768], addr_2942_7);

wire[31:0] addr_2943_7;

Selector_2 s2943_7(wires_735_6[3], addr_735_6, addr_positional[11775:11772], addr_2943_7);

wire[31:0] addr_2944_7;

Selector_2 s2944_7(wires_736_6[0], addr_736_6, addr_positional[11779:11776], addr_2944_7);

wire[31:0] addr_2945_7;

Selector_2 s2945_7(wires_736_6[1], addr_736_6, addr_positional[11783:11780], addr_2945_7);

wire[31:0] addr_2946_7;

Selector_2 s2946_7(wires_736_6[2], addr_736_6, addr_positional[11787:11784], addr_2946_7);

wire[31:0] addr_2947_7;

Selector_2 s2947_7(wires_736_6[3], addr_736_6, addr_positional[11791:11788], addr_2947_7);

wire[31:0] addr_2948_7;

Selector_2 s2948_7(wires_737_6[0], addr_737_6, addr_positional[11795:11792], addr_2948_7);

wire[31:0] addr_2949_7;

Selector_2 s2949_7(wires_737_6[1], addr_737_6, addr_positional[11799:11796], addr_2949_7);

wire[31:0] addr_2950_7;

Selector_2 s2950_7(wires_737_6[2], addr_737_6, addr_positional[11803:11800], addr_2950_7);

wire[31:0] addr_2951_7;

Selector_2 s2951_7(wires_737_6[3], addr_737_6, addr_positional[11807:11804], addr_2951_7);

wire[31:0] addr_2952_7;

Selector_2 s2952_7(wires_738_6[0], addr_738_6, addr_positional[11811:11808], addr_2952_7);

wire[31:0] addr_2953_7;

Selector_2 s2953_7(wires_738_6[1], addr_738_6, addr_positional[11815:11812], addr_2953_7);

wire[31:0] addr_2954_7;

Selector_2 s2954_7(wires_738_6[2], addr_738_6, addr_positional[11819:11816], addr_2954_7);

wire[31:0] addr_2955_7;

Selector_2 s2955_7(wires_738_6[3], addr_738_6, addr_positional[11823:11820], addr_2955_7);

wire[31:0] addr_2956_7;

Selector_2 s2956_7(wires_739_6[0], addr_739_6, addr_positional[11827:11824], addr_2956_7);

wire[31:0] addr_2957_7;

Selector_2 s2957_7(wires_739_6[1], addr_739_6, addr_positional[11831:11828], addr_2957_7);

wire[31:0] addr_2958_7;

Selector_2 s2958_7(wires_739_6[2], addr_739_6, addr_positional[11835:11832], addr_2958_7);

wire[31:0] addr_2959_7;

Selector_2 s2959_7(wires_739_6[3], addr_739_6, addr_positional[11839:11836], addr_2959_7);

wire[31:0] addr_2960_7;

Selector_2 s2960_7(wires_740_6[0], addr_740_6, addr_positional[11843:11840], addr_2960_7);

wire[31:0] addr_2961_7;

Selector_2 s2961_7(wires_740_6[1], addr_740_6, addr_positional[11847:11844], addr_2961_7);

wire[31:0] addr_2962_7;

Selector_2 s2962_7(wires_740_6[2], addr_740_6, addr_positional[11851:11848], addr_2962_7);

wire[31:0] addr_2963_7;

Selector_2 s2963_7(wires_740_6[3], addr_740_6, addr_positional[11855:11852], addr_2963_7);

wire[31:0] addr_2964_7;

Selector_2 s2964_7(wires_741_6[0], addr_741_6, addr_positional[11859:11856], addr_2964_7);

wire[31:0] addr_2965_7;

Selector_2 s2965_7(wires_741_6[1], addr_741_6, addr_positional[11863:11860], addr_2965_7);

wire[31:0] addr_2966_7;

Selector_2 s2966_7(wires_741_6[2], addr_741_6, addr_positional[11867:11864], addr_2966_7);

wire[31:0] addr_2967_7;

Selector_2 s2967_7(wires_741_6[3], addr_741_6, addr_positional[11871:11868], addr_2967_7);

wire[31:0] addr_2968_7;

Selector_2 s2968_7(wires_742_6[0], addr_742_6, addr_positional[11875:11872], addr_2968_7);

wire[31:0] addr_2969_7;

Selector_2 s2969_7(wires_742_6[1], addr_742_6, addr_positional[11879:11876], addr_2969_7);

wire[31:0] addr_2970_7;

Selector_2 s2970_7(wires_742_6[2], addr_742_6, addr_positional[11883:11880], addr_2970_7);

wire[31:0] addr_2971_7;

Selector_2 s2971_7(wires_742_6[3], addr_742_6, addr_positional[11887:11884], addr_2971_7);

wire[31:0] addr_2972_7;

Selector_2 s2972_7(wires_743_6[0], addr_743_6, addr_positional[11891:11888], addr_2972_7);

wire[31:0] addr_2973_7;

Selector_2 s2973_7(wires_743_6[1], addr_743_6, addr_positional[11895:11892], addr_2973_7);

wire[31:0] addr_2974_7;

Selector_2 s2974_7(wires_743_6[2], addr_743_6, addr_positional[11899:11896], addr_2974_7);

wire[31:0] addr_2975_7;

Selector_2 s2975_7(wires_743_6[3], addr_743_6, addr_positional[11903:11900], addr_2975_7);

wire[31:0] addr_2976_7;

Selector_2 s2976_7(wires_744_6[0], addr_744_6, addr_positional[11907:11904], addr_2976_7);

wire[31:0] addr_2977_7;

Selector_2 s2977_7(wires_744_6[1], addr_744_6, addr_positional[11911:11908], addr_2977_7);

wire[31:0] addr_2978_7;

Selector_2 s2978_7(wires_744_6[2], addr_744_6, addr_positional[11915:11912], addr_2978_7);

wire[31:0] addr_2979_7;

Selector_2 s2979_7(wires_744_6[3], addr_744_6, addr_positional[11919:11916], addr_2979_7);

wire[31:0] addr_2980_7;

Selector_2 s2980_7(wires_745_6[0], addr_745_6, addr_positional[11923:11920], addr_2980_7);

wire[31:0] addr_2981_7;

Selector_2 s2981_7(wires_745_6[1], addr_745_6, addr_positional[11927:11924], addr_2981_7);

wire[31:0] addr_2982_7;

Selector_2 s2982_7(wires_745_6[2], addr_745_6, addr_positional[11931:11928], addr_2982_7);

wire[31:0] addr_2983_7;

Selector_2 s2983_7(wires_745_6[3], addr_745_6, addr_positional[11935:11932], addr_2983_7);

wire[31:0] addr_2984_7;

Selector_2 s2984_7(wires_746_6[0], addr_746_6, addr_positional[11939:11936], addr_2984_7);

wire[31:0] addr_2985_7;

Selector_2 s2985_7(wires_746_6[1], addr_746_6, addr_positional[11943:11940], addr_2985_7);

wire[31:0] addr_2986_7;

Selector_2 s2986_7(wires_746_6[2], addr_746_6, addr_positional[11947:11944], addr_2986_7);

wire[31:0] addr_2987_7;

Selector_2 s2987_7(wires_746_6[3], addr_746_6, addr_positional[11951:11948], addr_2987_7);

wire[31:0] addr_2988_7;

Selector_2 s2988_7(wires_747_6[0], addr_747_6, addr_positional[11955:11952], addr_2988_7);

wire[31:0] addr_2989_7;

Selector_2 s2989_7(wires_747_6[1], addr_747_6, addr_positional[11959:11956], addr_2989_7);

wire[31:0] addr_2990_7;

Selector_2 s2990_7(wires_747_6[2], addr_747_6, addr_positional[11963:11960], addr_2990_7);

wire[31:0] addr_2991_7;

Selector_2 s2991_7(wires_747_6[3], addr_747_6, addr_positional[11967:11964], addr_2991_7);

wire[31:0] addr_2992_7;

Selector_2 s2992_7(wires_748_6[0], addr_748_6, addr_positional[11971:11968], addr_2992_7);

wire[31:0] addr_2993_7;

Selector_2 s2993_7(wires_748_6[1], addr_748_6, addr_positional[11975:11972], addr_2993_7);

wire[31:0] addr_2994_7;

Selector_2 s2994_7(wires_748_6[2], addr_748_6, addr_positional[11979:11976], addr_2994_7);

wire[31:0] addr_2995_7;

Selector_2 s2995_7(wires_748_6[3], addr_748_6, addr_positional[11983:11980], addr_2995_7);

wire[31:0] addr_2996_7;

Selector_2 s2996_7(wires_749_6[0], addr_749_6, addr_positional[11987:11984], addr_2996_7);

wire[31:0] addr_2997_7;

Selector_2 s2997_7(wires_749_6[1], addr_749_6, addr_positional[11991:11988], addr_2997_7);

wire[31:0] addr_2998_7;

Selector_2 s2998_7(wires_749_6[2], addr_749_6, addr_positional[11995:11992], addr_2998_7);

wire[31:0] addr_2999_7;

Selector_2 s2999_7(wires_749_6[3], addr_749_6, addr_positional[11999:11996], addr_2999_7);

wire[31:0] addr_3000_7;

Selector_2 s3000_7(wires_750_6[0], addr_750_6, addr_positional[12003:12000], addr_3000_7);

wire[31:0] addr_3001_7;

Selector_2 s3001_7(wires_750_6[1], addr_750_6, addr_positional[12007:12004], addr_3001_7);

wire[31:0] addr_3002_7;

Selector_2 s3002_7(wires_750_6[2], addr_750_6, addr_positional[12011:12008], addr_3002_7);

wire[31:0] addr_3003_7;

Selector_2 s3003_7(wires_750_6[3], addr_750_6, addr_positional[12015:12012], addr_3003_7);

wire[31:0] addr_3004_7;

Selector_2 s3004_7(wires_751_6[0], addr_751_6, addr_positional[12019:12016], addr_3004_7);

wire[31:0] addr_3005_7;

Selector_2 s3005_7(wires_751_6[1], addr_751_6, addr_positional[12023:12020], addr_3005_7);

wire[31:0] addr_3006_7;

Selector_2 s3006_7(wires_751_6[2], addr_751_6, addr_positional[12027:12024], addr_3006_7);

wire[31:0] addr_3007_7;

Selector_2 s3007_7(wires_751_6[3], addr_751_6, addr_positional[12031:12028], addr_3007_7);

wire[31:0] addr_3008_7;

Selector_2 s3008_7(wires_752_6[0], addr_752_6, addr_positional[12035:12032], addr_3008_7);

wire[31:0] addr_3009_7;

Selector_2 s3009_7(wires_752_6[1], addr_752_6, addr_positional[12039:12036], addr_3009_7);

wire[31:0] addr_3010_7;

Selector_2 s3010_7(wires_752_6[2], addr_752_6, addr_positional[12043:12040], addr_3010_7);

wire[31:0] addr_3011_7;

Selector_2 s3011_7(wires_752_6[3], addr_752_6, addr_positional[12047:12044], addr_3011_7);

wire[31:0] addr_3012_7;

Selector_2 s3012_7(wires_753_6[0], addr_753_6, addr_positional[12051:12048], addr_3012_7);

wire[31:0] addr_3013_7;

Selector_2 s3013_7(wires_753_6[1], addr_753_6, addr_positional[12055:12052], addr_3013_7);

wire[31:0] addr_3014_7;

Selector_2 s3014_7(wires_753_6[2], addr_753_6, addr_positional[12059:12056], addr_3014_7);

wire[31:0] addr_3015_7;

Selector_2 s3015_7(wires_753_6[3], addr_753_6, addr_positional[12063:12060], addr_3015_7);

wire[31:0] addr_3016_7;

Selector_2 s3016_7(wires_754_6[0], addr_754_6, addr_positional[12067:12064], addr_3016_7);

wire[31:0] addr_3017_7;

Selector_2 s3017_7(wires_754_6[1], addr_754_6, addr_positional[12071:12068], addr_3017_7);

wire[31:0] addr_3018_7;

Selector_2 s3018_7(wires_754_6[2], addr_754_6, addr_positional[12075:12072], addr_3018_7);

wire[31:0] addr_3019_7;

Selector_2 s3019_7(wires_754_6[3], addr_754_6, addr_positional[12079:12076], addr_3019_7);

wire[31:0] addr_3020_7;

Selector_2 s3020_7(wires_755_6[0], addr_755_6, addr_positional[12083:12080], addr_3020_7);

wire[31:0] addr_3021_7;

Selector_2 s3021_7(wires_755_6[1], addr_755_6, addr_positional[12087:12084], addr_3021_7);

wire[31:0] addr_3022_7;

Selector_2 s3022_7(wires_755_6[2], addr_755_6, addr_positional[12091:12088], addr_3022_7);

wire[31:0] addr_3023_7;

Selector_2 s3023_7(wires_755_6[3], addr_755_6, addr_positional[12095:12092], addr_3023_7);

wire[31:0] addr_3024_7;

Selector_2 s3024_7(wires_756_6[0], addr_756_6, addr_positional[12099:12096], addr_3024_7);

wire[31:0] addr_3025_7;

Selector_2 s3025_7(wires_756_6[1], addr_756_6, addr_positional[12103:12100], addr_3025_7);

wire[31:0] addr_3026_7;

Selector_2 s3026_7(wires_756_6[2], addr_756_6, addr_positional[12107:12104], addr_3026_7);

wire[31:0] addr_3027_7;

Selector_2 s3027_7(wires_756_6[3], addr_756_6, addr_positional[12111:12108], addr_3027_7);

wire[31:0] addr_3028_7;

Selector_2 s3028_7(wires_757_6[0], addr_757_6, addr_positional[12115:12112], addr_3028_7);

wire[31:0] addr_3029_7;

Selector_2 s3029_7(wires_757_6[1], addr_757_6, addr_positional[12119:12116], addr_3029_7);

wire[31:0] addr_3030_7;

Selector_2 s3030_7(wires_757_6[2], addr_757_6, addr_positional[12123:12120], addr_3030_7);

wire[31:0] addr_3031_7;

Selector_2 s3031_7(wires_757_6[3], addr_757_6, addr_positional[12127:12124], addr_3031_7);

wire[31:0] addr_3032_7;

Selector_2 s3032_7(wires_758_6[0], addr_758_6, addr_positional[12131:12128], addr_3032_7);

wire[31:0] addr_3033_7;

Selector_2 s3033_7(wires_758_6[1], addr_758_6, addr_positional[12135:12132], addr_3033_7);

wire[31:0] addr_3034_7;

Selector_2 s3034_7(wires_758_6[2], addr_758_6, addr_positional[12139:12136], addr_3034_7);

wire[31:0] addr_3035_7;

Selector_2 s3035_7(wires_758_6[3], addr_758_6, addr_positional[12143:12140], addr_3035_7);

wire[31:0] addr_3036_7;

Selector_2 s3036_7(wires_759_6[0], addr_759_6, addr_positional[12147:12144], addr_3036_7);

wire[31:0] addr_3037_7;

Selector_2 s3037_7(wires_759_6[1], addr_759_6, addr_positional[12151:12148], addr_3037_7);

wire[31:0] addr_3038_7;

Selector_2 s3038_7(wires_759_6[2], addr_759_6, addr_positional[12155:12152], addr_3038_7);

wire[31:0] addr_3039_7;

Selector_2 s3039_7(wires_759_6[3], addr_759_6, addr_positional[12159:12156], addr_3039_7);

wire[31:0] addr_3040_7;

Selector_2 s3040_7(wires_760_6[0], addr_760_6, addr_positional[12163:12160], addr_3040_7);

wire[31:0] addr_3041_7;

Selector_2 s3041_7(wires_760_6[1], addr_760_6, addr_positional[12167:12164], addr_3041_7);

wire[31:0] addr_3042_7;

Selector_2 s3042_7(wires_760_6[2], addr_760_6, addr_positional[12171:12168], addr_3042_7);

wire[31:0] addr_3043_7;

Selector_2 s3043_7(wires_760_6[3], addr_760_6, addr_positional[12175:12172], addr_3043_7);

wire[31:0] addr_3044_7;

Selector_2 s3044_7(wires_761_6[0], addr_761_6, addr_positional[12179:12176], addr_3044_7);

wire[31:0] addr_3045_7;

Selector_2 s3045_7(wires_761_6[1], addr_761_6, addr_positional[12183:12180], addr_3045_7);

wire[31:0] addr_3046_7;

Selector_2 s3046_7(wires_761_6[2], addr_761_6, addr_positional[12187:12184], addr_3046_7);

wire[31:0] addr_3047_7;

Selector_2 s3047_7(wires_761_6[3], addr_761_6, addr_positional[12191:12188], addr_3047_7);

wire[31:0] addr_3048_7;

Selector_2 s3048_7(wires_762_6[0], addr_762_6, addr_positional[12195:12192], addr_3048_7);

wire[31:0] addr_3049_7;

Selector_2 s3049_7(wires_762_6[1], addr_762_6, addr_positional[12199:12196], addr_3049_7);

wire[31:0] addr_3050_7;

Selector_2 s3050_7(wires_762_6[2], addr_762_6, addr_positional[12203:12200], addr_3050_7);

wire[31:0] addr_3051_7;

Selector_2 s3051_7(wires_762_6[3], addr_762_6, addr_positional[12207:12204], addr_3051_7);

wire[31:0] addr_3052_7;

Selector_2 s3052_7(wires_763_6[0], addr_763_6, addr_positional[12211:12208], addr_3052_7);

wire[31:0] addr_3053_7;

Selector_2 s3053_7(wires_763_6[1], addr_763_6, addr_positional[12215:12212], addr_3053_7);

wire[31:0] addr_3054_7;

Selector_2 s3054_7(wires_763_6[2], addr_763_6, addr_positional[12219:12216], addr_3054_7);

wire[31:0] addr_3055_7;

Selector_2 s3055_7(wires_763_6[3], addr_763_6, addr_positional[12223:12220], addr_3055_7);

wire[31:0] addr_3056_7;

Selector_2 s3056_7(wires_764_6[0], addr_764_6, addr_positional[12227:12224], addr_3056_7);

wire[31:0] addr_3057_7;

Selector_2 s3057_7(wires_764_6[1], addr_764_6, addr_positional[12231:12228], addr_3057_7);

wire[31:0] addr_3058_7;

Selector_2 s3058_7(wires_764_6[2], addr_764_6, addr_positional[12235:12232], addr_3058_7);

wire[31:0] addr_3059_7;

Selector_2 s3059_7(wires_764_6[3], addr_764_6, addr_positional[12239:12236], addr_3059_7);

wire[31:0] addr_3060_7;

Selector_2 s3060_7(wires_765_6[0], addr_765_6, addr_positional[12243:12240], addr_3060_7);

wire[31:0] addr_3061_7;

Selector_2 s3061_7(wires_765_6[1], addr_765_6, addr_positional[12247:12244], addr_3061_7);

wire[31:0] addr_3062_7;

Selector_2 s3062_7(wires_765_6[2], addr_765_6, addr_positional[12251:12248], addr_3062_7);

wire[31:0] addr_3063_7;

Selector_2 s3063_7(wires_765_6[3], addr_765_6, addr_positional[12255:12252], addr_3063_7);

wire[31:0] addr_3064_7;

Selector_2 s3064_7(wires_766_6[0], addr_766_6, addr_positional[12259:12256], addr_3064_7);

wire[31:0] addr_3065_7;

Selector_2 s3065_7(wires_766_6[1], addr_766_6, addr_positional[12263:12260], addr_3065_7);

wire[31:0] addr_3066_7;

Selector_2 s3066_7(wires_766_6[2], addr_766_6, addr_positional[12267:12264], addr_3066_7);

wire[31:0] addr_3067_7;

Selector_2 s3067_7(wires_766_6[3], addr_766_6, addr_positional[12271:12268], addr_3067_7);

wire[31:0] addr_3068_7;

Selector_2 s3068_7(wires_767_6[0], addr_767_6, addr_positional[12275:12272], addr_3068_7);

wire[31:0] addr_3069_7;

Selector_2 s3069_7(wires_767_6[1], addr_767_6, addr_positional[12279:12276], addr_3069_7);

wire[31:0] addr_3070_7;

Selector_2 s3070_7(wires_767_6[2], addr_767_6, addr_positional[12283:12280], addr_3070_7);

wire[31:0] addr_3071_7;

Selector_2 s3071_7(wires_767_6[3], addr_767_6, addr_positional[12287:12284], addr_3071_7);

wire[31:0] addr_3072_7;

Selector_2 s3072_7(wires_768_6[0], addr_768_6, addr_positional[12291:12288], addr_3072_7);

wire[31:0] addr_3073_7;

Selector_2 s3073_7(wires_768_6[1], addr_768_6, addr_positional[12295:12292], addr_3073_7);

wire[31:0] addr_3074_7;

Selector_2 s3074_7(wires_768_6[2], addr_768_6, addr_positional[12299:12296], addr_3074_7);

wire[31:0] addr_3075_7;

Selector_2 s3075_7(wires_768_6[3], addr_768_6, addr_positional[12303:12300], addr_3075_7);

wire[31:0] addr_3076_7;

Selector_2 s3076_7(wires_769_6[0], addr_769_6, addr_positional[12307:12304], addr_3076_7);

wire[31:0] addr_3077_7;

Selector_2 s3077_7(wires_769_6[1], addr_769_6, addr_positional[12311:12308], addr_3077_7);

wire[31:0] addr_3078_7;

Selector_2 s3078_7(wires_769_6[2], addr_769_6, addr_positional[12315:12312], addr_3078_7);

wire[31:0] addr_3079_7;

Selector_2 s3079_7(wires_769_6[3], addr_769_6, addr_positional[12319:12316], addr_3079_7);

wire[31:0] addr_3080_7;

Selector_2 s3080_7(wires_770_6[0], addr_770_6, addr_positional[12323:12320], addr_3080_7);

wire[31:0] addr_3081_7;

Selector_2 s3081_7(wires_770_6[1], addr_770_6, addr_positional[12327:12324], addr_3081_7);

wire[31:0] addr_3082_7;

Selector_2 s3082_7(wires_770_6[2], addr_770_6, addr_positional[12331:12328], addr_3082_7);

wire[31:0] addr_3083_7;

Selector_2 s3083_7(wires_770_6[3], addr_770_6, addr_positional[12335:12332], addr_3083_7);

wire[31:0] addr_3084_7;

Selector_2 s3084_7(wires_771_6[0], addr_771_6, addr_positional[12339:12336], addr_3084_7);

wire[31:0] addr_3085_7;

Selector_2 s3085_7(wires_771_6[1], addr_771_6, addr_positional[12343:12340], addr_3085_7);

wire[31:0] addr_3086_7;

Selector_2 s3086_7(wires_771_6[2], addr_771_6, addr_positional[12347:12344], addr_3086_7);

wire[31:0] addr_3087_7;

Selector_2 s3087_7(wires_771_6[3], addr_771_6, addr_positional[12351:12348], addr_3087_7);

wire[31:0] addr_3088_7;

Selector_2 s3088_7(wires_772_6[0], addr_772_6, addr_positional[12355:12352], addr_3088_7);

wire[31:0] addr_3089_7;

Selector_2 s3089_7(wires_772_6[1], addr_772_6, addr_positional[12359:12356], addr_3089_7);

wire[31:0] addr_3090_7;

Selector_2 s3090_7(wires_772_6[2], addr_772_6, addr_positional[12363:12360], addr_3090_7);

wire[31:0] addr_3091_7;

Selector_2 s3091_7(wires_772_6[3], addr_772_6, addr_positional[12367:12364], addr_3091_7);

wire[31:0] addr_3092_7;

Selector_2 s3092_7(wires_773_6[0], addr_773_6, addr_positional[12371:12368], addr_3092_7);

wire[31:0] addr_3093_7;

Selector_2 s3093_7(wires_773_6[1], addr_773_6, addr_positional[12375:12372], addr_3093_7);

wire[31:0] addr_3094_7;

Selector_2 s3094_7(wires_773_6[2], addr_773_6, addr_positional[12379:12376], addr_3094_7);

wire[31:0] addr_3095_7;

Selector_2 s3095_7(wires_773_6[3], addr_773_6, addr_positional[12383:12380], addr_3095_7);

wire[31:0] addr_3096_7;

Selector_2 s3096_7(wires_774_6[0], addr_774_6, addr_positional[12387:12384], addr_3096_7);

wire[31:0] addr_3097_7;

Selector_2 s3097_7(wires_774_6[1], addr_774_6, addr_positional[12391:12388], addr_3097_7);

wire[31:0] addr_3098_7;

Selector_2 s3098_7(wires_774_6[2], addr_774_6, addr_positional[12395:12392], addr_3098_7);

wire[31:0] addr_3099_7;

Selector_2 s3099_7(wires_774_6[3], addr_774_6, addr_positional[12399:12396], addr_3099_7);

wire[31:0] addr_3100_7;

Selector_2 s3100_7(wires_775_6[0], addr_775_6, addr_positional[12403:12400], addr_3100_7);

wire[31:0] addr_3101_7;

Selector_2 s3101_7(wires_775_6[1], addr_775_6, addr_positional[12407:12404], addr_3101_7);

wire[31:0] addr_3102_7;

Selector_2 s3102_7(wires_775_6[2], addr_775_6, addr_positional[12411:12408], addr_3102_7);

wire[31:0] addr_3103_7;

Selector_2 s3103_7(wires_775_6[3], addr_775_6, addr_positional[12415:12412], addr_3103_7);

wire[31:0] addr_3104_7;

Selector_2 s3104_7(wires_776_6[0], addr_776_6, addr_positional[12419:12416], addr_3104_7);

wire[31:0] addr_3105_7;

Selector_2 s3105_7(wires_776_6[1], addr_776_6, addr_positional[12423:12420], addr_3105_7);

wire[31:0] addr_3106_7;

Selector_2 s3106_7(wires_776_6[2], addr_776_6, addr_positional[12427:12424], addr_3106_7);

wire[31:0] addr_3107_7;

Selector_2 s3107_7(wires_776_6[3], addr_776_6, addr_positional[12431:12428], addr_3107_7);

wire[31:0] addr_3108_7;

Selector_2 s3108_7(wires_777_6[0], addr_777_6, addr_positional[12435:12432], addr_3108_7);

wire[31:0] addr_3109_7;

Selector_2 s3109_7(wires_777_6[1], addr_777_6, addr_positional[12439:12436], addr_3109_7);

wire[31:0] addr_3110_7;

Selector_2 s3110_7(wires_777_6[2], addr_777_6, addr_positional[12443:12440], addr_3110_7);

wire[31:0] addr_3111_7;

Selector_2 s3111_7(wires_777_6[3], addr_777_6, addr_positional[12447:12444], addr_3111_7);

wire[31:0] addr_3112_7;

Selector_2 s3112_7(wires_778_6[0], addr_778_6, addr_positional[12451:12448], addr_3112_7);

wire[31:0] addr_3113_7;

Selector_2 s3113_7(wires_778_6[1], addr_778_6, addr_positional[12455:12452], addr_3113_7);

wire[31:0] addr_3114_7;

Selector_2 s3114_7(wires_778_6[2], addr_778_6, addr_positional[12459:12456], addr_3114_7);

wire[31:0] addr_3115_7;

Selector_2 s3115_7(wires_778_6[3], addr_778_6, addr_positional[12463:12460], addr_3115_7);

wire[31:0] addr_3116_7;

Selector_2 s3116_7(wires_779_6[0], addr_779_6, addr_positional[12467:12464], addr_3116_7);

wire[31:0] addr_3117_7;

Selector_2 s3117_7(wires_779_6[1], addr_779_6, addr_positional[12471:12468], addr_3117_7);

wire[31:0] addr_3118_7;

Selector_2 s3118_7(wires_779_6[2], addr_779_6, addr_positional[12475:12472], addr_3118_7);

wire[31:0] addr_3119_7;

Selector_2 s3119_7(wires_779_6[3], addr_779_6, addr_positional[12479:12476], addr_3119_7);

wire[31:0] addr_3120_7;

Selector_2 s3120_7(wires_780_6[0], addr_780_6, addr_positional[12483:12480], addr_3120_7);

wire[31:0] addr_3121_7;

Selector_2 s3121_7(wires_780_6[1], addr_780_6, addr_positional[12487:12484], addr_3121_7);

wire[31:0] addr_3122_7;

Selector_2 s3122_7(wires_780_6[2], addr_780_6, addr_positional[12491:12488], addr_3122_7);

wire[31:0] addr_3123_7;

Selector_2 s3123_7(wires_780_6[3], addr_780_6, addr_positional[12495:12492], addr_3123_7);

wire[31:0] addr_3124_7;

Selector_2 s3124_7(wires_781_6[0], addr_781_6, addr_positional[12499:12496], addr_3124_7);

wire[31:0] addr_3125_7;

Selector_2 s3125_7(wires_781_6[1], addr_781_6, addr_positional[12503:12500], addr_3125_7);

wire[31:0] addr_3126_7;

Selector_2 s3126_7(wires_781_6[2], addr_781_6, addr_positional[12507:12504], addr_3126_7);

wire[31:0] addr_3127_7;

Selector_2 s3127_7(wires_781_6[3], addr_781_6, addr_positional[12511:12508], addr_3127_7);

wire[31:0] addr_3128_7;

Selector_2 s3128_7(wires_782_6[0], addr_782_6, addr_positional[12515:12512], addr_3128_7);

wire[31:0] addr_3129_7;

Selector_2 s3129_7(wires_782_6[1], addr_782_6, addr_positional[12519:12516], addr_3129_7);

wire[31:0] addr_3130_7;

Selector_2 s3130_7(wires_782_6[2], addr_782_6, addr_positional[12523:12520], addr_3130_7);

wire[31:0] addr_3131_7;

Selector_2 s3131_7(wires_782_6[3], addr_782_6, addr_positional[12527:12524], addr_3131_7);

wire[31:0] addr_3132_7;

Selector_2 s3132_7(wires_783_6[0], addr_783_6, addr_positional[12531:12528], addr_3132_7);

wire[31:0] addr_3133_7;

Selector_2 s3133_7(wires_783_6[1], addr_783_6, addr_positional[12535:12532], addr_3133_7);

wire[31:0] addr_3134_7;

Selector_2 s3134_7(wires_783_6[2], addr_783_6, addr_positional[12539:12536], addr_3134_7);

wire[31:0] addr_3135_7;

Selector_2 s3135_7(wires_783_6[3], addr_783_6, addr_positional[12543:12540], addr_3135_7);

wire[31:0] addr_3136_7;

Selector_2 s3136_7(wires_784_6[0], addr_784_6, addr_positional[12547:12544], addr_3136_7);

wire[31:0] addr_3137_7;

Selector_2 s3137_7(wires_784_6[1], addr_784_6, addr_positional[12551:12548], addr_3137_7);

wire[31:0] addr_3138_7;

Selector_2 s3138_7(wires_784_6[2], addr_784_6, addr_positional[12555:12552], addr_3138_7);

wire[31:0] addr_3139_7;

Selector_2 s3139_7(wires_784_6[3], addr_784_6, addr_positional[12559:12556], addr_3139_7);

wire[31:0] addr_3140_7;

Selector_2 s3140_7(wires_785_6[0], addr_785_6, addr_positional[12563:12560], addr_3140_7);

wire[31:0] addr_3141_7;

Selector_2 s3141_7(wires_785_6[1], addr_785_6, addr_positional[12567:12564], addr_3141_7);

wire[31:0] addr_3142_7;

Selector_2 s3142_7(wires_785_6[2], addr_785_6, addr_positional[12571:12568], addr_3142_7);

wire[31:0] addr_3143_7;

Selector_2 s3143_7(wires_785_6[3], addr_785_6, addr_positional[12575:12572], addr_3143_7);

wire[31:0] addr_3144_7;

Selector_2 s3144_7(wires_786_6[0], addr_786_6, addr_positional[12579:12576], addr_3144_7);

wire[31:0] addr_3145_7;

Selector_2 s3145_7(wires_786_6[1], addr_786_6, addr_positional[12583:12580], addr_3145_7);

wire[31:0] addr_3146_7;

Selector_2 s3146_7(wires_786_6[2], addr_786_6, addr_positional[12587:12584], addr_3146_7);

wire[31:0] addr_3147_7;

Selector_2 s3147_7(wires_786_6[3], addr_786_6, addr_positional[12591:12588], addr_3147_7);

wire[31:0] addr_3148_7;

Selector_2 s3148_7(wires_787_6[0], addr_787_6, addr_positional[12595:12592], addr_3148_7);

wire[31:0] addr_3149_7;

Selector_2 s3149_7(wires_787_6[1], addr_787_6, addr_positional[12599:12596], addr_3149_7);

wire[31:0] addr_3150_7;

Selector_2 s3150_7(wires_787_6[2], addr_787_6, addr_positional[12603:12600], addr_3150_7);

wire[31:0] addr_3151_7;

Selector_2 s3151_7(wires_787_6[3], addr_787_6, addr_positional[12607:12604], addr_3151_7);

wire[31:0] addr_3152_7;

Selector_2 s3152_7(wires_788_6[0], addr_788_6, addr_positional[12611:12608], addr_3152_7);

wire[31:0] addr_3153_7;

Selector_2 s3153_7(wires_788_6[1], addr_788_6, addr_positional[12615:12612], addr_3153_7);

wire[31:0] addr_3154_7;

Selector_2 s3154_7(wires_788_6[2], addr_788_6, addr_positional[12619:12616], addr_3154_7);

wire[31:0] addr_3155_7;

Selector_2 s3155_7(wires_788_6[3], addr_788_6, addr_positional[12623:12620], addr_3155_7);

wire[31:0] addr_3156_7;

Selector_2 s3156_7(wires_789_6[0], addr_789_6, addr_positional[12627:12624], addr_3156_7);

wire[31:0] addr_3157_7;

Selector_2 s3157_7(wires_789_6[1], addr_789_6, addr_positional[12631:12628], addr_3157_7);

wire[31:0] addr_3158_7;

Selector_2 s3158_7(wires_789_6[2], addr_789_6, addr_positional[12635:12632], addr_3158_7);

wire[31:0] addr_3159_7;

Selector_2 s3159_7(wires_789_6[3], addr_789_6, addr_positional[12639:12636], addr_3159_7);

wire[31:0] addr_3160_7;

Selector_2 s3160_7(wires_790_6[0], addr_790_6, addr_positional[12643:12640], addr_3160_7);

wire[31:0] addr_3161_7;

Selector_2 s3161_7(wires_790_6[1], addr_790_6, addr_positional[12647:12644], addr_3161_7);

wire[31:0] addr_3162_7;

Selector_2 s3162_7(wires_790_6[2], addr_790_6, addr_positional[12651:12648], addr_3162_7);

wire[31:0] addr_3163_7;

Selector_2 s3163_7(wires_790_6[3], addr_790_6, addr_positional[12655:12652], addr_3163_7);

wire[31:0] addr_3164_7;

Selector_2 s3164_7(wires_791_6[0], addr_791_6, addr_positional[12659:12656], addr_3164_7);

wire[31:0] addr_3165_7;

Selector_2 s3165_7(wires_791_6[1], addr_791_6, addr_positional[12663:12660], addr_3165_7);

wire[31:0] addr_3166_7;

Selector_2 s3166_7(wires_791_6[2], addr_791_6, addr_positional[12667:12664], addr_3166_7);

wire[31:0] addr_3167_7;

Selector_2 s3167_7(wires_791_6[3], addr_791_6, addr_positional[12671:12668], addr_3167_7);

wire[31:0] addr_3168_7;

Selector_2 s3168_7(wires_792_6[0], addr_792_6, addr_positional[12675:12672], addr_3168_7);

wire[31:0] addr_3169_7;

Selector_2 s3169_7(wires_792_6[1], addr_792_6, addr_positional[12679:12676], addr_3169_7);

wire[31:0] addr_3170_7;

Selector_2 s3170_7(wires_792_6[2], addr_792_6, addr_positional[12683:12680], addr_3170_7);

wire[31:0] addr_3171_7;

Selector_2 s3171_7(wires_792_6[3], addr_792_6, addr_positional[12687:12684], addr_3171_7);

wire[31:0] addr_3172_7;

Selector_2 s3172_7(wires_793_6[0], addr_793_6, addr_positional[12691:12688], addr_3172_7);

wire[31:0] addr_3173_7;

Selector_2 s3173_7(wires_793_6[1], addr_793_6, addr_positional[12695:12692], addr_3173_7);

wire[31:0] addr_3174_7;

Selector_2 s3174_7(wires_793_6[2], addr_793_6, addr_positional[12699:12696], addr_3174_7);

wire[31:0] addr_3175_7;

Selector_2 s3175_7(wires_793_6[3], addr_793_6, addr_positional[12703:12700], addr_3175_7);

wire[31:0] addr_3176_7;

Selector_2 s3176_7(wires_794_6[0], addr_794_6, addr_positional[12707:12704], addr_3176_7);

wire[31:0] addr_3177_7;

Selector_2 s3177_7(wires_794_6[1], addr_794_6, addr_positional[12711:12708], addr_3177_7);

wire[31:0] addr_3178_7;

Selector_2 s3178_7(wires_794_6[2], addr_794_6, addr_positional[12715:12712], addr_3178_7);

wire[31:0] addr_3179_7;

Selector_2 s3179_7(wires_794_6[3], addr_794_6, addr_positional[12719:12716], addr_3179_7);

wire[31:0] addr_3180_7;

Selector_2 s3180_7(wires_795_6[0], addr_795_6, addr_positional[12723:12720], addr_3180_7);

wire[31:0] addr_3181_7;

Selector_2 s3181_7(wires_795_6[1], addr_795_6, addr_positional[12727:12724], addr_3181_7);

wire[31:0] addr_3182_7;

Selector_2 s3182_7(wires_795_6[2], addr_795_6, addr_positional[12731:12728], addr_3182_7);

wire[31:0] addr_3183_7;

Selector_2 s3183_7(wires_795_6[3], addr_795_6, addr_positional[12735:12732], addr_3183_7);

wire[31:0] addr_3184_7;

Selector_2 s3184_7(wires_796_6[0], addr_796_6, addr_positional[12739:12736], addr_3184_7);

wire[31:0] addr_3185_7;

Selector_2 s3185_7(wires_796_6[1], addr_796_6, addr_positional[12743:12740], addr_3185_7);

wire[31:0] addr_3186_7;

Selector_2 s3186_7(wires_796_6[2], addr_796_6, addr_positional[12747:12744], addr_3186_7);

wire[31:0] addr_3187_7;

Selector_2 s3187_7(wires_796_6[3], addr_796_6, addr_positional[12751:12748], addr_3187_7);

wire[31:0] addr_3188_7;

Selector_2 s3188_7(wires_797_6[0], addr_797_6, addr_positional[12755:12752], addr_3188_7);

wire[31:0] addr_3189_7;

Selector_2 s3189_7(wires_797_6[1], addr_797_6, addr_positional[12759:12756], addr_3189_7);

wire[31:0] addr_3190_7;

Selector_2 s3190_7(wires_797_6[2], addr_797_6, addr_positional[12763:12760], addr_3190_7);

wire[31:0] addr_3191_7;

Selector_2 s3191_7(wires_797_6[3], addr_797_6, addr_positional[12767:12764], addr_3191_7);

wire[31:0] addr_3192_7;

Selector_2 s3192_7(wires_798_6[0], addr_798_6, addr_positional[12771:12768], addr_3192_7);

wire[31:0] addr_3193_7;

Selector_2 s3193_7(wires_798_6[1], addr_798_6, addr_positional[12775:12772], addr_3193_7);

wire[31:0] addr_3194_7;

Selector_2 s3194_7(wires_798_6[2], addr_798_6, addr_positional[12779:12776], addr_3194_7);

wire[31:0] addr_3195_7;

Selector_2 s3195_7(wires_798_6[3], addr_798_6, addr_positional[12783:12780], addr_3195_7);

wire[31:0] addr_3196_7;

Selector_2 s3196_7(wires_799_6[0], addr_799_6, addr_positional[12787:12784], addr_3196_7);

wire[31:0] addr_3197_7;

Selector_2 s3197_7(wires_799_6[1], addr_799_6, addr_positional[12791:12788], addr_3197_7);

wire[31:0] addr_3198_7;

Selector_2 s3198_7(wires_799_6[2], addr_799_6, addr_positional[12795:12792], addr_3198_7);

wire[31:0] addr_3199_7;

Selector_2 s3199_7(wires_799_6[3], addr_799_6, addr_positional[12799:12796], addr_3199_7);

wire[31:0] addr_3200_7;

Selector_2 s3200_7(wires_800_6[0], addr_800_6, addr_positional[12803:12800], addr_3200_7);

wire[31:0] addr_3201_7;

Selector_2 s3201_7(wires_800_6[1], addr_800_6, addr_positional[12807:12804], addr_3201_7);

wire[31:0] addr_3202_7;

Selector_2 s3202_7(wires_800_6[2], addr_800_6, addr_positional[12811:12808], addr_3202_7);

wire[31:0] addr_3203_7;

Selector_2 s3203_7(wires_800_6[3], addr_800_6, addr_positional[12815:12812], addr_3203_7);

wire[31:0] addr_3204_7;

Selector_2 s3204_7(wires_801_6[0], addr_801_6, addr_positional[12819:12816], addr_3204_7);

wire[31:0] addr_3205_7;

Selector_2 s3205_7(wires_801_6[1], addr_801_6, addr_positional[12823:12820], addr_3205_7);

wire[31:0] addr_3206_7;

Selector_2 s3206_7(wires_801_6[2], addr_801_6, addr_positional[12827:12824], addr_3206_7);

wire[31:0] addr_3207_7;

Selector_2 s3207_7(wires_801_6[3], addr_801_6, addr_positional[12831:12828], addr_3207_7);

wire[31:0] addr_3208_7;

Selector_2 s3208_7(wires_802_6[0], addr_802_6, addr_positional[12835:12832], addr_3208_7);

wire[31:0] addr_3209_7;

Selector_2 s3209_7(wires_802_6[1], addr_802_6, addr_positional[12839:12836], addr_3209_7);

wire[31:0] addr_3210_7;

Selector_2 s3210_7(wires_802_6[2], addr_802_6, addr_positional[12843:12840], addr_3210_7);

wire[31:0] addr_3211_7;

Selector_2 s3211_7(wires_802_6[3], addr_802_6, addr_positional[12847:12844], addr_3211_7);

wire[31:0] addr_3212_7;

Selector_2 s3212_7(wires_803_6[0], addr_803_6, addr_positional[12851:12848], addr_3212_7);

wire[31:0] addr_3213_7;

Selector_2 s3213_7(wires_803_6[1], addr_803_6, addr_positional[12855:12852], addr_3213_7);

wire[31:0] addr_3214_7;

Selector_2 s3214_7(wires_803_6[2], addr_803_6, addr_positional[12859:12856], addr_3214_7);

wire[31:0] addr_3215_7;

Selector_2 s3215_7(wires_803_6[3], addr_803_6, addr_positional[12863:12860], addr_3215_7);

wire[31:0] addr_3216_7;

Selector_2 s3216_7(wires_804_6[0], addr_804_6, addr_positional[12867:12864], addr_3216_7);

wire[31:0] addr_3217_7;

Selector_2 s3217_7(wires_804_6[1], addr_804_6, addr_positional[12871:12868], addr_3217_7);

wire[31:0] addr_3218_7;

Selector_2 s3218_7(wires_804_6[2], addr_804_6, addr_positional[12875:12872], addr_3218_7);

wire[31:0] addr_3219_7;

Selector_2 s3219_7(wires_804_6[3], addr_804_6, addr_positional[12879:12876], addr_3219_7);

wire[31:0] addr_3220_7;

Selector_2 s3220_7(wires_805_6[0], addr_805_6, addr_positional[12883:12880], addr_3220_7);

wire[31:0] addr_3221_7;

Selector_2 s3221_7(wires_805_6[1], addr_805_6, addr_positional[12887:12884], addr_3221_7);

wire[31:0] addr_3222_7;

Selector_2 s3222_7(wires_805_6[2], addr_805_6, addr_positional[12891:12888], addr_3222_7);

wire[31:0] addr_3223_7;

Selector_2 s3223_7(wires_805_6[3], addr_805_6, addr_positional[12895:12892], addr_3223_7);

wire[31:0] addr_3224_7;

Selector_2 s3224_7(wires_806_6[0], addr_806_6, addr_positional[12899:12896], addr_3224_7);

wire[31:0] addr_3225_7;

Selector_2 s3225_7(wires_806_6[1], addr_806_6, addr_positional[12903:12900], addr_3225_7);

wire[31:0] addr_3226_7;

Selector_2 s3226_7(wires_806_6[2], addr_806_6, addr_positional[12907:12904], addr_3226_7);

wire[31:0] addr_3227_7;

Selector_2 s3227_7(wires_806_6[3], addr_806_6, addr_positional[12911:12908], addr_3227_7);

wire[31:0] addr_3228_7;

Selector_2 s3228_7(wires_807_6[0], addr_807_6, addr_positional[12915:12912], addr_3228_7);

wire[31:0] addr_3229_7;

Selector_2 s3229_7(wires_807_6[1], addr_807_6, addr_positional[12919:12916], addr_3229_7);

wire[31:0] addr_3230_7;

Selector_2 s3230_7(wires_807_6[2], addr_807_6, addr_positional[12923:12920], addr_3230_7);

wire[31:0] addr_3231_7;

Selector_2 s3231_7(wires_807_6[3], addr_807_6, addr_positional[12927:12924], addr_3231_7);

wire[31:0] addr_3232_7;

Selector_2 s3232_7(wires_808_6[0], addr_808_6, addr_positional[12931:12928], addr_3232_7);

wire[31:0] addr_3233_7;

Selector_2 s3233_7(wires_808_6[1], addr_808_6, addr_positional[12935:12932], addr_3233_7);

wire[31:0] addr_3234_7;

Selector_2 s3234_7(wires_808_6[2], addr_808_6, addr_positional[12939:12936], addr_3234_7);

wire[31:0] addr_3235_7;

Selector_2 s3235_7(wires_808_6[3], addr_808_6, addr_positional[12943:12940], addr_3235_7);

wire[31:0] addr_3236_7;

Selector_2 s3236_7(wires_809_6[0], addr_809_6, addr_positional[12947:12944], addr_3236_7);

wire[31:0] addr_3237_7;

Selector_2 s3237_7(wires_809_6[1], addr_809_6, addr_positional[12951:12948], addr_3237_7);

wire[31:0] addr_3238_7;

Selector_2 s3238_7(wires_809_6[2], addr_809_6, addr_positional[12955:12952], addr_3238_7);

wire[31:0] addr_3239_7;

Selector_2 s3239_7(wires_809_6[3], addr_809_6, addr_positional[12959:12956], addr_3239_7);

wire[31:0] addr_3240_7;

Selector_2 s3240_7(wires_810_6[0], addr_810_6, addr_positional[12963:12960], addr_3240_7);

wire[31:0] addr_3241_7;

Selector_2 s3241_7(wires_810_6[1], addr_810_6, addr_positional[12967:12964], addr_3241_7);

wire[31:0] addr_3242_7;

Selector_2 s3242_7(wires_810_6[2], addr_810_6, addr_positional[12971:12968], addr_3242_7);

wire[31:0] addr_3243_7;

Selector_2 s3243_7(wires_810_6[3], addr_810_6, addr_positional[12975:12972], addr_3243_7);

wire[31:0] addr_3244_7;

Selector_2 s3244_7(wires_811_6[0], addr_811_6, addr_positional[12979:12976], addr_3244_7);

wire[31:0] addr_3245_7;

Selector_2 s3245_7(wires_811_6[1], addr_811_6, addr_positional[12983:12980], addr_3245_7);

wire[31:0] addr_3246_7;

Selector_2 s3246_7(wires_811_6[2], addr_811_6, addr_positional[12987:12984], addr_3246_7);

wire[31:0] addr_3247_7;

Selector_2 s3247_7(wires_811_6[3], addr_811_6, addr_positional[12991:12988], addr_3247_7);

wire[31:0] addr_3248_7;

Selector_2 s3248_7(wires_812_6[0], addr_812_6, addr_positional[12995:12992], addr_3248_7);

wire[31:0] addr_3249_7;

Selector_2 s3249_7(wires_812_6[1], addr_812_6, addr_positional[12999:12996], addr_3249_7);

wire[31:0] addr_3250_7;

Selector_2 s3250_7(wires_812_6[2], addr_812_6, addr_positional[13003:13000], addr_3250_7);

wire[31:0] addr_3251_7;

Selector_2 s3251_7(wires_812_6[3], addr_812_6, addr_positional[13007:13004], addr_3251_7);

wire[31:0] addr_3252_7;

Selector_2 s3252_7(wires_813_6[0], addr_813_6, addr_positional[13011:13008], addr_3252_7);

wire[31:0] addr_3253_7;

Selector_2 s3253_7(wires_813_6[1], addr_813_6, addr_positional[13015:13012], addr_3253_7);

wire[31:0] addr_3254_7;

Selector_2 s3254_7(wires_813_6[2], addr_813_6, addr_positional[13019:13016], addr_3254_7);

wire[31:0] addr_3255_7;

Selector_2 s3255_7(wires_813_6[3], addr_813_6, addr_positional[13023:13020], addr_3255_7);

wire[31:0] addr_3256_7;

Selector_2 s3256_7(wires_814_6[0], addr_814_6, addr_positional[13027:13024], addr_3256_7);

wire[31:0] addr_3257_7;

Selector_2 s3257_7(wires_814_6[1], addr_814_6, addr_positional[13031:13028], addr_3257_7);

wire[31:0] addr_3258_7;

Selector_2 s3258_7(wires_814_6[2], addr_814_6, addr_positional[13035:13032], addr_3258_7);

wire[31:0] addr_3259_7;

Selector_2 s3259_7(wires_814_6[3], addr_814_6, addr_positional[13039:13036], addr_3259_7);

wire[31:0] addr_3260_7;

Selector_2 s3260_7(wires_815_6[0], addr_815_6, addr_positional[13043:13040], addr_3260_7);

wire[31:0] addr_3261_7;

Selector_2 s3261_7(wires_815_6[1], addr_815_6, addr_positional[13047:13044], addr_3261_7);

wire[31:0] addr_3262_7;

Selector_2 s3262_7(wires_815_6[2], addr_815_6, addr_positional[13051:13048], addr_3262_7);

wire[31:0] addr_3263_7;

Selector_2 s3263_7(wires_815_6[3], addr_815_6, addr_positional[13055:13052], addr_3263_7);

wire[31:0] addr_3264_7;

Selector_2 s3264_7(wires_816_6[0], addr_816_6, addr_positional[13059:13056], addr_3264_7);

wire[31:0] addr_3265_7;

Selector_2 s3265_7(wires_816_6[1], addr_816_6, addr_positional[13063:13060], addr_3265_7);

wire[31:0] addr_3266_7;

Selector_2 s3266_7(wires_816_6[2], addr_816_6, addr_positional[13067:13064], addr_3266_7);

wire[31:0] addr_3267_7;

Selector_2 s3267_7(wires_816_6[3], addr_816_6, addr_positional[13071:13068], addr_3267_7);

wire[31:0] addr_3268_7;

Selector_2 s3268_7(wires_817_6[0], addr_817_6, addr_positional[13075:13072], addr_3268_7);

wire[31:0] addr_3269_7;

Selector_2 s3269_7(wires_817_6[1], addr_817_6, addr_positional[13079:13076], addr_3269_7);

wire[31:0] addr_3270_7;

Selector_2 s3270_7(wires_817_6[2], addr_817_6, addr_positional[13083:13080], addr_3270_7);

wire[31:0] addr_3271_7;

Selector_2 s3271_7(wires_817_6[3], addr_817_6, addr_positional[13087:13084], addr_3271_7);

wire[31:0] addr_3272_7;

Selector_2 s3272_7(wires_818_6[0], addr_818_6, addr_positional[13091:13088], addr_3272_7);

wire[31:0] addr_3273_7;

Selector_2 s3273_7(wires_818_6[1], addr_818_6, addr_positional[13095:13092], addr_3273_7);

wire[31:0] addr_3274_7;

Selector_2 s3274_7(wires_818_6[2], addr_818_6, addr_positional[13099:13096], addr_3274_7);

wire[31:0] addr_3275_7;

Selector_2 s3275_7(wires_818_6[3], addr_818_6, addr_positional[13103:13100], addr_3275_7);

wire[31:0] addr_3276_7;

Selector_2 s3276_7(wires_819_6[0], addr_819_6, addr_positional[13107:13104], addr_3276_7);

wire[31:0] addr_3277_7;

Selector_2 s3277_7(wires_819_6[1], addr_819_6, addr_positional[13111:13108], addr_3277_7);

wire[31:0] addr_3278_7;

Selector_2 s3278_7(wires_819_6[2], addr_819_6, addr_positional[13115:13112], addr_3278_7);

wire[31:0] addr_3279_7;

Selector_2 s3279_7(wires_819_6[3], addr_819_6, addr_positional[13119:13116], addr_3279_7);

wire[31:0] addr_3280_7;

Selector_2 s3280_7(wires_820_6[0], addr_820_6, addr_positional[13123:13120], addr_3280_7);

wire[31:0] addr_3281_7;

Selector_2 s3281_7(wires_820_6[1], addr_820_6, addr_positional[13127:13124], addr_3281_7);

wire[31:0] addr_3282_7;

Selector_2 s3282_7(wires_820_6[2], addr_820_6, addr_positional[13131:13128], addr_3282_7);

wire[31:0] addr_3283_7;

Selector_2 s3283_7(wires_820_6[3], addr_820_6, addr_positional[13135:13132], addr_3283_7);

wire[31:0] addr_3284_7;

Selector_2 s3284_7(wires_821_6[0], addr_821_6, addr_positional[13139:13136], addr_3284_7);

wire[31:0] addr_3285_7;

Selector_2 s3285_7(wires_821_6[1], addr_821_6, addr_positional[13143:13140], addr_3285_7);

wire[31:0] addr_3286_7;

Selector_2 s3286_7(wires_821_6[2], addr_821_6, addr_positional[13147:13144], addr_3286_7);

wire[31:0] addr_3287_7;

Selector_2 s3287_7(wires_821_6[3], addr_821_6, addr_positional[13151:13148], addr_3287_7);

wire[31:0] addr_3288_7;

Selector_2 s3288_7(wires_822_6[0], addr_822_6, addr_positional[13155:13152], addr_3288_7);

wire[31:0] addr_3289_7;

Selector_2 s3289_7(wires_822_6[1], addr_822_6, addr_positional[13159:13156], addr_3289_7);

wire[31:0] addr_3290_7;

Selector_2 s3290_7(wires_822_6[2], addr_822_6, addr_positional[13163:13160], addr_3290_7);

wire[31:0] addr_3291_7;

Selector_2 s3291_7(wires_822_6[3], addr_822_6, addr_positional[13167:13164], addr_3291_7);

wire[31:0] addr_3292_7;

Selector_2 s3292_7(wires_823_6[0], addr_823_6, addr_positional[13171:13168], addr_3292_7);

wire[31:0] addr_3293_7;

Selector_2 s3293_7(wires_823_6[1], addr_823_6, addr_positional[13175:13172], addr_3293_7);

wire[31:0] addr_3294_7;

Selector_2 s3294_7(wires_823_6[2], addr_823_6, addr_positional[13179:13176], addr_3294_7);

wire[31:0] addr_3295_7;

Selector_2 s3295_7(wires_823_6[3], addr_823_6, addr_positional[13183:13180], addr_3295_7);

wire[31:0] addr_3296_7;

Selector_2 s3296_7(wires_824_6[0], addr_824_6, addr_positional[13187:13184], addr_3296_7);

wire[31:0] addr_3297_7;

Selector_2 s3297_7(wires_824_6[1], addr_824_6, addr_positional[13191:13188], addr_3297_7);

wire[31:0] addr_3298_7;

Selector_2 s3298_7(wires_824_6[2], addr_824_6, addr_positional[13195:13192], addr_3298_7);

wire[31:0] addr_3299_7;

Selector_2 s3299_7(wires_824_6[3], addr_824_6, addr_positional[13199:13196], addr_3299_7);

wire[31:0] addr_3300_7;

Selector_2 s3300_7(wires_825_6[0], addr_825_6, addr_positional[13203:13200], addr_3300_7);

wire[31:0] addr_3301_7;

Selector_2 s3301_7(wires_825_6[1], addr_825_6, addr_positional[13207:13204], addr_3301_7);

wire[31:0] addr_3302_7;

Selector_2 s3302_7(wires_825_6[2], addr_825_6, addr_positional[13211:13208], addr_3302_7);

wire[31:0] addr_3303_7;

Selector_2 s3303_7(wires_825_6[3], addr_825_6, addr_positional[13215:13212], addr_3303_7);

wire[31:0] addr_3304_7;

Selector_2 s3304_7(wires_826_6[0], addr_826_6, addr_positional[13219:13216], addr_3304_7);

wire[31:0] addr_3305_7;

Selector_2 s3305_7(wires_826_6[1], addr_826_6, addr_positional[13223:13220], addr_3305_7);

wire[31:0] addr_3306_7;

Selector_2 s3306_7(wires_826_6[2], addr_826_6, addr_positional[13227:13224], addr_3306_7);

wire[31:0] addr_3307_7;

Selector_2 s3307_7(wires_826_6[3], addr_826_6, addr_positional[13231:13228], addr_3307_7);

wire[31:0] addr_3308_7;

Selector_2 s3308_7(wires_827_6[0], addr_827_6, addr_positional[13235:13232], addr_3308_7);

wire[31:0] addr_3309_7;

Selector_2 s3309_7(wires_827_6[1], addr_827_6, addr_positional[13239:13236], addr_3309_7);

wire[31:0] addr_3310_7;

Selector_2 s3310_7(wires_827_6[2], addr_827_6, addr_positional[13243:13240], addr_3310_7);

wire[31:0] addr_3311_7;

Selector_2 s3311_7(wires_827_6[3], addr_827_6, addr_positional[13247:13244], addr_3311_7);

wire[31:0] addr_3312_7;

Selector_2 s3312_7(wires_828_6[0], addr_828_6, addr_positional[13251:13248], addr_3312_7);

wire[31:0] addr_3313_7;

Selector_2 s3313_7(wires_828_6[1], addr_828_6, addr_positional[13255:13252], addr_3313_7);

wire[31:0] addr_3314_7;

Selector_2 s3314_7(wires_828_6[2], addr_828_6, addr_positional[13259:13256], addr_3314_7);

wire[31:0] addr_3315_7;

Selector_2 s3315_7(wires_828_6[3], addr_828_6, addr_positional[13263:13260], addr_3315_7);

wire[31:0] addr_3316_7;

Selector_2 s3316_7(wires_829_6[0], addr_829_6, addr_positional[13267:13264], addr_3316_7);

wire[31:0] addr_3317_7;

Selector_2 s3317_7(wires_829_6[1], addr_829_6, addr_positional[13271:13268], addr_3317_7);

wire[31:0] addr_3318_7;

Selector_2 s3318_7(wires_829_6[2], addr_829_6, addr_positional[13275:13272], addr_3318_7);

wire[31:0] addr_3319_7;

Selector_2 s3319_7(wires_829_6[3], addr_829_6, addr_positional[13279:13276], addr_3319_7);

wire[31:0] addr_3320_7;

Selector_2 s3320_7(wires_830_6[0], addr_830_6, addr_positional[13283:13280], addr_3320_7);

wire[31:0] addr_3321_7;

Selector_2 s3321_7(wires_830_6[1], addr_830_6, addr_positional[13287:13284], addr_3321_7);

wire[31:0] addr_3322_7;

Selector_2 s3322_7(wires_830_6[2], addr_830_6, addr_positional[13291:13288], addr_3322_7);

wire[31:0] addr_3323_7;

Selector_2 s3323_7(wires_830_6[3], addr_830_6, addr_positional[13295:13292], addr_3323_7);

wire[31:0] addr_3324_7;

Selector_2 s3324_7(wires_831_6[0], addr_831_6, addr_positional[13299:13296], addr_3324_7);

wire[31:0] addr_3325_7;

Selector_2 s3325_7(wires_831_6[1], addr_831_6, addr_positional[13303:13300], addr_3325_7);

wire[31:0] addr_3326_7;

Selector_2 s3326_7(wires_831_6[2], addr_831_6, addr_positional[13307:13304], addr_3326_7);

wire[31:0] addr_3327_7;

Selector_2 s3327_7(wires_831_6[3], addr_831_6, addr_positional[13311:13308], addr_3327_7);

wire[31:0] addr_3328_7;

Selector_2 s3328_7(wires_832_6[0], addr_832_6, addr_positional[13315:13312], addr_3328_7);

wire[31:0] addr_3329_7;

Selector_2 s3329_7(wires_832_6[1], addr_832_6, addr_positional[13319:13316], addr_3329_7);

wire[31:0] addr_3330_7;

Selector_2 s3330_7(wires_832_6[2], addr_832_6, addr_positional[13323:13320], addr_3330_7);

wire[31:0] addr_3331_7;

Selector_2 s3331_7(wires_832_6[3], addr_832_6, addr_positional[13327:13324], addr_3331_7);

wire[31:0] addr_3332_7;

Selector_2 s3332_7(wires_833_6[0], addr_833_6, addr_positional[13331:13328], addr_3332_7);

wire[31:0] addr_3333_7;

Selector_2 s3333_7(wires_833_6[1], addr_833_6, addr_positional[13335:13332], addr_3333_7);

wire[31:0] addr_3334_7;

Selector_2 s3334_7(wires_833_6[2], addr_833_6, addr_positional[13339:13336], addr_3334_7);

wire[31:0] addr_3335_7;

Selector_2 s3335_7(wires_833_6[3], addr_833_6, addr_positional[13343:13340], addr_3335_7);

wire[31:0] addr_3336_7;

Selector_2 s3336_7(wires_834_6[0], addr_834_6, addr_positional[13347:13344], addr_3336_7);

wire[31:0] addr_3337_7;

Selector_2 s3337_7(wires_834_6[1], addr_834_6, addr_positional[13351:13348], addr_3337_7);

wire[31:0] addr_3338_7;

Selector_2 s3338_7(wires_834_6[2], addr_834_6, addr_positional[13355:13352], addr_3338_7);

wire[31:0] addr_3339_7;

Selector_2 s3339_7(wires_834_6[3], addr_834_6, addr_positional[13359:13356], addr_3339_7);

wire[31:0] addr_3340_7;

Selector_2 s3340_7(wires_835_6[0], addr_835_6, addr_positional[13363:13360], addr_3340_7);

wire[31:0] addr_3341_7;

Selector_2 s3341_7(wires_835_6[1], addr_835_6, addr_positional[13367:13364], addr_3341_7);

wire[31:0] addr_3342_7;

Selector_2 s3342_7(wires_835_6[2], addr_835_6, addr_positional[13371:13368], addr_3342_7);

wire[31:0] addr_3343_7;

Selector_2 s3343_7(wires_835_6[3], addr_835_6, addr_positional[13375:13372], addr_3343_7);

wire[31:0] addr_3344_7;

Selector_2 s3344_7(wires_836_6[0], addr_836_6, addr_positional[13379:13376], addr_3344_7);

wire[31:0] addr_3345_7;

Selector_2 s3345_7(wires_836_6[1], addr_836_6, addr_positional[13383:13380], addr_3345_7);

wire[31:0] addr_3346_7;

Selector_2 s3346_7(wires_836_6[2], addr_836_6, addr_positional[13387:13384], addr_3346_7);

wire[31:0] addr_3347_7;

Selector_2 s3347_7(wires_836_6[3], addr_836_6, addr_positional[13391:13388], addr_3347_7);

wire[31:0] addr_3348_7;

Selector_2 s3348_7(wires_837_6[0], addr_837_6, addr_positional[13395:13392], addr_3348_7);

wire[31:0] addr_3349_7;

Selector_2 s3349_7(wires_837_6[1], addr_837_6, addr_positional[13399:13396], addr_3349_7);

wire[31:0] addr_3350_7;

Selector_2 s3350_7(wires_837_6[2], addr_837_6, addr_positional[13403:13400], addr_3350_7);

wire[31:0] addr_3351_7;

Selector_2 s3351_7(wires_837_6[3], addr_837_6, addr_positional[13407:13404], addr_3351_7);

wire[31:0] addr_3352_7;

Selector_2 s3352_7(wires_838_6[0], addr_838_6, addr_positional[13411:13408], addr_3352_7);

wire[31:0] addr_3353_7;

Selector_2 s3353_7(wires_838_6[1], addr_838_6, addr_positional[13415:13412], addr_3353_7);

wire[31:0] addr_3354_7;

Selector_2 s3354_7(wires_838_6[2], addr_838_6, addr_positional[13419:13416], addr_3354_7);

wire[31:0] addr_3355_7;

Selector_2 s3355_7(wires_838_6[3], addr_838_6, addr_positional[13423:13420], addr_3355_7);

wire[31:0] addr_3356_7;

Selector_2 s3356_7(wires_839_6[0], addr_839_6, addr_positional[13427:13424], addr_3356_7);

wire[31:0] addr_3357_7;

Selector_2 s3357_7(wires_839_6[1], addr_839_6, addr_positional[13431:13428], addr_3357_7);

wire[31:0] addr_3358_7;

Selector_2 s3358_7(wires_839_6[2], addr_839_6, addr_positional[13435:13432], addr_3358_7);

wire[31:0] addr_3359_7;

Selector_2 s3359_7(wires_839_6[3], addr_839_6, addr_positional[13439:13436], addr_3359_7);

wire[31:0] addr_3360_7;

Selector_2 s3360_7(wires_840_6[0], addr_840_6, addr_positional[13443:13440], addr_3360_7);

wire[31:0] addr_3361_7;

Selector_2 s3361_7(wires_840_6[1], addr_840_6, addr_positional[13447:13444], addr_3361_7);

wire[31:0] addr_3362_7;

Selector_2 s3362_7(wires_840_6[2], addr_840_6, addr_positional[13451:13448], addr_3362_7);

wire[31:0] addr_3363_7;

Selector_2 s3363_7(wires_840_6[3], addr_840_6, addr_positional[13455:13452], addr_3363_7);

wire[31:0] addr_3364_7;

Selector_2 s3364_7(wires_841_6[0], addr_841_6, addr_positional[13459:13456], addr_3364_7);

wire[31:0] addr_3365_7;

Selector_2 s3365_7(wires_841_6[1], addr_841_6, addr_positional[13463:13460], addr_3365_7);

wire[31:0] addr_3366_7;

Selector_2 s3366_7(wires_841_6[2], addr_841_6, addr_positional[13467:13464], addr_3366_7);

wire[31:0] addr_3367_7;

Selector_2 s3367_7(wires_841_6[3], addr_841_6, addr_positional[13471:13468], addr_3367_7);

wire[31:0] addr_3368_7;

Selector_2 s3368_7(wires_842_6[0], addr_842_6, addr_positional[13475:13472], addr_3368_7);

wire[31:0] addr_3369_7;

Selector_2 s3369_7(wires_842_6[1], addr_842_6, addr_positional[13479:13476], addr_3369_7);

wire[31:0] addr_3370_7;

Selector_2 s3370_7(wires_842_6[2], addr_842_6, addr_positional[13483:13480], addr_3370_7);

wire[31:0] addr_3371_7;

Selector_2 s3371_7(wires_842_6[3], addr_842_6, addr_positional[13487:13484], addr_3371_7);

wire[31:0] addr_3372_7;

Selector_2 s3372_7(wires_843_6[0], addr_843_6, addr_positional[13491:13488], addr_3372_7);

wire[31:0] addr_3373_7;

Selector_2 s3373_7(wires_843_6[1], addr_843_6, addr_positional[13495:13492], addr_3373_7);

wire[31:0] addr_3374_7;

Selector_2 s3374_7(wires_843_6[2], addr_843_6, addr_positional[13499:13496], addr_3374_7);

wire[31:0] addr_3375_7;

Selector_2 s3375_7(wires_843_6[3], addr_843_6, addr_positional[13503:13500], addr_3375_7);

wire[31:0] addr_3376_7;

Selector_2 s3376_7(wires_844_6[0], addr_844_6, addr_positional[13507:13504], addr_3376_7);

wire[31:0] addr_3377_7;

Selector_2 s3377_7(wires_844_6[1], addr_844_6, addr_positional[13511:13508], addr_3377_7);

wire[31:0] addr_3378_7;

Selector_2 s3378_7(wires_844_6[2], addr_844_6, addr_positional[13515:13512], addr_3378_7);

wire[31:0] addr_3379_7;

Selector_2 s3379_7(wires_844_6[3], addr_844_6, addr_positional[13519:13516], addr_3379_7);

wire[31:0] addr_3380_7;

Selector_2 s3380_7(wires_845_6[0], addr_845_6, addr_positional[13523:13520], addr_3380_7);

wire[31:0] addr_3381_7;

Selector_2 s3381_7(wires_845_6[1], addr_845_6, addr_positional[13527:13524], addr_3381_7);

wire[31:0] addr_3382_7;

Selector_2 s3382_7(wires_845_6[2], addr_845_6, addr_positional[13531:13528], addr_3382_7);

wire[31:0] addr_3383_7;

Selector_2 s3383_7(wires_845_6[3], addr_845_6, addr_positional[13535:13532], addr_3383_7);

wire[31:0] addr_3384_7;

Selector_2 s3384_7(wires_846_6[0], addr_846_6, addr_positional[13539:13536], addr_3384_7);

wire[31:0] addr_3385_7;

Selector_2 s3385_7(wires_846_6[1], addr_846_6, addr_positional[13543:13540], addr_3385_7);

wire[31:0] addr_3386_7;

Selector_2 s3386_7(wires_846_6[2], addr_846_6, addr_positional[13547:13544], addr_3386_7);

wire[31:0] addr_3387_7;

Selector_2 s3387_7(wires_846_6[3], addr_846_6, addr_positional[13551:13548], addr_3387_7);

wire[31:0] addr_3388_7;

Selector_2 s3388_7(wires_847_6[0], addr_847_6, addr_positional[13555:13552], addr_3388_7);

wire[31:0] addr_3389_7;

Selector_2 s3389_7(wires_847_6[1], addr_847_6, addr_positional[13559:13556], addr_3389_7);

wire[31:0] addr_3390_7;

Selector_2 s3390_7(wires_847_6[2], addr_847_6, addr_positional[13563:13560], addr_3390_7);

wire[31:0] addr_3391_7;

Selector_2 s3391_7(wires_847_6[3], addr_847_6, addr_positional[13567:13564], addr_3391_7);

wire[31:0] addr_3392_7;

Selector_2 s3392_7(wires_848_6[0], addr_848_6, addr_positional[13571:13568], addr_3392_7);

wire[31:0] addr_3393_7;

Selector_2 s3393_7(wires_848_6[1], addr_848_6, addr_positional[13575:13572], addr_3393_7);

wire[31:0] addr_3394_7;

Selector_2 s3394_7(wires_848_6[2], addr_848_6, addr_positional[13579:13576], addr_3394_7);

wire[31:0] addr_3395_7;

Selector_2 s3395_7(wires_848_6[3], addr_848_6, addr_positional[13583:13580], addr_3395_7);

wire[31:0] addr_3396_7;

Selector_2 s3396_7(wires_849_6[0], addr_849_6, addr_positional[13587:13584], addr_3396_7);

wire[31:0] addr_3397_7;

Selector_2 s3397_7(wires_849_6[1], addr_849_6, addr_positional[13591:13588], addr_3397_7);

wire[31:0] addr_3398_7;

Selector_2 s3398_7(wires_849_6[2], addr_849_6, addr_positional[13595:13592], addr_3398_7);

wire[31:0] addr_3399_7;

Selector_2 s3399_7(wires_849_6[3], addr_849_6, addr_positional[13599:13596], addr_3399_7);

wire[31:0] addr_3400_7;

Selector_2 s3400_7(wires_850_6[0], addr_850_6, addr_positional[13603:13600], addr_3400_7);

wire[31:0] addr_3401_7;

Selector_2 s3401_7(wires_850_6[1], addr_850_6, addr_positional[13607:13604], addr_3401_7);

wire[31:0] addr_3402_7;

Selector_2 s3402_7(wires_850_6[2], addr_850_6, addr_positional[13611:13608], addr_3402_7);

wire[31:0] addr_3403_7;

Selector_2 s3403_7(wires_850_6[3], addr_850_6, addr_positional[13615:13612], addr_3403_7);

wire[31:0] addr_3404_7;

Selector_2 s3404_7(wires_851_6[0], addr_851_6, addr_positional[13619:13616], addr_3404_7);

wire[31:0] addr_3405_7;

Selector_2 s3405_7(wires_851_6[1], addr_851_6, addr_positional[13623:13620], addr_3405_7);

wire[31:0] addr_3406_7;

Selector_2 s3406_7(wires_851_6[2], addr_851_6, addr_positional[13627:13624], addr_3406_7);

wire[31:0] addr_3407_7;

Selector_2 s3407_7(wires_851_6[3], addr_851_6, addr_positional[13631:13628], addr_3407_7);

wire[31:0] addr_3408_7;

Selector_2 s3408_7(wires_852_6[0], addr_852_6, addr_positional[13635:13632], addr_3408_7);

wire[31:0] addr_3409_7;

Selector_2 s3409_7(wires_852_6[1], addr_852_6, addr_positional[13639:13636], addr_3409_7);

wire[31:0] addr_3410_7;

Selector_2 s3410_7(wires_852_6[2], addr_852_6, addr_positional[13643:13640], addr_3410_7);

wire[31:0] addr_3411_7;

Selector_2 s3411_7(wires_852_6[3], addr_852_6, addr_positional[13647:13644], addr_3411_7);

wire[31:0] addr_3412_7;

Selector_2 s3412_7(wires_853_6[0], addr_853_6, addr_positional[13651:13648], addr_3412_7);

wire[31:0] addr_3413_7;

Selector_2 s3413_7(wires_853_6[1], addr_853_6, addr_positional[13655:13652], addr_3413_7);

wire[31:0] addr_3414_7;

Selector_2 s3414_7(wires_853_6[2], addr_853_6, addr_positional[13659:13656], addr_3414_7);

wire[31:0] addr_3415_7;

Selector_2 s3415_7(wires_853_6[3], addr_853_6, addr_positional[13663:13660], addr_3415_7);

wire[31:0] addr_3416_7;

Selector_2 s3416_7(wires_854_6[0], addr_854_6, addr_positional[13667:13664], addr_3416_7);

wire[31:0] addr_3417_7;

Selector_2 s3417_7(wires_854_6[1], addr_854_6, addr_positional[13671:13668], addr_3417_7);

wire[31:0] addr_3418_7;

Selector_2 s3418_7(wires_854_6[2], addr_854_6, addr_positional[13675:13672], addr_3418_7);

wire[31:0] addr_3419_7;

Selector_2 s3419_7(wires_854_6[3], addr_854_6, addr_positional[13679:13676], addr_3419_7);

wire[31:0] addr_3420_7;

Selector_2 s3420_7(wires_855_6[0], addr_855_6, addr_positional[13683:13680], addr_3420_7);

wire[31:0] addr_3421_7;

Selector_2 s3421_7(wires_855_6[1], addr_855_6, addr_positional[13687:13684], addr_3421_7);

wire[31:0] addr_3422_7;

Selector_2 s3422_7(wires_855_6[2], addr_855_6, addr_positional[13691:13688], addr_3422_7);

wire[31:0] addr_3423_7;

Selector_2 s3423_7(wires_855_6[3], addr_855_6, addr_positional[13695:13692], addr_3423_7);

wire[31:0] addr_3424_7;

Selector_2 s3424_7(wires_856_6[0], addr_856_6, addr_positional[13699:13696], addr_3424_7);

wire[31:0] addr_3425_7;

Selector_2 s3425_7(wires_856_6[1], addr_856_6, addr_positional[13703:13700], addr_3425_7);

wire[31:0] addr_3426_7;

Selector_2 s3426_7(wires_856_6[2], addr_856_6, addr_positional[13707:13704], addr_3426_7);

wire[31:0] addr_3427_7;

Selector_2 s3427_7(wires_856_6[3], addr_856_6, addr_positional[13711:13708], addr_3427_7);

wire[31:0] addr_3428_7;

Selector_2 s3428_7(wires_857_6[0], addr_857_6, addr_positional[13715:13712], addr_3428_7);

wire[31:0] addr_3429_7;

Selector_2 s3429_7(wires_857_6[1], addr_857_6, addr_positional[13719:13716], addr_3429_7);

wire[31:0] addr_3430_7;

Selector_2 s3430_7(wires_857_6[2], addr_857_6, addr_positional[13723:13720], addr_3430_7);

wire[31:0] addr_3431_7;

Selector_2 s3431_7(wires_857_6[3], addr_857_6, addr_positional[13727:13724], addr_3431_7);

wire[31:0] addr_3432_7;

Selector_2 s3432_7(wires_858_6[0], addr_858_6, addr_positional[13731:13728], addr_3432_7);

wire[31:0] addr_3433_7;

Selector_2 s3433_7(wires_858_6[1], addr_858_6, addr_positional[13735:13732], addr_3433_7);

wire[31:0] addr_3434_7;

Selector_2 s3434_7(wires_858_6[2], addr_858_6, addr_positional[13739:13736], addr_3434_7);

wire[31:0] addr_3435_7;

Selector_2 s3435_7(wires_858_6[3], addr_858_6, addr_positional[13743:13740], addr_3435_7);

wire[31:0] addr_3436_7;

Selector_2 s3436_7(wires_859_6[0], addr_859_6, addr_positional[13747:13744], addr_3436_7);

wire[31:0] addr_3437_7;

Selector_2 s3437_7(wires_859_6[1], addr_859_6, addr_positional[13751:13748], addr_3437_7);

wire[31:0] addr_3438_7;

Selector_2 s3438_7(wires_859_6[2], addr_859_6, addr_positional[13755:13752], addr_3438_7);

wire[31:0] addr_3439_7;

Selector_2 s3439_7(wires_859_6[3], addr_859_6, addr_positional[13759:13756], addr_3439_7);

wire[31:0] addr_3440_7;

Selector_2 s3440_7(wires_860_6[0], addr_860_6, addr_positional[13763:13760], addr_3440_7);

wire[31:0] addr_3441_7;

Selector_2 s3441_7(wires_860_6[1], addr_860_6, addr_positional[13767:13764], addr_3441_7);

wire[31:0] addr_3442_7;

Selector_2 s3442_7(wires_860_6[2], addr_860_6, addr_positional[13771:13768], addr_3442_7);

wire[31:0] addr_3443_7;

Selector_2 s3443_7(wires_860_6[3], addr_860_6, addr_positional[13775:13772], addr_3443_7);

wire[31:0] addr_3444_7;

Selector_2 s3444_7(wires_861_6[0], addr_861_6, addr_positional[13779:13776], addr_3444_7);

wire[31:0] addr_3445_7;

Selector_2 s3445_7(wires_861_6[1], addr_861_6, addr_positional[13783:13780], addr_3445_7);

wire[31:0] addr_3446_7;

Selector_2 s3446_7(wires_861_6[2], addr_861_6, addr_positional[13787:13784], addr_3446_7);

wire[31:0] addr_3447_7;

Selector_2 s3447_7(wires_861_6[3], addr_861_6, addr_positional[13791:13788], addr_3447_7);

wire[31:0] addr_3448_7;

Selector_2 s3448_7(wires_862_6[0], addr_862_6, addr_positional[13795:13792], addr_3448_7);

wire[31:0] addr_3449_7;

Selector_2 s3449_7(wires_862_6[1], addr_862_6, addr_positional[13799:13796], addr_3449_7);

wire[31:0] addr_3450_7;

Selector_2 s3450_7(wires_862_6[2], addr_862_6, addr_positional[13803:13800], addr_3450_7);

wire[31:0] addr_3451_7;

Selector_2 s3451_7(wires_862_6[3], addr_862_6, addr_positional[13807:13804], addr_3451_7);

wire[31:0] addr_3452_7;

Selector_2 s3452_7(wires_863_6[0], addr_863_6, addr_positional[13811:13808], addr_3452_7);

wire[31:0] addr_3453_7;

Selector_2 s3453_7(wires_863_6[1], addr_863_6, addr_positional[13815:13812], addr_3453_7);

wire[31:0] addr_3454_7;

Selector_2 s3454_7(wires_863_6[2], addr_863_6, addr_positional[13819:13816], addr_3454_7);

wire[31:0] addr_3455_7;

Selector_2 s3455_7(wires_863_6[3], addr_863_6, addr_positional[13823:13820], addr_3455_7);

wire[31:0] addr_3456_7;

Selector_2 s3456_7(wires_864_6[0], addr_864_6, addr_positional[13827:13824], addr_3456_7);

wire[31:0] addr_3457_7;

Selector_2 s3457_7(wires_864_6[1], addr_864_6, addr_positional[13831:13828], addr_3457_7);

wire[31:0] addr_3458_7;

Selector_2 s3458_7(wires_864_6[2], addr_864_6, addr_positional[13835:13832], addr_3458_7);

wire[31:0] addr_3459_7;

Selector_2 s3459_7(wires_864_6[3], addr_864_6, addr_positional[13839:13836], addr_3459_7);

wire[31:0] addr_3460_7;

Selector_2 s3460_7(wires_865_6[0], addr_865_6, addr_positional[13843:13840], addr_3460_7);

wire[31:0] addr_3461_7;

Selector_2 s3461_7(wires_865_6[1], addr_865_6, addr_positional[13847:13844], addr_3461_7);

wire[31:0] addr_3462_7;

Selector_2 s3462_7(wires_865_6[2], addr_865_6, addr_positional[13851:13848], addr_3462_7);

wire[31:0] addr_3463_7;

Selector_2 s3463_7(wires_865_6[3], addr_865_6, addr_positional[13855:13852], addr_3463_7);

wire[31:0] addr_3464_7;

Selector_2 s3464_7(wires_866_6[0], addr_866_6, addr_positional[13859:13856], addr_3464_7);

wire[31:0] addr_3465_7;

Selector_2 s3465_7(wires_866_6[1], addr_866_6, addr_positional[13863:13860], addr_3465_7);

wire[31:0] addr_3466_7;

Selector_2 s3466_7(wires_866_6[2], addr_866_6, addr_positional[13867:13864], addr_3466_7);

wire[31:0] addr_3467_7;

Selector_2 s3467_7(wires_866_6[3], addr_866_6, addr_positional[13871:13868], addr_3467_7);

wire[31:0] addr_3468_7;

Selector_2 s3468_7(wires_867_6[0], addr_867_6, addr_positional[13875:13872], addr_3468_7);

wire[31:0] addr_3469_7;

Selector_2 s3469_7(wires_867_6[1], addr_867_6, addr_positional[13879:13876], addr_3469_7);

wire[31:0] addr_3470_7;

Selector_2 s3470_7(wires_867_6[2], addr_867_6, addr_positional[13883:13880], addr_3470_7);

wire[31:0] addr_3471_7;

Selector_2 s3471_7(wires_867_6[3], addr_867_6, addr_positional[13887:13884], addr_3471_7);

wire[31:0] addr_3472_7;

Selector_2 s3472_7(wires_868_6[0], addr_868_6, addr_positional[13891:13888], addr_3472_7);

wire[31:0] addr_3473_7;

Selector_2 s3473_7(wires_868_6[1], addr_868_6, addr_positional[13895:13892], addr_3473_7);

wire[31:0] addr_3474_7;

Selector_2 s3474_7(wires_868_6[2], addr_868_6, addr_positional[13899:13896], addr_3474_7);

wire[31:0] addr_3475_7;

Selector_2 s3475_7(wires_868_6[3], addr_868_6, addr_positional[13903:13900], addr_3475_7);

wire[31:0] addr_3476_7;

Selector_2 s3476_7(wires_869_6[0], addr_869_6, addr_positional[13907:13904], addr_3476_7);

wire[31:0] addr_3477_7;

Selector_2 s3477_7(wires_869_6[1], addr_869_6, addr_positional[13911:13908], addr_3477_7);

wire[31:0] addr_3478_7;

Selector_2 s3478_7(wires_869_6[2], addr_869_6, addr_positional[13915:13912], addr_3478_7);

wire[31:0] addr_3479_7;

Selector_2 s3479_7(wires_869_6[3], addr_869_6, addr_positional[13919:13916], addr_3479_7);

wire[31:0] addr_3480_7;

Selector_2 s3480_7(wires_870_6[0], addr_870_6, addr_positional[13923:13920], addr_3480_7);

wire[31:0] addr_3481_7;

Selector_2 s3481_7(wires_870_6[1], addr_870_6, addr_positional[13927:13924], addr_3481_7);

wire[31:0] addr_3482_7;

Selector_2 s3482_7(wires_870_6[2], addr_870_6, addr_positional[13931:13928], addr_3482_7);

wire[31:0] addr_3483_7;

Selector_2 s3483_7(wires_870_6[3], addr_870_6, addr_positional[13935:13932], addr_3483_7);

wire[31:0] addr_3484_7;

Selector_2 s3484_7(wires_871_6[0], addr_871_6, addr_positional[13939:13936], addr_3484_7);

wire[31:0] addr_3485_7;

Selector_2 s3485_7(wires_871_6[1], addr_871_6, addr_positional[13943:13940], addr_3485_7);

wire[31:0] addr_3486_7;

Selector_2 s3486_7(wires_871_6[2], addr_871_6, addr_positional[13947:13944], addr_3486_7);

wire[31:0] addr_3487_7;

Selector_2 s3487_7(wires_871_6[3], addr_871_6, addr_positional[13951:13948], addr_3487_7);

wire[31:0] addr_3488_7;

Selector_2 s3488_7(wires_872_6[0], addr_872_6, addr_positional[13955:13952], addr_3488_7);

wire[31:0] addr_3489_7;

Selector_2 s3489_7(wires_872_6[1], addr_872_6, addr_positional[13959:13956], addr_3489_7);

wire[31:0] addr_3490_7;

Selector_2 s3490_7(wires_872_6[2], addr_872_6, addr_positional[13963:13960], addr_3490_7);

wire[31:0] addr_3491_7;

Selector_2 s3491_7(wires_872_6[3], addr_872_6, addr_positional[13967:13964], addr_3491_7);

wire[31:0] addr_3492_7;

Selector_2 s3492_7(wires_873_6[0], addr_873_6, addr_positional[13971:13968], addr_3492_7);

wire[31:0] addr_3493_7;

Selector_2 s3493_7(wires_873_6[1], addr_873_6, addr_positional[13975:13972], addr_3493_7);

wire[31:0] addr_3494_7;

Selector_2 s3494_7(wires_873_6[2], addr_873_6, addr_positional[13979:13976], addr_3494_7);

wire[31:0] addr_3495_7;

Selector_2 s3495_7(wires_873_6[3], addr_873_6, addr_positional[13983:13980], addr_3495_7);

wire[31:0] addr_3496_7;

Selector_2 s3496_7(wires_874_6[0], addr_874_6, addr_positional[13987:13984], addr_3496_7);

wire[31:0] addr_3497_7;

Selector_2 s3497_7(wires_874_6[1], addr_874_6, addr_positional[13991:13988], addr_3497_7);

wire[31:0] addr_3498_7;

Selector_2 s3498_7(wires_874_6[2], addr_874_6, addr_positional[13995:13992], addr_3498_7);

wire[31:0] addr_3499_7;

Selector_2 s3499_7(wires_874_6[3], addr_874_6, addr_positional[13999:13996], addr_3499_7);

wire[31:0] addr_3500_7;

Selector_2 s3500_7(wires_875_6[0], addr_875_6, addr_positional[14003:14000], addr_3500_7);

wire[31:0] addr_3501_7;

Selector_2 s3501_7(wires_875_6[1], addr_875_6, addr_positional[14007:14004], addr_3501_7);

wire[31:0] addr_3502_7;

Selector_2 s3502_7(wires_875_6[2], addr_875_6, addr_positional[14011:14008], addr_3502_7);

wire[31:0] addr_3503_7;

Selector_2 s3503_7(wires_875_6[3], addr_875_6, addr_positional[14015:14012], addr_3503_7);

wire[31:0] addr_3504_7;

Selector_2 s3504_7(wires_876_6[0], addr_876_6, addr_positional[14019:14016], addr_3504_7);

wire[31:0] addr_3505_7;

Selector_2 s3505_7(wires_876_6[1], addr_876_6, addr_positional[14023:14020], addr_3505_7);

wire[31:0] addr_3506_7;

Selector_2 s3506_7(wires_876_6[2], addr_876_6, addr_positional[14027:14024], addr_3506_7);

wire[31:0] addr_3507_7;

Selector_2 s3507_7(wires_876_6[3], addr_876_6, addr_positional[14031:14028], addr_3507_7);

wire[31:0] addr_3508_7;

Selector_2 s3508_7(wires_877_6[0], addr_877_6, addr_positional[14035:14032], addr_3508_7);

wire[31:0] addr_3509_7;

Selector_2 s3509_7(wires_877_6[1], addr_877_6, addr_positional[14039:14036], addr_3509_7);

wire[31:0] addr_3510_7;

Selector_2 s3510_7(wires_877_6[2], addr_877_6, addr_positional[14043:14040], addr_3510_7);

wire[31:0] addr_3511_7;

Selector_2 s3511_7(wires_877_6[3], addr_877_6, addr_positional[14047:14044], addr_3511_7);

wire[31:0] addr_3512_7;

Selector_2 s3512_7(wires_878_6[0], addr_878_6, addr_positional[14051:14048], addr_3512_7);

wire[31:0] addr_3513_7;

Selector_2 s3513_7(wires_878_6[1], addr_878_6, addr_positional[14055:14052], addr_3513_7);

wire[31:0] addr_3514_7;

Selector_2 s3514_7(wires_878_6[2], addr_878_6, addr_positional[14059:14056], addr_3514_7);

wire[31:0] addr_3515_7;

Selector_2 s3515_7(wires_878_6[3], addr_878_6, addr_positional[14063:14060], addr_3515_7);

wire[31:0] addr_3516_7;

Selector_2 s3516_7(wires_879_6[0], addr_879_6, addr_positional[14067:14064], addr_3516_7);

wire[31:0] addr_3517_7;

Selector_2 s3517_7(wires_879_6[1], addr_879_6, addr_positional[14071:14068], addr_3517_7);

wire[31:0] addr_3518_7;

Selector_2 s3518_7(wires_879_6[2], addr_879_6, addr_positional[14075:14072], addr_3518_7);

wire[31:0] addr_3519_7;

Selector_2 s3519_7(wires_879_6[3], addr_879_6, addr_positional[14079:14076], addr_3519_7);

wire[31:0] addr_3520_7;

Selector_2 s3520_7(wires_880_6[0], addr_880_6, addr_positional[14083:14080], addr_3520_7);

wire[31:0] addr_3521_7;

Selector_2 s3521_7(wires_880_6[1], addr_880_6, addr_positional[14087:14084], addr_3521_7);

wire[31:0] addr_3522_7;

Selector_2 s3522_7(wires_880_6[2], addr_880_6, addr_positional[14091:14088], addr_3522_7);

wire[31:0] addr_3523_7;

Selector_2 s3523_7(wires_880_6[3], addr_880_6, addr_positional[14095:14092], addr_3523_7);

wire[31:0] addr_3524_7;

Selector_2 s3524_7(wires_881_6[0], addr_881_6, addr_positional[14099:14096], addr_3524_7);

wire[31:0] addr_3525_7;

Selector_2 s3525_7(wires_881_6[1], addr_881_6, addr_positional[14103:14100], addr_3525_7);

wire[31:0] addr_3526_7;

Selector_2 s3526_7(wires_881_6[2], addr_881_6, addr_positional[14107:14104], addr_3526_7);

wire[31:0] addr_3527_7;

Selector_2 s3527_7(wires_881_6[3], addr_881_6, addr_positional[14111:14108], addr_3527_7);

wire[31:0] addr_3528_7;

Selector_2 s3528_7(wires_882_6[0], addr_882_6, addr_positional[14115:14112], addr_3528_7);

wire[31:0] addr_3529_7;

Selector_2 s3529_7(wires_882_6[1], addr_882_6, addr_positional[14119:14116], addr_3529_7);

wire[31:0] addr_3530_7;

Selector_2 s3530_7(wires_882_6[2], addr_882_6, addr_positional[14123:14120], addr_3530_7);

wire[31:0] addr_3531_7;

Selector_2 s3531_7(wires_882_6[3], addr_882_6, addr_positional[14127:14124], addr_3531_7);

wire[31:0] addr_3532_7;

Selector_2 s3532_7(wires_883_6[0], addr_883_6, addr_positional[14131:14128], addr_3532_7);

wire[31:0] addr_3533_7;

Selector_2 s3533_7(wires_883_6[1], addr_883_6, addr_positional[14135:14132], addr_3533_7);

wire[31:0] addr_3534_7;

Selector_2 s3534_7(wires_883_6[2], addr_883_6, addr_positional[14139:14136], addr_3534_7);

wire[31:0] addr_3535_7;

Selector_2 s3535_7(wires_883_6[3], addr_883_6, addr_positional[14143:14140], addr_3535_7);

wire[31:0] addr_3536_7;

Selector_2 s3536_7(wires_884_6[0], addr_884_6, addr_positional[14147:14144], addr_3536_7);

wire[31:0] addr_3537_7;

Selector_2 s3537_7(wires_884_6[1], addr_884_6, addr_positional[14151:14148], addr_3537_7);

wire[31:0] addr_3538_7;

Selector_2 s3538_7(wires_884_6[2], addr_884_6, addr_positional[14155:14152], addr_3538_7);

wire[31:0] addr_3539_7;

Selector_2 s3539_7(wires_884_6[3], addr_884_6, addr_positional[14159:14156], addr_3539_7);

wire[31:0] addr_3540_7;

Selector_2 s3540_7(wires_885_6[0], addr_885_6, addr_positional[14163:14160], addr_3540_7);

wire[31:0] addr_3541_7;

Selector_2 s3541_7(wires_885_6[1], addr_885_6, addr_positional[14167:14164], addr_3541_7);

wire[31:0] addr_3542_7;

Selector_2 s3542_7(wires_885_6[2], addr_885_6, addr_positional[14171:14168], addr_3542_7);

wire[31:0] addr_3543_7;

Selector_2 s3543_7(wires_885_6[3], addr_885_6, addr_positional[14175:14172], addr_3543_7);

wire[31:0] addr_3544_7;

Selector_2 s3544_7(wires_886_6[0], addr_886_6, addr_positional[14179:14176], addr_3544_7);

wire[31:0] addr_3545_7;

Selector_2 s3545_7(wires_886_6[1], addr_886_6, addr_positional[14183:14180], addr_3545_7);

wire[31:0] addr_3546_7;

Selector_2 s3546_7(wires_886_6[2], addr_886_6, addr_positional[14187:14184], addr_3546_7);

wire[31:0] addr_3547_7;

Selector_2 s3547_7(wires_886_6[3], addr_886_6, addr_positional[14191:14188], addr_3547_7);

wire[31:0] addr_3548_7;

Selector_2 s3548_7(wires_887_6[0], addr_887_6, addr_positional[14195:14192], addr_3548_7);

wire[31:0] addr_3549_7;

Selector_2 s3549_7(wires_887_6[1], addr_887_6, addr_positional[14199:14196], addr_3549_7);

wire[31:0] addr_3550_7;

Selector_2 s3550_7(wires_887_6[2], addr_887_6, addr_positional[14203:14200], addr_3550_7);

wire[31:0] addr_3551_7;

Selector_2 s3551_7(wires_887_6[3], addr_887_6, addr_positional[14207:14204], addr_3551_7);

wire[31:0] addr_3552_7;

Selector_2 s3552_7(wires_888_6[0], addr_888_6, addr_positional[14211:14208], addr_3552_7);

wire[31:0] addr_3553_7;

Selector_2 s3553_7(wires_888_6[1], addr_888_6, addr_positional[14215:14212], addr_3553_7);

wire[31:0] addr_3554_7;

Selector_2 s3554_7(wires_888_6[2], addr_888_6, addr_positional[14219:14216], addr_3554_7);

wire[31:0] addr_3555_7;

Selector_2 s3555_7(wires_888_6[3], addr_888_6, addr_positional[14223:14220], addr_3555_7);

wire[31:0] addr_3556_7;

Selector_2 s3556_7(wires_889_6[0], addr_889_6, addr_positional[14227:14224], addr_3556_7);

wire[31:0] addr_3557_7;

Selector_2 s3557_7(wires_889_6[1], addr_889_6, addr_positional[14231:14228], addr_3557_7);

wire[31:0] addr_3558_7;

Selector_2 s3558_7(wires_889_6[2], addr_889_6, addr_positional[14235:14232], addr_3558_7);

wire[31:0] addr_3559_7;

Selector_2 s3559_7(wires_889_6[3], addr_889_6, addr_positional[14239:14236], addr_3559_7);

wire[31:0] addr_3560_7;

Selector_2 s3560_7(wires_890_6[0], addr_890_6, addr_positional[14243:14240], addr_3560_7);

wire[31:0] addr_3561_7;

Selector_2 s3561_7(wires_890_6[1], addr_890_6, addr_positional[14247:14244], addr_3561_7);

wire[31:0] addr_3562_7;

Selector_2 s3562_7(wires_890_6[2], addr_890_6, addr_positional[14251:14248], addr_3562_7);

wire[31:0] addr_3563_7;

Selector_2 s3563_7(wires_890_6[3], addr_890_6, addr_positional[14255:14252], addr_3563_7);

wire[31:0] addr_3564_7;

Selector_2 s3564_7(wires_891_6[0], addr_891_6, addr_positional[14259:14256], addr_3564_7);

wire[31:0] addr_3565_7;

Selector_2 s3565_7(wires_891_6[1], addr_891_6, addr_positional[14263:14260], addr_3565_7);

wire[31:0] addr_3566_7;

Selector_2 s3566_7(wires_891_6[2], addr_891_6, addr_positional[14267:14264], addr_3566_7);

wire[31:0] addr_3567_7;

Selector_2 s3567_7(wires_891_6[3], addr_891_6, addr_positional[14271:14268], addr_3567_7);

wire[31:0] addr_3568_7;

Selector_2 s3568_7(wires_892_6[0], addr_892_6, addr_positional[14275:14272], addr_3568_7);

wire[31:0] addr_3569_7;

Selector_2 s3569_7(wires_892_6[1], addr_892_6, addr_positional[14279:14276], addr_3569_7);

wire[31:0] addr_3570_7;

Selector_2 s3570_7(wires_892_6[2], addr_892_6, addr_positional[14283:14280], addr_3570_7);

wire[31:0] addr_3571_7;

Selector_2 s3571_7(wires_892_6[3], addr_892_6, addr_positional[14287:14284], addr_3571_7);

wire[31:0] addr_3572_7;

Selector_2 s3572_7(wires_893_6[0], addr_893_6, addr_positional[14291:14288], addr_3572_7);

wire[31:0] addr_3573_7;

Selector_2 s3573_7(wires_893_6[1], addr_893_6, addr_positional[14295:14292], addr_3573_7);

wire[31:0] addr_3574_7;

Selector_2 s3574_7(wires_893_6[2], addr_893_6, addr_positional[14299:14296], addr_3574_7);

wire[31:0] addr_3575_7;

Selector_2 s3575_7(wires_893_6[3], addr_893_6, addr_positional[14303:14300], addr_3575_7);

wire[31:0] addr_3576_7;

Selector_2 s3576_7(wires_894_6[0], addr_894_6, addr_positional[14307:14304], addr_3576_7);

wire[31:0] addr_3577_7;

Selector_2 s3577_7(wires_894_6[1], addr_894_6, addr_positional[14311:14308], addr_3577_7);

wire[31:0] addr_3578_7;

Selector_2 s3578_7(wires_894_6[2], addr_894_6, addr_positional[14315:14312], addr_3578_7);

wire[31:0] addr_3579_7;

Selector_2 s3579_7(wires_894_6[3], addr_894_6, addr_positional[14319:14316], addr_3579_7);

wire[31:0] addr_3580_7;

Selector_2 s3580_7(wires_895_6[0], addr_895_6, addr_positional[14323:14320], addr_3580_7);

wire[31:0] addr_3581_7;

Selector_2 s3581_7(wires_895_6[1], addr_895_6, addr_positional[14327:14324], addr_3581_7);

wire[31:0] addr_3582_7;

Selector_2 s3582_7(wires_895_6[2], addr_895_6, addr_positional[14331:14328], addr_3582_7);

wire[31:0] addr_3583_7;

Selector_2 s3583_7(wires_895_6[3], addr_895_6, addr_positional[14335:14332], addr_3583_7);

wire[31:0] addr_3584_7;

Selector_2 s3584_7(wires_896_6[0], addr_896_6, addr_positional[14339:14336], addr_3584_7);

wire[31:0] addr_3585_7;

Selector_2 s3585_7(wires_896_6[1], addr_896_6, addr_positional[14343:14340], addr_3585_7);

wire[31:0] addr_3586_7;

Selector_2 s3586_7(wires_896_6[2], addr_896_6, addr_positional[14347:14344], addr_3586_7);

wire[31:0] addr_3587_7;

Selector_2 s3587_7(wires_896_6[3], addr_896_6, addr_positional[14351:14348], addr_3587_7);

wire[31:0] addr_3588_7;

Selector_2 s3588_7(wires_897_6[0], addr_897_6, addr_positional[14355:14352], addr_3588_7);

wire[31:0] addr_3589_7;

Selector_2 s3589_7(wires_897_6[1], addr_897_6, addr_positional[14359:14356], addr_3589_7);

wire[31:0] addr_3590_7;

Selector_2 s3590_7(wires_897_6[2], addr_897_6, addr_positional[14363:14360], addr_3590_7);

wire[31:0] addr_3591_7;

Selector_2 s3591_7(wires_897_6[3], addr_897_6, addr_positional[14367:14364], addr_3591_7);

wire[31:0] addr_3592_7;

Selector_2 s3592_7(wires_898_6[0], addr_898_6, addr_positional[14371:14368], addr_3592_7);

wire[31:0] addr_3593_7;

Selector_2 s3593_7(wires_898_6[1], addr_898_6, addr_positional[14375:14372], addr_3593_7);

wire[31:0] addr_3594_7;

Selector_2 s3594_7(wires_898_6[2], addr_898_6, addr_positional[14379:14376], addr_3594_7);

wire[31:0] addr_3595_7;

Selector_2 s3595_7(wires_898_6[3], addr_898_6, addr_positional[14383:14380], addr_3595_7);

wire[31:0] addr_3596_7;

Selector_2 s3596_7(wires_899_6[0], addr_899_6, addr_positional[14387:14384], addr_3596_7);

wire[31:0] addr_3597_7;

Selector_2 s3597_7(wires_899_6[1], addr_899_6, addr_positional[14391:14388], addr_3597_7);

wire[31:0] addr_3598_7;

Selector_2 s3598_7(wires_899_6[2], addr_899_6, addr_positional[14395:14392], addr_3598_7);

wire[31:0] addr_3599_7;

Selector_2 s3599_7(wires_899_6[3], addr_899_6, addr_positional[14399:14396], addr_3599_7);

wire[31:0] addr_3600_7;

Selector_2 s3600_7(wires_900_6[0], addr_900_6, addr_positional[14403:14400], addr_3600_7);

wire[31:0] addr_3601_7;

Selector_2 s3601_7(wires_900_6[1], addr_900_6, addr_positional[14407:14404], addr_3601_7);

wire[31:0] addr_3602_7;

Selector_2 s3602_7(wires_900_6[2], addr_900_6, addr_positional[14411:14408], addr_3602_7);

wire[31:0] addr_3603_7;

Selector_2 s3603_7(wires_900_6[3], addr_900_6, addr_positional[14415:14412], addr_3603_7);

wire[31:0] addr_3604_7;

Selector_2 s3604_7(wires_901_6[0], addr_901_6, addr_positional[14419:14416], addr_3604_7);

wire[31:0] addr_3605_7;

Selector_2 s3605_7(wires_901_6[1], addr_901_6, addr_positional[14423:14420], addr_3605_7);

wire[31:0] addr_3606_7;

Selector_2 s3606_7(wires_901_6[2], addr_901_6, addr_positional[14427:14424], addr_3606_7);

wire[31:0] addr_3607_7;

Selector_2 s3607_7(wires_901_6[3], addr_901_6, addr_positional[14431:14428], addr_3607_7);

wire[31:0] addr_3608_7;

Selector_2 s3608_7(wires_902_6[0], addr_902_6, addr_positional[14435:14432], addr_3608_7);

wire[31:0] addr_3609_7;

Selector_2 s3609_7(wires_902_6[1], addr_902_6, addr_positional[14439:14436], addr_3609_7);

wire[31:0] addr_3610_7;

Selector_2 s3610_7(wires_902_6[2], addr_902_6, addr_positional[14443:14440], addr_3610_7);

wire[31:0] addr_3611_7;

Selector_2 s3611_7(wires_902_6[3], addr_902_6, addr_positional[14447:14444], addr_3611_7);

wire[31:0] addr_3612_7;

Selector_2 s3612_7(wires_903_6[0], addr_903_6, addr_positional[14451:14448], addr_3612_7);

wire[31:0] addr_3613_7;

Selector_2 s3613_7(wires_903_6[1], addr_903_6, addr_positional[14455:14452], addr_3613_7);

wire[31:0] addr_3614_7;

Selector_2 s3614_7(wires_903_6[2], addr_903_6, addr_positional[14459:14456], addr_3614_7);

wire[31:0] addr_3615_7;

Selector_2 s3615_7(wires_903_6[3], addr_903_6, addr_positional[14463:14460], addr_3615_7);

wire[31:0] addr_3616_7;

Selector_2 s3616_7(wires_904_6[0], addr_904_6, addr_positional[14467:14464], addr_3616_7);

wire[31:0] addr_3617_7;

Selector_2 s3617_7(wires_904_6[1], addr_904_6, addr_positional[14471:14468], addr_3617_7);

wire[31:0] addr_3618_7;

Selector_2 s3618_7(wires_904_6[2], addr_904_6, addr_positional[14475:14472], addr_3618_7);

wire[31:0] addr_3619_7;

Selector_2 s3619_7(wires_904_6[3], addr_904_6, addr_positional[14479:14476], addr_3619_7);

wire[31:0] addr_3620_7;

Selector_2 s3620_7(wires_905_6[0], addr_905_6, addr_positional[14483:14480], addr_3620_7);

wire[31:0] addr_3621_7;

Selector_2 s3621_7(wires_905_6[1], addr_905_6, addr_positional[14487:14484], addr_3621_7);

wire[31:0] addr_3622_7;

Selector_2 s3622_7(wires_905_6[2], addr_905_6, addr_positional[14491:14488], addr_3622_7);

wire[31:0] addr_3623_7;

Selector_2 s3623_7(wires_905_6[3], addr_905_6, addr_positional[14495:14492], addr_3623_7);

wire[31:0] addr_3624_7;

Selector_2 s3624_7(wires_906_6[0], addr_906_6, addr_positional[14499:14496], addr_3624_7);

wire[31:0] addr_3625_7;

Selector_2 s3625_7(wires_906_6[1], addr_906_6, addr_positional[14503:14500], addr_3625_7);

wire[31:0] addr_3626_7;

Selector_2 s3626_7(wires_906_6[2], addr_906_6, addr_positional[14507:14504], addr_3626_7);

wire[31:0] addr_3627_7;

Selector_2 s3627_7(wires_906_6[3], addr_906_6, addr_positional[14511:14508], addr_3627_7);

wire[31:0] addr_3628_7;

Selector_2 s3628_7(wires_907_6[0], addr_907_6, addr_positional[14515:14512], addr_3628_7);

wire[31:0] addr_3629_7;

Selector_2 s3629_7(wires_907_6[1], addr_907_6, addr_positional[14519:14516], addr_3629_7);

wire[31:0] addr_3630_7;

Selector_2 s3630_7(wires_907_6[2], addr_907_6, addr_positional[14523:14520], addr_3630_7);

wire[31:0] addr_3631_7;

Selector_2 s3631_7(wires_907_6[3], addr_907_6, addr_positional[14527:14524], addr_3631_7);

wire[31:0] addr_3632_7;

Selector_2 s3632_7(wires_908_6[0], addr_908_6, addr_positional[14531:14528], addr_3632_7);

wire[31:0] addr_3633_7;

Selector_2 s3633_7(wires_908_6[1], addr_908_6, addr_positional[14535:14532], addr_3633_7);

wire[31:0] addr_3634_7;

Selector_2 s3634_7(wires_908_6[2], addr_908_6, addr_positional[14539:14536], addr_3634_7);

wire[31:0] addr_3635_7;

Selector_2 s3635_7(wires_908_6[3], addr_908_6, addr_positional[14543:14540], addr_3635_7);

wire[31:0] addr_3636_7;

Selector_2 s3636_7(wires_909_6[0], addr_909_6, addr_positional[14547:14544], addr_3636_7);

wire[31:0] addr_3637_7;

Selector_2 s3637_7(wires_909_6[1], addr_909_6, addr_positional[14551:14548], addr_3637_7);

wire[31:0] addr_3638_7;

Selector_2 s3638_7(wires_909_6[2], addr_909_6, addr_positional[14555:14552], addr_3638_7);

wire[31:0] addr_3639_7;

Selector_2 s3639_7(wires_909_6[3], addr_909_6, addr_positional[14559:14556], addr_3639_7);

wire[31:0] addr_3640_7;

Selector_2 s3640_7(wires_910_6[0], addr_910_6, addr_positional[14563:14560], addr_3640_7);

wire[31:0] addr_3641_7;

Selector_2 s3641_7(wires_910_6[1], addr_910_6, addr_positional[14567:14564], addr_3641_7);

wire[31:0] addr_3642_7;

Selector_2 s3642_7(wires_910_6[2], addr_910_6, addr_positional[14571:14568], addr_3642_7);

wire[31:0] addr_3643_7;

Selector_2 s3643_7(wires_910_6[3], addr_910_6, addr_positional[14575:14572], addr_3643_7);

wire[31:0] addr_3644_7;

Selector_2 s3644_7(wires_911_6[0], addr_911_6, addr_positional[14579:14576], addr_3644_7);

wire[31:0] addr_3645_7;

Selector_2 s3645_7(wires_911_6[1], addr_911_6, addr_positional[14583:14580], addr_3645_7);

wire[31:0] addr_3646_7;

Selector_2 s3646_7(wires_911_6[2], addr_911_6, addr_positional[14587:14584], addr_3646_7);

wire[31:0] addr_3647_7;

Selector_2 s3647_7(wires_911_6[3], addr_911_6, addr_positional[14591:14588], addr_3647_7);

wire[31:0] addr_3648_7;

Selector_2 s3648_7(wires_912_6[0], addr_912_6, addr_positional[14595:14592], addr_3648_7);

wire[31:0] addr_3649_7;

Selector_2 s3649_7(wires_912_6[1], addr_912_6, addr_positional[14599:14596], addr_3649_7);

wire[31:0] addr_3650_7;

Selector_2 s3650_7(wires_912_6[2], addr_912_6, addr_positional[14603:14600], addr_3650_7);

wire[31:0] addr_3651_7;

Selector_2 s3651_7(wires_912_6[3], addr_912_6, addr_positional[14607:14604], addr_3651_7);

wire[31:0] addr_3652_7;

Selector_2 s3652_7(wires_913_6[0], addr_913_6, addr_positional[14611:14608], addr_3652_7);

wire[31:0] addr_3653_7;

Selector_2 s3653_7(wires_913_6[1], addr_913_6, addr_positional[14615:14612], addr_3653_7);

wire[31:0] addr_3654_7;

Selector_2 s3654_7(wires_913_6[2], addr_913_6, addr_positional[14619:14616], addr_3654_7);

wire[31:0] addr_3655_7;

Selector_2 s3655_7(wires_913_6[3], addr_913_6, addr_positional[14623:14620], addr_3655_7);

wire[31:0] addr_3656_7;

Selector_2 s3656_7(wires_914_6[0], addr_914_6, addr_positional[14627:14624], addr_3656_7);

wire[31:0] addr_3657_7;

Selector_2 s3657_7(wires_914_6[1], addr_914_6, addr_positional[14631:14628], addr_3657_7);

wire[31:0] addr_3658_7;

Selector_2 s3658_7(wires_914_6[2], addr_914_6, addr_positional[14635:14632], addr_3658_7);

wire[31:0] addr_3659_7;

Selector_2 s3659_7(wires_914_6[3], addr_914_6, addr_positional[14639:14636], addr_3659_7);

wire[31:0] addr_3660_7;

Selector_2 s3660_7(wires_915_6[0], addr_915_6, addr_positional[14643:14640], addr_3660_7);

wire[31:0] addr_3661_7;

Selector_2 s3661_7(wires_915_6[1], addr_915_6, addr_positional[14647:14644], addr_3661_7);

wire[31:0] addr_3662_7;

Selector_2 s3662_7(wires_915_6[2], addr_915_6, addr_positional[14651:14648], addr_3662_7);

wire[31:0] addr_3663_7;

Selector_2 s3663_7(wires_915_6[3], addr_915_6, addr_positional[14655:14652], addr_3663_7);

wire[31:0] addr_3664_7;

Selector_2 s3664_7(wires_916_6[0], addr_916_6, addr_positional[14659:14656], addr_3664_7);

wire[31:0] addr_3665_7;

Selector_2 s3665_7(wires_916_6[1], addr_916_6, addr_positional[14663:14660], addr_3665_7);

wire[31:0] addr_3666_7;

Selector_2 s3666_7(wires_916_6[2], addr_916_6, addr_positional[14667:14664], addr_3666_7);

wire[31:0] addr_3667_7;

Selector_2 s3667_7(wires_916_6[3], addr_916_6, addr_positional[14671:14668], addr_3667_7);

wire[31:0] addr_3668_7;

Selector_2 s3668_7(wires_917_6[0], addr_917_6, addr_positional[14675:14672], addr_3668_7);

wire[31:0] addr_3669_7;

Selector_2 s3669_7(wires_917_6[1], addr_917_6, addr_positional[14679:14676], addr_3669_7);

wire[31:0] addr_3670_7;

Selector_2 s3670_7(wires_917_6[2], addr_917_6, addr_positional[14683:14680], addr_3670_7);

wire[31:0] addr_3671_7;

Selector_2 s3671_7(wires_917_6[3], addr_917_6, addr_positional[14687:14684], addr_3671_7);

wire[31:0] addr_3672_7;

Selector_2 s3672_7(wires_918_6[0], addr_918_6, addr_positional[14691:14688], addr_3672_7);

wire[31:0] addr_3673_7;

Selector_2 s3673_7(wires_918_6[1], addr_918_6, addr_positional[14695:14692], addr_3673_7);

wire[31:0] addr_3674_7;

Selector_2 s3674_7(wires_918_6[2], addr_918_6, addr_positional[14699:14696], addr_3674_7);

wire[31:0] addr_3675_7;

Selector_2 s3675_7(wires_918_6[3], addr_918_6, addr_positional[14703:14700], addr_3675_7);

wire[31:0] addr_3676_7;

Selector_2 s3676_7(wires_919_6[0], addr_919_6, addr_positional[14707:14704], addr_3676_7);

wire[31:0] addr_3677_7;

Selector_2 s3677_7(wires_919_6[1], addr_919_6, addr_positional[14711:14708], addr_3677_7);

wire[31:0] addr_3678_7;

Selector_2 s3678_7(wires_919_6[2], addr_919_6, addr_positional[14715:14712], addr_3678_7);

wire[31:0] addr_3679_7;

Selector_2 s3679_7(wires_919_6[3], addr_919_6, addr_positional[14719:14716], addr_3679_7);

wire[31:0] addr_3680_7;

Selector_2 s3680_7(wires_920_6[0], addr_920_6, addr_positional[14723:14720], addr_3680_7);

wire[31:0] addr_3681_7;

Selector_2 s3681_7(wires_920_6[1], addr_920_6, addr_positional[14727:14724], addr_3681_7);

wire[31:0] addr_3682_7;

Selector_2 s3682_7(wires_920_6[2], addr_920_6, addr_positional[14731:14728], addr_3682_7);

wire[31:0] addr_3683_7;

Selector_2 s3683_7(wires_920_6[3], addr_920_6, addr_positional[14735:14732], addr_3683_7);

wire[31:0] addr_3684_7;

Selector_2 s3684_7(wires_921_6[0], addr_921_6, addr_positional[14739:14736], addr_3684_7);

wire[31:0] addr_3685_7;

Selector_2 s3685_7(wires_921_6[1], addr_921_6, addr_positional[14743:14740], addr_3685_7);

wire[31:0] addr_3686_7;

Selector_2 s3686_7(wires_921_6[2], addr_921_6, addr_positional[14747:14744], addr_3686_7);

wire[31:0] addr_3687_7;

Selector_2 s3687_7(wires_921_6[3], addr_921_6, addr_positional[14751:14748], addr_3687_7);

wire[31:0] addr_3688_7;

Selector_2 s3688_7(wires_922_6[0], addr_922_6, addr_positional[14755:14752], addr_3688_7);

wire[31:0] addr_3689_7;

Selector_2 s3689_7(wires_922_6[1], addr_922_6, addr_positional[14759:14756], addr_3689_7);

wire[31:0] addr_3690_7;

Selector_2 s3690_7(wires_922_6[2], addr_922_6, addr_positional[14763:14760], addr_3690_7);

wire[31:0] addr_3691_7;

Selector_2 s3691_7(wires_922_6[3], addr_922_6, addr_positional[14767:14764], addr_3691_7);

wire[31:0] addr_3692_7;

Selector_2 s3692_7(wires_923_6[0], addr_923_6, addr_positional[14771:14768], addr_3692_7);

wire[31:0] addr_3693_7;

Selector_2 s3693_7(wires_923_6[1], addr_923_6, addr_positional[14775:14772], addr_3693_7);

wire[31:0] addr_3694_7;

Selector_2 s3694_7(wires_923_6[2], addr_923_6, addr_positional[14779:14776], addr_3694_7);

wire[31:0] addr_3695_7;

Selector_2 s3695_7(wires_923_6[3], addr_923_6, addr_positional[14783:14780], addr_3695_7);

wire[31:0] addr_3696_7;

Selector_2 s3696_7(wires_924_6[0], addr_924_6, addr_positional[14787:14784], addr_3696_7);

wire[31:0] addr_3697_7;

Selector_2 s3697_7(wires_924_6[1], addr_924_6, addr_positional[14791:14788], addr_3697_7);

wire[31:0] addr_3698_7;

Selector_2 s3698_7(wires_924_6[2], addr_924_6, addr_positional[14795:14792], addr_3698_7);

wire[31:0] addr_3699_7;

Selector_2 s3699_7(wires_924_6[3], addr_924_6, addr_positional[14799:14796], addr_3699_7);

wire[31:0] addr_3700_7;

Selector_2 s3700_7(wires_925_6[0], addr_925_6, addr_positional[14803:14800], addr_3700_7);

wire[31:0] addr_3701_7;

Selector_2 s3701_7(wires_925_6[1], addr_925_6, addr_positional[14807:14804], addr_3701_7);

wire[31:0] addr_3702_7;

Selector_2 s3702_7(wires_925_6[2], addr_925_6, addr_positional[14811:14808], addr_3702_7);

wire[31:0] addr_3703_7;

Selector_2 s3703_7(wires_925_6[3], addr_925_6, addr_positional[14815:14812], addr_3703_7);

wire[31:0] addr_3704_7;

Selector_2 s3704_7(wires_926_6[0], addr_926_6, addr_positional[14819:14816], addr_3704_7);

wire[31:0] addr_3705_7;

Selector_2 s3705_7(wires_926_6[1], addr_926_6, addr_positional[14823:14820], addr_3705_7);

wire[31:0] addr_3706_7;

Selector_2 s3706_7(wires_926_6[2], addr_926_6, addr_positional[14827:14824], addr_3706_7);

wire[31:0] addr_3707_7;

Selector_2 s3707_7(wires_926_6[3], addr_926_6, addr_positional[14831:14828], addr_3707_7);

wire[31:0] addr_3708_7;

Selector_2 s3708_7(wires_927_6[0], addr_927_6, addr_positional[14835:14832], addr_3708_7);

wire[31:0] addr_3709_7;

Selector_2 s3709_7(wires_927_6[1], addr_927_6, addr_positional[14839:14836], addr_3709_7);

wire[31:0] addr_3710_7;

Selector_2 s3710_7(wires_927_6[2], addr_927_6, addr_positional[14843:14840], addr_3710_7);

wire[31:0] addr_3711_7;

Selector_2 s3711_7(wires_927_6[3], addr_927_6, addr_positional[14847:14844], addr_3711_7);

wire[31:0] addr_3712_7;

Selector_2 s3712_7(wires_928_6[0], addr_928_6, addr_positional[14851:14848], addr_3712_7);

wire[31:0] addr_3713_7;

Selector_2 s3713_7(wires_928_6[1], addr_928_6, addr_positional[14855:14852], addr_3713_7);

wire[31:0] addr_3714_7;

Selector_2 s3714_7(wires_928_6[2], addr_928_6, addr_positional[14859:14856], addr_3714_7);

wire[31:0] addr_3715_7;

Selector_2 s3715_7(wires_928_6[3], addr_928_6, addr_positional[14863:14860], addr_3715_7);

wire[31:0] addr_3716_7;

Selector_2 s3716_7(wires_929_6[0], addr_929_6, addr_positional[14867:14864], addr_3716_7);

wire[31:0] addr_3717_7;

Selector_2 s3717_7(wires_929_6[1], addr_929_6, addr_positional[14871:14868], addr_3717_7);

wire[31:0] addr_3718_7;

Selector_2 s3718_7(wires_929_6[2], addr_929_6, addr_positional[14875:14872], addr_3718_7);

wire[31:0] addr_3719_7;

Selector_2 s3719_7(wires_929_6[3], addr_929_6, addr_positional[14879:14876], addr_3719_7);

wire[31:0] addr_3720_7;

Selector_2 s3720_7(wires_930_6[0], addr_930_6, addr_positional[14883:14880], addr_3720_7);

wire[31:0] addr_3721_7;

Selector_2 s3721_7(wires_930_6[1], addr_930_6, addr_positional[14887:14884], addr_3721_7);

wire[31:0] addr_3722_7;

Selector_2 s3722_7(wires_930_6[2], addr_930_6, addr_positional[14891:14888], addr_3722_7);

wire[31:0] addr_3723_7;

Selector_2 s3723_7(wires_930_6[3], addr_930_6, addr_positional[14895:14892], addr_3723_7);

wire[31:0] addr_3724_7;

Selector_2 s3724_7(wires_931_6[0], addr_931_6, addr_positional[14899:14896], addr_3724_7);

wire[31:0] addr_3725_7;

Selector_2 s3725_7(wires_931_6[1], addr_931_6, addr_positional[14903:14900], addr_3725_7);

wire[31:0] addr_3726_7;

Selector_2 s3726_7(wires_931_6[2], addr_931_6, addr_positional[14907:14904], addr_3726_7);

wire[31:0] addr_3727_7;

Selector_2 s3727_7(wires_931_6[3], addr_931_6, addr_positional[14911:14908], addr_3727_7);

wire[31:0] addr_3728_7;

Selector_2 s3728_7(wires_932_6[0], addr_932_6, addr_positional[14915:14912], addr_3728_7);

wire[31:0] addr_3729_7;

Selector_2 s3729_7(wires_932_6[1], addr_932_6, addr_positional[14919:14916], addr_3729_7);

wire[31:0] addr_3730_7;

Selector_2 s3730_7(wires_932_6[2], addr_932_6, addr_positional[14923:14920], addr_3730_7);

wire[31:0] addr_3731_7;

Selector_2 s3731_7(wires_932_6[3], addr_932_6, addr_positional[14927:14924], addr_3731_7);

wire[31:0] addr_3732_7;

Selector_2 s3732_7(wires_933_6[0], addr_933_6, addr_positional[14931:14928], addr_3732_7);

wire[31:0] addr_3733_7;

Selector_2 s3733_7(wires_933_6[1], addr_933_6, addr_positional[14935:14932], addr_3733_7);

wire[31:0] addr_3734_7;

Selector_2 s3734_7(wires_933_6[2], addr_933_6, addr_positional[14939:14936], addr_3734_7);

wire[31:0] addr_3735_7;

Selector_2 s3735_7(wires_933_6[3], addr_933_6, addr_positional[14943:14940], addr_3735_7);

wire[31:0] addr_3736_7;

Selector_2 s3736_7(wires_934_6[0], addr_934_6, addr_positional[14947:14944], addr_3736_7);

wire[31:0] addr_3737_7;

Selector_2 s3737_7(wires_934_6[1], addr_934_6, addr_positional[14951:14948], addr_3737_7);

wire[31:0] addr_3738_7;

Selector_2 s3738_7(wires_934_6[2], addr_934_6, addr_positional[14955:14952], addr_3738_7);

wire[31:0] addr_3739_7;

Selector_2 s3739_7(wires_934_6[3], addr_934_6, addr_positional[14959:14956], addr_3739_7);

wire[31:0] addr_3740_7;

Selector_2 s3740_7(wires_935_6[0], addr_935_6, addr_positional[14963:14960], addr_3740_7);

wire[31:0] addr_3741_7;

Selector_2 s3741_7(wires_935_6[1], addr_935_6, addr_positional[14967:14964], addr_3741_7);

wire[31:0] addr_3742_7;

Selector_2 s3742_7(wires_935_6[2], addr_935_6, addr_positional[14971:14968], addr_3742_7);

wire[31:0] addr_3743_7;

Selector_2 s3743_7(wires_935_6[3], addr_935_6, addr_positional[14975:14972], addr_3743_7);

wire[31:0] addr_3744_7;

Selector_2 s3744_7(wires_936_6[0], addr_936_6, addr_positional[14979:14976], addr_3744_7);

wire[31:0] addr_3745_7;

Selector_2 s3745_7(wires_936_6[1], addr_936_6, addr_positional[14983:14980], addr_3745_7);

wire[31:0] addr_3746_7;

Selector_2 s3746_7(wires_936_6[2], addr_936_6, addr_positional[14987:14984], addr_3746_7);

wire[31:0] addr_3747_7;

Selector_2 s3747_7(wires_936_6[3], addr_936_6, addr_positional[14991:14988], addr_3747_7);

wire[31:0] addr_3748_7;

Selector_2 s3748_7(wires_937_6[0], addr_937_6, addr_positional[14995:14992], addr_3748_7);

wire[31:0] addr_3749_7;

Selector_2 s3749_7(wires_937_6[1], addr_937_6, addr_positional[14999:14996], addr_3749_7);

wire[31:0] addr_3750_7;

Selector_2 s3750_7(wires_937_6[2], addr_937_6, addr_positional[15003:15000], addr_3750_7);

wire[31:0] addr_3751_7;

Selector_2 s3751_7(wires_937_6[3], addr_937_6, addr_positional[15007:15004], addr_3751_7);

wire[31:0] addr_3752_7;

Selector_2 s3752_7(wires_938_6[0], addr_938_6, addr_positional[15011:15008], addr_3752_7);

wire[31:0] addr_3753_7;

Selector_2 s3753_7(wires_938_6[1], addr_938_6, addr_positional[15015:15012], addr_3753_7);

wire[31:0] addr_3754_7;

Selector_2 s3754_7(wires_938_6[2], addr_938_6, addr_positional[15019:15016], addr_3754_7);

wire[31:0] addr_3755_7;

Selector_2 s3755_7(wires_938_6[3], addr_938_6, addr_positional[15023:15020], addr_3755_7);

wire[31:0] addr_3756_7;

Selector_2 s3756_7(wires_939_6[0], addr_939_6, addr_positional[15027:15024], addr_3756_7);

wire[31:0] addr_3757_7;

Selector_2 s3757_7(wires_939_6[1], addr_939_6, addr_positional[15031:15028], addr_3757_7);

wire[31:0] addr_3758_7;

Selector_2 s3758_7(wires_939_6[2], addr_939_6, addr_positional[15035:15032], addr_3758_7);

wire[31:0] addr_3759_7;

Selector_2 s3759_7(wires_939_6[3], addr_939_6, addr_positional[15039:15036], addr_3759_7);

wire[31:0] addr_3760_7;

Selector_2 s3760_7(wires_940_6[0], addr_940_6, addr_positional[15043:15040], addr_3760_7);

wire[31:0] addr_3761_7;

Selector_2 s3761_7(wires_940_6[1], addr_940_6, addr_positional[15047:15044], addr_3761_7);

wire[31:0] addr_3762_7;

Selector_2 s3762_7(wires_940_6[2], addr_940_6, addr_positional[15051:15048], addr_3762_7);

wire[31:0] addr_3763_7;

Selector_2 s3763_7(wires_940_6[3], addr_940_6, addr_positional[15055:15052], addr_3763_7);

wire[31:0] addr_3764_7;

Selector_2 s3764_7(wires_941_6[0], addr_941_6, addr_positional[15059:15056], addr_3764_7);

wire[31:0] addr_3765_7;

Selector_2 s3765_7(wires_941_6[1], addr_941_6, addr_positional[15063:15060], addr_3765_7);

wire[31:0] addr_3766_7;

Selector_2 s3766_7(wires_941_6[2], addr_941_6, addr_positional[15067:15064], addr_3766_7);

wire[31:0] addr_3767_7;

Selector_2 s3767_7(wires_941_6[3], addr_941_6, addr_positional[15071:15068], addr_3767_7);

wire[31:0] addr_3768_7;

Selector_2 s3768_7(wires_942_6[0], addr_942_6, addr_positional[15075:15072], addr_3768_7);

wire[31:0] addr_3769_7;

Selector_2 s3769_7(wires_942_6[1], addr_942_6, addr_positional[15079:15076], addr_3769_7);

wire[31:0] addr_3770_7;

Selector_2 s3770_7(wires_942_6[2], addr_942_6, addr_positional[15083:15080], addr_3770_7);

wire[31:0] addr_3771_7;

Selector_2 s3771_7(wires_942_6[3], addr_942_6, addr_positional[15087:15084], addr_3771_7);

wire[31:0] addr_3772_7;

Selector_2 s3772_7(wires_943_6[0], addr_943_6, addr_positional[15091:15088], addr_3772_7);

wire[31:0] addr_3773_7;

Selector_2 s3773_7(wires_943_6[1], addr_943_6, addr_positional[15095:15092], addr_3773_7);

wire[31:0] addr_3774_7;

Selector_2 s3774_7(wires_943_6[2], addr_943_6, addr_positional[15099:15096], addr_3774_7);

wire[31:0] addr_3775_7;

Selector_2 s3775_7(wires_943_6[3], addr_943_6, addr_positional[15103:15100], addr_3775_7);

wire[31:0] addr_3776_7;

Selector_2 s3776_7(wires_944_6[0], addr_944_6, addr_positional[15107:15104], addr_3776_7);

wire[31:0] addr_3777_7;

Selector_2 s3777_7(wires_944_6[1], addr_944_6, addr_positional[15111:15108], addr_3777_7);

wire[31:0] addr_3778_7;

Selector_2 s3778_7(wires_944_6[2], addr_944_6, addr_positional[15115:15112], addr_3778_7);

wire[31:0] addr_3779_7;

Selector_2 s3779_7(wires_944_6[3], addr_944_6, addr_positional[15119:15116], addr_3779_7);

wire[31:0] addr_3780_7;

Selector_2 s3780_7(wires_945_6[0], addr_945_6, addr_positional[15123:15120], addr_3780_7);

wire[31:0] addr_3781_7;

Selector_2 s3781_7(wires_945_6[1], addr_945_6, addr_positional[15127:15124], addr_3781_7);

wire[31:0] addr_3782_7;

Selector_2 s3782_7(wires_945_6[2], addr_945_6, addr_positional[15131:15128], addr_3782_7);

wire[31:0] addr_3783_7;

Selector_2 s3783_7(wires_945_6[3], addr_945_6, addr_positional[15135:15132], addr_3783_7);

wire[31:0] addr_3784_7;

Selector_2 s3784_7(wires_946_6[0], addr_946_6, addr_positional[15139:15136], addr_3784_7);

wire[31:0] addr_3785_7;

Selector_2 s3785_7(wires_946_6[1], addr_946_6, addr_positional[15143:15140], addr_3785_7);

wire[31:0] addr_3786_7;

Selector_2 s3786_7(wires_946_6[2], addr_946_6, addr_positional[15147:15144], addr_3786_7);

wire[31:0] addr_3787_7;

Selector_2 s3787_7(wires_946_6[3], addr_946_6, addr_positional[15151:15148], addr_3787_7);

wire[31:0] addr_3788_7;

Selector_2 s3788_7(wires_947_6[0], addr_947_6, addr_positional[15155:15152], addr_3788_7);

wire[31:0] addr_3789_7;

Selector_2 s3789_7(wires_947_6[1], addr_947_6, addr_positional[15159:15156], addr_3789_7);

wire[31:0] addr_3790_7;

Selector_2 s3790_7(wires_947_6[2], addr_947_6, addr_positional[15163:15160], addr_3790_7);

wire[31:0] addr_3791_7;

Selector_2 s3791_7(wires_947_6[3], addr_947_6, addr_positional[15167:15164], addr_3791_7);

wire[31:0] addr_3792_7;

Selector_2 s3792_7(wires_948_6[0], addr_948_6, addr_positional[15171:15168], addr_3792_7);

wire[31:0] addr_3793_7;

Selector_2 s3793_7(wires_948_6[1], addr_948_6, addr_positional[15175:15172], addr_3793_7);

wire[31:0] addr_3794_7;

Selector_2 s3794_7(wires_948_6[2], addr_948_6, addr_positional[15179:15176], addr_3794_7);

wire[31:0] addr_3795_7;

Selector_2 s3795_7(wires_948_6[3], addr_948_6, addr_positional[15183:15180], addr_3795_7);

wire[31:0] addr_3796_7;

Selector_2 s3796_7(wires_949_6[0], addr_949_6, addr_positional[15187:15184], addr_3796_7);

wire[31:0] addr_3797_7;

Selector_2 s3797_7(wires_949_6[1], addr_949_6, addr_positional[15191:15188], addr_3797_7);

wire[31:0] addr_3798_7;

Selector_2 s3798_7(wires_949_6[2], addr_949_6, addr_positional[15195:15192], addr_3798_7);

wire[31:0] addr_3799_7;

Selector_2 s3799_7(wires_949_6[3], addr_949_6, addr_positional[15199:15196], addr_3799_7);

wire[31:0] addr_3800_7;

Selector_2 s3800_7(wires_950_6[0], addr_950_6, addr_positional[15203:15200], addr_3800_7);

wire[31:0] addr_3801_7;

Selector_2 s3801_7(wires_950_6[1], addr_950_6, addr_positional[15207:15204], addr_3801_7);

wire[31:0] addr_3802_7;

Selector_2 s3802_7(wires_950_6[2], addr_950_6, addr_positional[15211:15208], addr_3802_7);

wire[31:0] addr_3803_7;

Selector_2 s3803_7(wires_950_6[3], addr_950_6, addr_positional[15215:15212], addr_3803_7);

wire[31:0] addr_3804_7;

Selector_2 s3804_7(wires_951_6[0], addr_951_6, addr_positional[15219:15216], addr_3804_7);

wire[31:0] addr_3805_7;

Selector_2 s3805_7(wires_951_6[1], addr_951_6, addr_positional[15223:15220], addr_3805_7);

wire[31:0] addr_3806_7;

Selector_2 s3806_7(wires_951_6[2], addr_951_6, addr_positional[15227:15224], addr_3806_7);

wire[31:0] addr_3807_7;

Selector_2 s3807_7(wires_951_6[3], addr_951_6, addr_positional[15231:15228], addr_3807_7);

wire[31:0] addr_3808_7;

Selector_2 s3808_7(wires_952_6[0], addr_952_6, addr_positional[15235:15232], addr_3808_7);

wire[31:0] addr_3809_7;

Selector_2 s3809_7(wires_952_6[1], addr_952_6, addr_positional[15239:15236], addr_3809_7);

wire[31:0] addr_3810_7;

Selector_2 s3810_7(wires_952_6[2], addr_952_6, addr_positional[15243:15240], addr_3810_7);

wire[31:0] addr_3811_7;

Selector_2 s3811_7(wires_952_6[3], addr_952_6, addr_positional[15247:15244], addr_3811_7);

wire[31:0] addr_3812_7;

Selector_2 s3812_7(wires_953_6[0], addr_953_6, addr_positional[15251:15248], addr_3812_7);

wire[31:0] addr_3813_7;

Selector_2 s3813_7(wires_953_6[1], addr_953_6, addr_positional[15255:15252], addr_3813_7);

wire[31:0] addr_3814_7;

Selector_2 s3814_7(wires_953_6[2], addr_953_6, addr_positional[15259:15256], addr_3814_7);

wire[31:0] addr_3815_7;

Selector_2 s3815_7(wires_953_6[3], addr_953_6, addr_positional[15263:15260], addr_3815_7);

wire[31:0] addr_3816_7;

Selector_2 s3816_7(wires_954_6[0], addr_954_6, addr_positional[15267:15264], addr_3816_7);

wire[31:0] addr_3817_7;

Selector_2 s3817_7(wires_954_6[1], addr_954_6, addr_positional[15271:15268], addr_3817_7);

wire[31:0] addr_3818_7;

Selector_2 s3818_7(wires_954_6[2], addr_954_6, addr_positional[15275:15272], addr_3818_7);

wire[31:0] addr_3819_7;

Selector_2 s3819_7(wires_954_6[3], addr_954_6, addr_positional[15279:15276], addr_3819_7);

wire[31:0] addr_3820_7;

Selector_2 s3820_7(wires_955_6[0], addr_955_6, addr_positional[15283:15280], addr_3820_7);

wire[31:0] addr_3821_7;

Selector_2 s3821_7(wires_955_6[1], addr_955_6, addr_positional[15287:15284], addr_3821_7);

wire[31:0] addr_3822_7;

Selector_2 s3822_7(wires_955_6[2], addr_955_6, addr_positional[15291:15288], addr_3822_7);

wire[31:0] addr_3823_7;

Selector_2 s3823_7(wires_955_6[3], addr_955_6, addr_positional[15295:15292], addr_3823_7);

wire[31:0] addr_3824_7;

Selector_2 s3824_7(wires_956_6[0], addr_956_6, addr_positional[15299:15296], addr_3824_7);

wire[31:0] addr_3825_7;

Selector_2 s3825_7(wires_956_6[1], addr_956_6, addr_positional[15303:15300], addr_3825_7);

wire[31:0] addr_3826_7;

Selector_2 s3826_7(wires_956_6[2], addr_956_6, addr_positional[15307:15304], addr_3826_7);

wire[31:0] addr_3827_7;

Selector_2 s3827_7(wires_956_6[3], addr_956_6, addr_positional[15311:15308], addr_3827_7);

wire[31:0] addr_3828_7;

Selector_2 s3828_7(wires_957_6[0], addr_957_6, addr_positional[15315:15312], addr_3828_7);

wire[31:0] addr_3829_7;

Selector_2 s3829_7(wires_957_6[1], addr_957_6, addr_positional[15319:15316], addr_3829_7);

wire[31:0] addr_3830_7;

Selector_2 s3830_7(wires_957_6[2], addr_957_6, addr_positional[15323:15320], addr_3830_7);

wire[31:0] addr_3831_7;

Selector_2 s3831_7(wires_957_6[3], addr_957_6, addr_positional[15327:15324], addr_3831_7);

wire[31:0] addr_3832_7;

Selector_2 s3832_7(wires_958_6[0], addr_958_6, addr_positional[15331:15328], addr_3832_7);

wire[31:0] addr_3833_7;

Selector_2 s3833_7(wires_958_6[1], addr_958_6, addr_positional[15335:15332], addr_3833_7);

wire[31:0] addr_3834_7;

Selector_2 s3834_7(wires_958_6[2], addr_958_6, addr_positional[15339:15336], addr_3834_7);

wire[31:0] addr_3835_7;

Selector_2 s3835_7(wires_958_6[3], addr_958_6, addr_positional[15343:15340], addr_3835_7);

wire[31:0] addr_3836_7;

Selector_2 s3836_7(wires_959_6[0], addr_959_6, addr_positional[15347:15344], addr_3836_7);

wire[31:0] addr_3837_7;

Selector_2 s3837_7(wires_959_6[1], addr_959_6, addr_positional[15351:15348], addr_3837_7);

wire[31:0] addr_3838_7;

Selector_2 s3838_7(wires_959_6[2], addr_959_6, addr_positional[15355:15352], addr_3838_7);

wire[31:0] addr_3839_7;

Selector_2 s3839_7(wires_959_6[3], addr_959_6, addr_positional[15359:15356], addr_3839_7);

wire[31:0] addr_3840_7;

Selector_2 s3840_7(wires_960_6[0], addr_960_6, addr_positional[15363:15360], addr_3840_7);

wire[31:0] addr_3841_7;

Selector_2 s3841_7(wires_960_6[1], addr_960_6, addr_positional[15367:15364], addr_3841_7);

wire[31:0] addr_3842_7;

Selector_2 s3842_7(wires_960_6[2], addr_960_6, addr_positional[15371:15368], addr_3842_7);

wire[31:0] addr_3843_7;

Selector_2 s3843_7(wires_960_6[3], addr_960_6, addr_positional[15375:15372], addr_3843_7);

wire[31:0] addr_3844_7;

Selector_2 s3844_7(wires_961_6[0], addr_961_6, addr_positional[15379:15376], addr_3844_7);

wire[31:0] addr_3845_7;

Selector_2 s3845_7(wires_961_6[1], addr_961_6, addr_positional[15383:15380], addr_3845_7);

wire[31:0] addr_3846_7;

Selector_2 s3846_7(wires_961_6[2], addr_961_6, addr_positional[15387:15384], addr_3846_7);

wire[31:0] addr_3847_7;

Selector_2 s3847_7(wires_961_6[3], addr_961_6, addr_positional[15391:15388], addr_3847_7);

wire[31:0] addr_3848_7;

Selector_2 s3848_7(wires_962_6[0], addr_962_6, addr_positional[15395:15392], addr_3848_7);

wire[31:0] addr_3849_7;

Selector_2 s3849_7(wires_962_6[1], addr_962_6, addr_positional[15399:15396], addr_3849_7);

wire[31:0] addr_3850_7;

Selector_2 s3850_7(wires_962_6[2], addr_962_6, addr_positional[15403:15400], addr_3850_7);

wire[31:0] addr_3851_7;

Selector_2 s3851_7(wires_962_6[3], addr_962_6, addr_positional[15407:15404], addr_3851_7);

wire[31:0] addr_3852_7;

Selector_2 s3852_7(wires_963_6[0], addr_963_6, addr_positional[15411:15408], addr_3852_7);

wire[31:0] addr_3853_7;

Selector_2 s3853_7(wires_963_6[1], addr_963_6, addr_positional[15415:15412], addr_3853_7);

wire[31:0] addr_3854_7;

Selector_2 s3854_7(wires_963_6[2], addr_963_6, addr_positional[15419:15416], addr_3854_7);

wire[31:0] addr_3855_7;

Selector_2 s3855_7(wires_963_6[3], addr_963_6, addr_positional[15423:15420], addr_3855_7);

wire[31:0] addr_3856_7;

Selector_2 s3856_7(wires_964_6[0], addr_964_6, addr_positional[15427:15424], addr_3856_7);

wire[31:0] addr_3857_7;

Selector_2 s3857_7(wires_964_6[1], addr_964_6, addr_positional[15431:15428], addr_3857_7);

wire[31:0] addr_3858_7;

Selector_2 s3858_7(wires_964_6[2], addr_964_6, addr_positional[15435:15432], addr_3858_7);

wire[31:0] addr_3859_7;

Selector_2 s3859_7(wires_964_6[3], addr_964_6, addr_positional[15439:15436], addr_3859_7);

wire[31:0] addr_3860_7;

Selector_2 s3860_7(wires_965_6[0], addr_965_6, addr_positional[15443:15440], addr_3860_7);

wire[31:0] addr_3861_7;

Selector_2 s3861_7(wires_965_6[1], addr_965_6, addr_positional[15447:15444], addr_3861_7);

wire[31:0] addr_3862_7;

Selector_2 s3862_7(wires_965_6[2], addr_965_6, addr_positional[15451:15448], addr_3862_7);

wire[31:0] addr_3863_7;

Selector_2 s3863_7(wires_965_6[3], addr_965_6, addr_positional[15455:15452], addr_3863_7);

wire[31:0] addr_3864_7;

Selector_2 s3864_7(wires_966_6[0], addr_966_6, addr_positional[15459:15456], addr_3864_7);

wire[31:0] addr_3865_7;

Selector_2 s3865_7(wires_966_6[1], addr_966_6, addr_positional[15463:15460], addr_3865_7);

wire[31:0] addr_3866_7;

Selector_2 s3866_7(wires_966_6[2], addr_966_6, addr_positional[15467:15464], addr_3866_7);

wire[31:0] addr_3867_7;

Selector_2 s3867_7(wires_966_6[3], addr_966_6, addr_positional[15471:15468], addr_3867_7);

wire[31:0] addr_3868_7;

Selector_2 s3868_7(wires_967_6[0], addr_967_6, addr_positional[15475:15472], addr_3868_7);

wire[31:0] addr_3869_7;

Selector_2 s3869_7(wires_967_6[1], addr_967_6, addr_positional[15479:15476], addr_3869_7);

wire[31:0] addr_3870_7;

Selector_2 s3870_7(wires_967_6[2], addr_967_6, addr_positional[15483:15480], addr_3870_7);

wire[31:0] addr_3871_7;

Selector_2 s3871_7(wires_967_6[3], addr_967_6, addr_positional[15487:15484], addr_3871_7);

wire[31:0] addr_3872_7;

Selector_2 s3872_7(wires_968_6[0], addr_968_6, addr_positional[15491:15488], addr_3872_7);

wire[31:0] addr_3873_7;

Selector_2 s3873_7(wires_968_6[1], addr_968_6, addr_positional[15495:15492], addr_3873_7);

wire[31:0] addr_3874_7;

Selector_2 s3874_7(wires_968_6[2], addr_968_6, addr_positional[15499:15496], addr_3874_7);

wire[31:0] addr_3875_7;

Selector_2 s3875_7(wires_968_6[3], addr_968_6, addr_positional[15503:15500], addr_3875_7);

wire[31:0] addr_3876_7;

Selector_2 s3876_7(wires_969_6[0], addr_969_6, addr_positional[15507:15504], addr_3876_7);

wire[31:0] addr_3877_7;

Selector_2 s3877_7(wires_969_6[1], addr_969_6, addr_positional[15511:15508], addr_3877_7);

wire[31:0] addr_3878_7;

Selector_2 s3878_7(wires_969_6[2], addr_969_6, addr_positional[15515:15512], addr_3878_7);

wire[31:0] addr_3879_7;

Selector_2 s3879_7(wires_969_6[3], addr_969_6, addr_positional[15519:15516], addr_3879_7);

wire[31:0] addr_3880_7;

Selector_2 s3880_7(wires_970_6[0], addr_970_6, addr_positional[15523:15520], addr_3880_7);

wire[31:0] addr_3881_7;

Selector_2 s3881_7(wires_970_6[1], addr_970_6, addr_positional[15527:15524], addr_3881_7);

wire[31:0] addr_3882_7;

Selector_2 s3882_7(wires_970_6[2], addr_970_6, addr_positional[15531:15528], addr_3882_7);

wire[31:0] addr_3883_7;

Selector_2 s3883_7(wires_970_6[3], addr_970_6, addr_positional[15535:15532], addr_3883_7);

wire[31:0] addr_3884_7;

Selector_2 s3884_7(wires_971_6[0], addr_971_6, addr_positional[15539:15536], addr_3884_7);

wire[31:0] addr_3885_7;

Selector_2 s3885_7(wires_971_6[1], addr_971_6, addr_positional[15543:15540], addr_3885_7);

wire[31:0] addr_3886_7;

Selector_2 s3886_7(wires_971_6[2], addr_971_6, addr_positional[15547:15544], addr_3886_7);

wire[31:0] addr_3887_7;

Selector_2 s3887_7(wires_971_6[3], addr_971_6, addr_positional[15551:15548], addr_3887_7);

wire[31:0] addr_3888_7;

Selector_2 s3888_7(wires_972_6[0], addr_972_6, addr_positional[15555:15552], addr_3888_7);

wire[31:0] addr_3889_7;

Selector_2 s3889_7(wires_972_6[1], addr_972_6, addr_positional[15559:15556], addr_3889_7);

wire[31:0] addr_3890_7;

Selector_2 s3890_7(wires_972_6[2], addr_972_6, addr_positional[15563:15560], addr_3890_7);

wire[31:0] addr_3891_7;

Selector_2 s3891_7(wires_972_6[3], addr_972_6, addr_positional[15567:15564], addr_3891_7);

wire[31:0] addr_3892_7;

Selector_2 s3892_7(wires_973_6[0], addr_973_6, addr_positional[15571:15568], addr_3892_7);

wire[31:0] addr_3893_7;

Selector_2 s3893_7(wires_973_6[1], addr_973_6, addr_positional[15575:15572], addr_3893_7);

wire[31:0] addr_3894_7;

Selector_2 s3894_7(wires_973_6[2], addr_973_6, addr_positional[15579:15576], addr_3894_7);

wire[31:0] addr_3895_7;

Selector_2 s3895_7(wires_973_6[3], addr_973_6, addr_positional[15583:15580], addr_3895_7);

wire[31:0] addr_3896_7;

Selector_2 s3896_7(wires_974_6[0], addr_974_6, addr_positional[15587:15584], addr_3896_7);

wire[31:0] addr_3897_7;

Selector_2 s3897_7(wires_974_6[1], addr_974_6, addr_positional[15591:15588], addr_3897_7);

wire[31:0] addr_3898_7;

Selector_2 s3898_7(wires_974_6[2], addr_974_6, addr_positional[15595:15592], addr_3898_7);

wire[31:0] addr_3899_7;

Selector_2 s3899_7(wires_974_6[3], addr_974_6, addr_positional[15599:15596], addr_3899_7);

wire[31:0] addr_3900_7;

Selector_2 s3900_7(wires_975_6[0], addr_975_6, addr_positional[15603:15600], addr_3900_7);

wire[31:0] addr_3901_7;

Selector_2 s3901_7(wires_975_6[1], addr_975_6, addr_positional[15607:15604], addr_3901_7);

wire[31:0] addr_3902_7;

Selector_2 s3902_7(wires_975_6[2], addr_975_6, addr_positional[15611:15608], addr_3902_7);

wire[31:0] addr_3903_7;

Selector_2 s3903_7(wires_975_6[3], addr_975_6, addr_positional[15615:15612], addr_3903_7);

wire[31:0] addr_3904_7;

Selector_2 s3904_7(wires_976_6[0], addr_976_6, addr_positional[15619:15616], addr_3904_7);

wire[31:0] addr_3905_7;

Selector_2 s3905_7(wires_976_6[1], addr_976_6, addr_positional[15623:15620], addr_3905_7);

wire[31:0] addr_3906_7;

Selector_2 s3906_7(wires_976_6[2], addr_976_6, addr_positional[15627:15624], addr_3906_7);

wire[31:0] addr_3907_7;

Selector_2 s3907_7(wires_976_6[3], addr_976_6, addr_positional[15631:15628], addr_3907_7);

wire[31:0] addr_3908_7;

Selector_2 s3908_7(wires_977_6[0], addr_977_6, addr_positional[15635:15632], addr_3908_7);

wire[31:0] addr_3909_7;

Selector_2 s3909_7(wires_977_6[1], addr_977_6, addr_positional[15639:15636], addr_3909_7);

wire[31:0] addr_3910_7;

Selector_2 s3910_7(wires_977_6[2], addr_977_6, addr_positional[15643:15640], addr_3910_7);

wire[31:0] addr_3911_7;

Selector_2 s3911_7(wires_977_6[3], addr_977_6, addr_positional[15647:15644], addr_3911_7);

wire[31:0] addr_3912_7;

Selector_2 s3912_7(wires_978_6[0], addr_978_6, addr_positional[15651:15648], addr_3912_7);

wire[31:0] addr_3913_7;

Selector_2 s3913_7(wires_978_6[1], addr_978_6, addr_positional[15655:15652], addr_3913_7);

wire[31:0] addr_3914_7;

Selector_2 s3914_7(wires_978_6[2], addr_978_6, addr_positional[15659:15656], addr_3914_7);

wire[31:0] addr_3915_7;

Selector_2 s3915_7(wires_978_6[3], addr_978_6, addr_positional[15663:15660], addr_3915_7);

wire[31:0] addr_3916_7;

Selector_2 s3916_7(wires_979_6[0], addr_979_6, addr_positional[15667:15664], addr_3916_7);

wire[31:0] addr_3917_7;

Selector_2 s3917_7(wires_979_6[1], addr_979_6, addr_positional[15671:15668], addr_3917_7);

wire[31:0] addr_3918_7;

Selector_2 s3918_7(wires_979_6[2], addr_979_6, addr_positional[15675:15672], addr_3918_7);

wire[31:0] addr_3919_7;

Selector_2 s3919_7(wires_979_6[3], addr_979_6, addr_positional[15679:15676], addr_3919_7);

wire[31:0] addr_3920_7;

Selector_2 s3920_7(wires_980_6[0], addr_980_6, addr_positional[15683:15680], addr_3920_7);

wire[31:0] addr_3921_7;

Selector_2 s3921_7(wires_980_6[1], addr_980_6, addr_positional[15687:15684], addr_3921_7);

wire[31:0] addr_3922_7;

Selector_2 s3922_7(wires_980_6[2], addr_980_6, addr_positional[15691:15688], addr_3922_7);

wire[31:0] addr_3923_7;

Selector_2 s3923_7(wires_980_6[3], addr_980_6, addr_positional[15695:15692], addr_3923_7);

wire[31:0] addr_3924_7;

Selector_2 s3924_7(wires_981_6[0], addr_981_6, addr_positional[15699:15696], addr_3924_7);

wire[31:0] addr_3925_7;

Selector_2 s3925_7(wires_981_6[1], addr_981_6, addr_positional[15703:15700], addr_3925_7);

wire[31:0] addr_3926_7;

Selector_2 s3926_7(wires_981_6[2], addr_981_6, addr_positional[15707:15704], addr_3926_7);

wire[31:0] addr_3927_7;

Selector_2 s3927_7(wires_981_6[3], addr_981_6, addr_positional[15711:15708], addr_3927_7);

wire[31:0] addr_3928_7;

Selector_2 s3928_7(wires_982_6[0], addr_982_6, addr_positional[15715:15712], addr_3928_7);

wire[31:0] addr_3929_7;

Selector_2 s3929_7(wires_982_6[1], addr_982_6, addr_positional[15719:15716], addr_3929_7);

wire[31:0] addr_3930_7;

Selector_2 s3930_7(wires_982_6[2], addr_982_6, addr_positional[15723:15720], addr_3930_7);

wire[31:0] addr_3931_7;

Selector_2 s3931_7(wires_982_6[3], addr_982_6, addr_positional[15727:15724], addr_3931_7);

wire[31:0] addr_3932_7;

Selector_2 s3932_7(wires_983_6[0], addr_983_6, addr_positional[15731:15728], addr_3932_7);

wire[31:0] addr_3933_7;

Selector_2 s3933_7(wires_983_6[1], addr_983_6, addr_positional[15735:15732], addr_3933_7);

wire[31:0] addr_3934_7;

Selector_2 s3934_7(wires_983_6[2], addr_983_6, addr_positional[15739:15736], addr_3934_7);

wire[31:0] addr_3935_7;

Selector_2 s3935_7(wires_983_6[3], addr_983_6, addr_positional[15743:15740], addr_3935_7);

wire[31:0] addr_3936_7;

Selector_2 s3936_7(wires_984_6[0], addr_984_6, addr_positional[15747:15744], addr_3936_7);

wire[31:0] addr_3937_7;

Selector_2 s3937_7(wires_984_6[1], addr_984_6, addr_positional[15751:15748], addr_3937_7);

wire[31:0] addr_3938_7;

Selector_2 s3938_7(wires_984_6[2], addr_984_6, addr_positional[15755:15752], addr_3938_7);

wire[31:0] addr_3939_7;

Selector_2 s3939_7(wires_984_6[3], addr_984_6, addr_positional[15759:15756], addr_3939_7);

wire[31:0] addr_3940_7;

Selector_2 s3940_7(wires_985_6[0], addr_985_6, addr_positional[15763:15760], addr_3940_7);

wire[31:0] addr_3941_7;

Selector_2 s3941_7(wires_985_6[1], addr_985_6, addr_positional[15767:15764], addr_3941_7);

wire[31:0] addr_3942_7;

Selector_2 s3942_7(wires_985_6[2], addr_985_6, addr_positional[15771:15768], addr_3942_7);

wire[31:0] addr_3943_7;

Selector_2 s3943_7(wires_985_6[3], addr_985_6, addr_positional[15775:15772], addr_3943_7);

wire[31:0] addr_3944_7;

Selector_2 s3944_7(wires_986_6[0], addr_986_6, addr_positional[15779:15776], addr_3944_7);

wire[31:0] addr_3945_7;

Selector_2 s3945_7(wires_986_6[1], addr_986_6, addr_positional[15783:15780], addr_3945_7);

wire[31:0] addr_3946_7;

Selector_2 s3946_7(wires_986_6[2], addr_986_6, addr_positional[15787:15784], addr_3946_7);

wire[31:0] addr_3947_7;

Selector_2 s3947_7(wires_986_6[3], addr_986_6, addr_positional[15791:15788], addr_3947_7);

wire[31:0] addr_3948_7;

Selector_2 s3948_7(wires_987_6[0], addr_987_6, addr_positional[15795:15792], addr_3948_7);

wire[31:0] addr_3949_7;

Selector_2 s3949_7(wires_987_6[1], addr_987_6, addr_positional[15799:15796], addr_3949_7);

wire[31:0] addr_3950_7;

Selector_2 s3950_7(wires_987_6[2], addr_987_6, addr_positional[15803:15800], addr_3950_7);

wire[31:0] addr_3951_7;

Selector_2 s3951_7(wires_987_6[3], addr_987_6, addr_positional[15807:15804], addr_3951_7);

wire[31:0] addr_3952_7;

Selector_2 s3952_7(wires_988_6[0], addr_988_6, addr_positional[15811:15808], addr_3952_7);

wire[31:0] addr_3953_7;

Selector_2 s3953_7(wires_988_6[1], addr_988_6, addr_positional[15815:15812], addr_3953_7);

wire[31:0] addr_3954_7;

Selector_2 s3954_7(wires_988_6[2], addr_988_6, addr_positional[15819:15816], addr_3954_7);

wire[31:0] addr_3955_7;

Selector_2 s3955_7(wires_988_6[3], addr_988_6, addr_positional[15823:15820], addr_3955_7);

wire[31:0] addr_3956_7;

Selector_2 s3956_7(wires_989_6[0], addr_989_6, addr_positional[15827:15824], addr_3956_7);

wire[31:0] addr_3957_7;

Selector_2 s3957_7(wires_989_6[1], addr_989_6, addr_positional[15831:15828], addr_3957_7);

wire[31:0] addr_3958_7;

Selector_2 s3958_7(wires_989_6[2], addr_989_6, addr_positional[15835:15832], addr_3958_7);

wire[31:0] addr_3959_7;

Selector_2 s3959_7(wires_989_6[3], addr_989_6, addr_positional[15839:15836], addr_3959_7);

wire[31:0] addr_3960_7;

Selector_2 s3960_7(wires_990_6[0], addr_990_6, addr_positional[15843:15840], addr_3960_7);

wire[31:0] addr_3961_7;

Selector_2 s3961_7(wires_990_6[1], addr_990_6, addr_positional[15847:15844], addr_3961_7);

wire[31:0] addr_3962_7;

Selector_2 s3962_7(wires_990_6[2], addr_990_6, addr_positional[15851:15848], addr_3962_7);

wire[31:0] addr_3963_7;

Selector_2 s3963_7(wires_990_6[3], addr_990_6, addr_positional[15855:15852], addr_3963_7);

wire[31:0] addr_3964_7;

Selector_2 s3964_7(wires_991_6[0], addr_991_6, addr_positional[15859:15856], addr_3964_7);

wire[31:0] addr_3965_7;

Selector_2 s3965_7(wires_991_6[1], addr_991_6, addr_positional[15863:15860], addr_3965_7);

wire[31:0] addr_3966_7;

Selector_2 s3966_7(wires_991_6[2], addr_991_6, addr_positional[15867:15864], addr_3966_7);

wire[31:0] addr_3967_7;

Selector_2 s3967_7(wires_991_6[3], addr_991_6, addr_positional[15871:15868], addr_3967_7);

wire[31:0] addr_3968_7;

Selector_2 s3968_7(wires_992_6[0], addr_992_6, addr_positional[15875:15872], addr_3968_7);

wire[31:0] addr_3969_7;

Selector_2 s3969_7(wires_992_6[1], addr_992_6, addr_positional[15879:15876], addr_3969_7);

wire[31:0] addr_3970_7;

Selector_2 s3970_7(wires_992_6[2], addr_992_6, addr_positional[15883:15880], addr_3970_7);

wire[31:0] addr_3971_7;

Selector_2 s3971_7(wires_992_6[3], addr_992_6, addr_positional[15887:15884], addr_3971_7);

wire[31:0] addr_3972_7;

Selector_2 s3972_7(wires_993_6[0], addr_993_6, addr_positional[15891:15888], addr_3972_7);

wire[31:0] addr_3973_7;

Selector_2 s3973_7(wires_993_6[1], addr_993_6, addr_positional[15895:15892], addr_3973_7);

wire[31:0] addr_3974_7;

Selector_2 s3974_7(wires_993_6[2], addr_993_6, addr_positional[15899:15896], addr_3974_7);

wire[31:0] addr_3975_7;

Selector_2 s3975_7(wires_993_6[3], addr_993_6, addr_positional[15903:15900], addr_3975_7);

wire[31:0] addr_3976_7;

Selector_2 s3976_7(wires_994_6[0], addr_994_6, addr_positional[15907:15904], addr_3976_7);

wire[31:0] addr_3977_7;

Selector_2 s3977_7(wires_994_6[1], addr_994_6, addr_positional[15911:15908], addr_3977_7);

wire[31:0] addr_3978_7;

Selector_2 s3978_7(wires_994_6[2], addr_994_6, addr_positional[15915:15912], addr_3978_7);

wire[31:0] addr_3979_7;

Selector_2 s3979_7(wires_994_6[3], addr_994_6, addr_positional[15919:15916], addr_3979_7);

wire[31:0] addr_3980_7;

Selector_2 s3980_7(wires_995_6[0], addr_995_6, addr_positional[15923:15920], addr_3980_7);

wire[31:0] addr_3981_7;

Selector_2 s3981_7(wires_995_6[1], addr_995_6, addr_positional[15927:15924], addr_3981_7);

wire[31:0] addr_3982_7;

Selector_2 s3982_7(wires_995_6[2], addr_995_6, addr_positional[15931:15928], addr_3982_7);

wire[31:0] addr_3983_7;

Selector_2 s3983_7(wires_995_6[3], addr_995_6, addr_positional[15935:15932], addr_3983_7);

wire[31:0] addr_3984_7;

Selector_2 s3984_7(wires_996_6[0], addr_996_6, addr_positional[15939:15936], addr_3984_7);

wire[31:0] addr_3985_7;

Selector_2 s3985_7(wires_996_6[1], addr_996_6, addr_positional[15943:15940], addr_3985_7);

wire[31:0] addr_3986_7;

Selector_2 s3986_7(wires_996_6[2], addr_996_6, addr_positional[15947:15944], addr_3986_7);

wire[31:0] addr_3987_7;

Selector_2 s3987_7(wires_996_6[3], addr_996_6, addr_positional[15951:15948], addr_3987_7);

wire[31:0] addr_3988_7;

Selector_2 s3988_7(wires_997_6[0], addr_997_6, addr_positional[15955:15952], addr_3988_7);

wire[31:0] addr_3989_7;

Selector_2 s3989_7(wires_997_6[1], addr_997_6, addr_positional[15959:15956], addr_3989_7);

wire[31:0] addr_3990_7;

Selector_2 s3990_7(wires_997_6[2], addr_997_6, addr_positional[15963:15960], addr_3990_7);

wire[31:0] addr_3991_7;

Selector_2 s3991_7(wires_997_6[3], addr_997_6, addr_positional[15967:15964], addr_3991_7);

wire[31:0] addr_3992_7;

Selector_2 s3992_7(wires_998_6[0], addr_998_6, addr_positional[15971:15968], addr_3992_7);

wire[31:0] addr_3993_7;

Selector_2 s3993_7(wires_998_6[1], addr_998_6, addr_positional[15975:15972], addr_3993_7);

wire[31:0] addr_3994_7;

Selector_2 s3994_7(wires_998_6[2], addr_998_6, addr_positional[15979:15976], addr_3994_7);

wire[31:0] addr_3995_7;

Selector_2 s3995_7(wires_998_6[3], addr_998_6, addr_positional[15983:15980], addr_3995_7);

wire[31:0] addr_3996_7;

Selector_2 s3996_7(wires_999_6[0], addr_999_6, addr_positional[15987:15984], addr_3996_7);

wire[31:0] addr_3997_7;

Selector_2 s3997_7(wires_999_6[1], addr_999_6, addr_positional[15991:15988], addr_3997_7);

wire[31:0] addr_3998_7;

Selector_2 s3998_7(wires_999_6[2], addr_999_6, addr_positional[15995:15992], addr_3998_7);

wire[31:0] addr_3999_7;

Selector_2 s3999_7(wires_999_6[3], addr_999_6, addr_positional[15999:15996], addr_3999_7);

wire[31:0] addr_4000_7;

Selector_2 s4000_7(wires_1000_6[0], addr_1000_6, addr_positional[16003:16000], addr_4000_7);

wire[31:0] addr_4001_7;

Selector_2 s4001_7(wires_1000_6[1], addr_1000_6, addr_positional[16007:16004], addr_4001_7);

wire[31:0] addr_4002_7;

Selector_2 s4002_7(wires_1000_6[2], addr_1000_6, addr_positional[16011:16008], addr_4002_7);

wire[31:0] addr_4003_7;

Selector_2 s4003_7(wires_1000_6[3], addr_1000_6, addr_positional[16015:16012], addr_4003_7);

wire[31:0] addr_4004_7;

Selector_2 s4004_7(wires_1001_6[0], addr_1001_6, addr_positional[16019:16016], addr_4004_7);

wire[31:0] addr_4005_7;

Selector_2 s4005_7(wires_1001_6[1], addr_1001_6, addr_positional[16023:16020], addr_4005_7);

wire[31:0] addr_4006_7;

Selector_2 s4006_7(wires_1001_6[2], addr_1001_6, addr_positional[16027:16024], addr_4006_7);

wire[31:0] addr_4007_7;

Selector_2 s4007_7(wires_1001_6[3], addr_1001_6, addr_positional[16031:16028], addr_4007_7);

wire[31:0] addr_4008_7;

Selector_2 s4008_7(wires_1002_6[0], addr_1002_6, addr_positional[16035:16032], addr_4008_7);

wire[31:0] addr_4009_7;

Selector_2 s4009_7(wires_1002_6[1], addr_1002_6, addr_positional[16039:16036], addr_4009_7);

wire[31:0] addr_4010_7;

Selector_2 s4010_7(wires_1002_6[2], addr_1002_6, addr_positional[16043:16040], addr_4010_7);

wire[31:0] addr_4011_7;

Selector_2 s4011_7(wires_1002_6[3], addr_1002_6, addr_positional[16047:16044], addr_4011_7);

wire[31:0] addr_4012_7;

Selector_2 s4012_7(wires_1003_6[0], addr_1003_6, addr_positional[16051:16048], addr_4012_7);

wire[31:0] addr_4013_7;

Selector_2 s4013_7(wires_1003_6[1], addr_1003_6, addr_positional[16055:16052], addr_4013_7);

wire[31:0] addr_4014_7;

Selector_2 s4014_7(wires_1003_6[2], addr_1003_6, addr_positional[16059:16056], addr_4014_7);

wire[31:0] addr_4015_7;

Selector_2 s4015_7(wires_1003_6[3], addr_1003_6, addr_positional[16063:16060], addr_4015_7);

wire[31:0] addr_4016_7;

Selector_2 s4016_7(wires_1004_6[0], addr_1004_6, addr_positional[16067:16064], addr_4016_7);

wire[31:0] addr_4017_7;

Selector_2 s4017_7(wires_1004_6[1], addr_1004_6, addr_positional[16071:16068], addr_4017_7);

wire[31:0] addr_4018_7;

Selector_2 s4018_7(wires_1004_6[2], addr_1004_6, addr_positional[16075:16072], addr_4018_7);

wire[31:0] addr_4019_7;

Selector_2 s4019_7(wires_1004_6[3], addr_1004_6, addr_positional[16079:16076], addr_4019_7);

wire[31:0] addr_4020_7;

Selector_2 s4020_7(wires_1005_6[0], addr_1005_6, addr_positional[16083:16080], addr_4020_7);

wire[31:0] addr_4021_7;

Selector_2 s4021_7(wires_1005_6[1], addr_1005_6, addr_positional[16087:16084], addr_4021_7);

wire[31:0] addr_4022_7;

Selector_2 s4022_7(wires_1005_6[2], addr_1005_6, addr_positional[16091:16088], addr_4022_7);

wire[31:0] addr_4023_7;

Selector_2 s4023_7(wires_1005_6[3], addr_1005_6, addr_positional[16095:16092], addr_4023_7);

wire[31:0] addr_4024_7;

Selector_2 s4024_7(wires_1006_6[0], addr_1006_6, addr_positional[16099:16096], addr_4024_7);

wire[31:0] addr_4025_7;

Selector_2 s4025_7(wires_1006_6[1], addr_1006_6, addr_positional[16103:16100], addr_4025_7);

wire[31:0] addr_4026_7;

Selector_2 s4026_7(wires_1006_6[2], addr_1006_6, addr_positional[16107:16104], addr_4026_7);

wire[31:0] addr_4027_7;

Selector_2 s4027_7(wires_1006_6[3], addr_1006_6, addr_positional[16111:16108], addr_4027_7);

wire[31:0] addr_4028_7;

Selector_2 s4028_7(wires_1007_6[0], addr_1007_6, addr_positional[16115:16112], addr_4028_7);

wire[31:0] addr_4029_7;

Selector_2 s4029_7(wires_1007_6[1], addr_1007_6, addr_positional[16119:16116], addr_4029_7);

wire[31:0] addr_4030_7;

Selector_2 s4030_7(wires_1007_6[2], addr_1007_6, addr_positional[16123:16120], addr_4030_7);

wire[31:0] addr_4031_7;

Selector_2 s4031_7(wires_1007_6[3], addr_1007_6, addr_positional[16127:16124], addr_4031_7);

wire[31:0] addr_4032_7;

Selector_2 s4032_7(wires_1008_6[0], addr_1008_6, addr_positional[16131:16128], addr_4032_7);

wire[31:0] addr_4033_7;

Selector_2 s4033_7(wires_1008_6[1], addr_1008_6, addr_positional[16135:16132], addr_4033_7);

wire[31:0] addr_4034_7;

Selector_2 s4034_7(wires_1008_6[2], addr_1008_6, addr_positional[16139:16136], addr_4034_7);

wire[31:0] addr_4035_7;

Selector_2 s4035_7(wires_1008_6[3], addr_1008_6, addr_positional[16143:16140], addr_4035_7);

wire[31:0] addr_4036_7;

Selector_2 s4036_7(wires_1009_6[0], addr_1009_6, addr_positional[16147:16144], addr_4036_7);

wire[31:0] addr_4037_7;

Selector_2 s4037_7(wires_1009_6[1], addr_1009_6, addr_positional[16151:16148], addr_4037_7);

wire[31:0] addr_4038_7;

Selector_2 s4038_7(wires_1009_6[2], addr_1009_6, addr_positional[16155:16152], addr_4038_7);

wire[31:0] addr_4039_7;

Selector_2 s4039_7(wires_1009_6[3], addr_1009_6, addr_positional[16159:16156], addr_4039_7);

wire[31:0] addr_4040_7;

Selector_2 s4040_7(wires_1010_6[0], addr_1010_6, addr_positional[16163:16160], addr_4040_7);

wire[31:0] addr_4041_7;

Selector_2 s4041_7(wires_1010_6[1], addr_1010_6, addr_positional[16167:16164], addr_4041_7);

wire[31:0] addr_4042_7;

Selector_2 s4042_7(wires_1010_6[2], addr_1010_6, addr_positional[16171:16168], addr_4042_7);

wire[31:0] addr_4043_7;

Selector_2 s4043_7(wires_1010_6[3], addr_1010_6, addr_positional[16175:16172], addr_4043_7);

wire[31:0] addr_4044_7;

Selector_2 s4044_7(wires_1011_6[0], addr_1011_6, addr_positional[16179:16176], addr_4044_7);

wire[31:0] addr_4045_7;

Selector_2 s4045_7(wires_1011_6[1], addr_1011_6, addr_positional[16183:16180], addr_4045_7);

wire[31:0] addr_4046_7;

Selector_2 s4046_7(wires_1011_6[2], addr_1011_6, addr_positional[16187:16184], addr_4046_7);

wire[31:0] addr_4047_7;

Selector_2 s4047_7(wires_1011_6[3], addr_1011_6, addr_positional[16191:16188], addr_4047_7);

wire[31:0] addr_4048_7;

Selector_2 s4048_7(wires_1012_6[0], addr_1012_6, addr_positional[16195:16192], addr_4048_7);

wire[31:0] addr_4049_7;

Selector_2 s4049_7(wires_1012_6[1], addr_1012_6, addr_positional[16199:16196], addr_4049_7);

wire[31:0] addr_4050_7;

Selector_2 s4050_7(wires_1012_6[2], addr_1012_6, addr_positional[16203:16200], addr_4050_7);

wire[31:0] addr_4051_7;

Selector_2 s4051_7(wires_1012_6[3], addr_1012_6, addr_positional[16207:16204], addr_4051_7);

wire[31:0] addr_4052_7;

Selector_2 s4052_7(wires_1013_6[0], addr_1013_6, addr_positional[16211:16208], addr_4052_7);

wire[31:0] addr_4053_7;

Selector_2 s4053_7(wires_1013_6[1], addr_1013_6, addr_positional[16215:16212], addr_4053_7);

wire[31:0] addr_4054_7;

Selector_2 s4054_7(wires_1013_6[2], addr_1013_6, addr_positional[16219:16216], addr_4054_7);

wire[31:0] addr_4055_7;

Selector_2 s4055_7(wires_1013_6[3], addr_1013_6, addr_positional[16223:16220], addr_4055_7);

wire[31:0] addr_4056_7;

Selector_2 s4056_7(wires_1014_6[0], addr_1014_6, addr_positional[16227:16224], addr_4056_7);

wire[31:0] addr_4057_7;

Selector_2 s4057_7(wires_1014_6[1], addr_1014_6, addr_positional[16231:16228], addr_4057_7);

wire[31:0] addr_4058_7;

Selector_2 s4058_7(wires_1014_6[2], addr_1014_6, addr_positional[16235:16232], addr_4058_7);

wire[31:0] addr_4059_7;

Selector_2 s4059_7(wires_1014_6[3], addr_1014_6, addr_positional[16239:16236], addr_4059_7);

wire[31:0] addr_4060_7;

Selector_2 s4060_7(wires_1015_6[0], addr_1015_6, addr_positional[16243:16240], addr_4060_7);

wire[31:0] addr_4061_7;

Selector_2 s4061_7(wires_1015_6[1], addr_1015_6, addr_positional[16247:16244], addr_4061_7);

wire[31:0] addr_4062_7;

Selector_2 s4062_7(wires_1015_6[2], addr_1015_6, addr_positional[16251:16248], addr_4062_7);

wire[31:0] addr_4063_7;

Selector_2 s4063_7(wires_1015_6[3], addr_1015_6, addr_positional[16255:16252], addr_4063_7);

wire[31:0] addr_4064_7;

Selector_2 s4064_7(wires_1016_6[0], addr_1016_6, addr_positional[16259:16256], addr_4064_7);

wire[31:0] addr_4065_7;

Selector_2 s4065_7(wires_1016_6[1], addr_1016_6, addr_positional[16263:16260], addr_4065_7);

wire[31:0] addr_4066_7;

Selector_2 s4066_7(wires_1016_6[2], addr_1016_6, addr_positional[16267:16264], addr_4066_7);

wire[31:0] addr_4067_7;

Selector_2 s4067_7(wires_1016_6[3], addr_1016_6, addr_positional[16271:16268], addr_4067_7);

wire[31:0] addr_4068_7;

Selector_2 s4068_7(wires_1017_6[0], addr_1017_6, addr_positional[16275:16272], addr_4068_7);

wire[31:0] addr_4069_7;

Selector_2 s4069_7(wires_1017_6[1], addr_1017_6, addr_positional[16279:16276], addr_4069_7);

wire[31:0] addr_4070_7;

Selector_2 s4070_7(wires_1017_6[2], addr_1017_6, addr_positional[16283:16280], addr_4070_7);

wire[31:0] addr_4071_7;

Selector_2 s4071_7(wires_1017_6[3], addr_1017_6, addr_positional[16287:16284], addr_4071_7);

wire[31:0] addr_4072_7;

Selector_2 s4072_7(wires_1018_6[0], addr_1018_6, addr_positional[16291:16288], addr_4072_7);

wire[31:0] addr_4073_7;

Selector_2 s4073_7(wires_1018_6[1], addr_1018_6, addr_positional[16295:16292], addr_4073_7);

wire[31:0] addr_4074_7;

Selector_2 s4074_7(wires_1018_6[2], addr_1018_6, addr_positional[16299:16296], addr_4074_7);

wire[31:0] addr_4075_7;

Selector_2 s4075_7(wires_1018_6[3], addr_1018_6, addr_positional[16303:16300], addr_4075_7);

wire[31:0] addr_4076_7;

Selector_2 s4076_7(wires_1019_6[0], addr_1019_6, addr_positional[16307:16304], addr_4076_7);

wire[31:0] addr_4077_7;

Selector_2 s4077_7(wires_1019_6[1], addr_1019_6, addr_positional[16311:16308], addr_4077_7);

wire[31:0] addr_4078_7;

Selector_2 s4078_7(wires_1019_6[2], addr_1019_6, addr_positional[16315:16312], addr_4078_7);

wire[31:0] addr_4079_7;

Selector_2 s4079_7(wires_1019_6[3], addr_1019_6, addr_positional[16319:16316], addr_4079_7);

wire[31:0] addr_4080_7;

Selector_2 s4080_7(wires_1020_6[0], addr_1020_6, addr_positional[16323:16320], addr_4080_7);

wire[31:0] addr_4081_7;

Selector_2 s4081_7(wires_1020_6[1], addr_1020_6, addr_positional[16327:16324], addr_4081_7);

wire[31:0] addr_4082_7;

Selector_2 s4082_7(wires_1020_6[2], addr_1020_6, addr_positional[16331:16328], addr_4082_7);

wire[31:0] addr_4083_7;

Selector_2 s4083_7(wires_1020_6[3], addr_1020_6, addr_positional[16335:16332], addr_4083_7);

wire[31:0] addr_4084_7;

Selector_2 s4084_7(wires_1021_6[0], addr_1021_6, addr_positional[16339:16336], addr_4084_7);

wire[31:0] addr_4085_7;

Selector_2 s4085_7(wires_1021_6[1], addr_1021_6, addr_positional[16343:16340], addr_4085_7);

wire[31:0] addr_4086_7;

Selector_2 s4086_7(wires_1021_6[2], addr_1021_6, addr_positional[16347:16344], addr_4086_7);

wire[31:0] addr_4087_7;

Selector_2 s4087_7(wires_1021_6[3], addr_1021_6, addr_positional[16351:16348], addr_4087_7);

wire[31:0] addr_4088_7;

Selector_2 s4088_7(wires_1022_6[0], addr_1022_6, addr_positional[16355:16352], addr_4088_7);

wire[31:0] addr_4089_7;

Selector_2 s4089_7(wires_1022_6[1], addr_1022_6, addr_positional[16359:16356], addr_4089_7);

wire[31:0] addr_4090_7;

Selector_2 s4090_7(wires_1022_6[2], addr_1022_6, addr_positional[16363:16360], addr_4090_7);

wire[31:0] addr_4091_7;

Selector_2 s4091_7(wires_1022_6[3], addr_1022_6, addr_positional[16367:16364], addr_4091_7);

wire[31:0] addr_4092_7;

Selector_2 s4092_7(wires_1023_6[0], addr_1023_6, addr_positional[16371:16368], addr_4092_7);

wire[31:0] addr_4093_7;

Selector_2 s4093_7(wires_1023_6[1], addr_1023_6, addr_positional[16375:16372], addr_4093_7);

wire[31:0] addr_4094_7;

Selector_2 s4094_7(wires_1023_6[2], addr_1023_6, addr_positional[16379:16376], addr_4094_7);

wire[31:0] addr_4095_7;

Selector_2 s4095_7(wires_1023_6[3], addr_1023_6, addr_positional[16383:16380], addr_4095_7);

wire[31:0] addr_4096_7;

Selector_2 s4096_7(wires_1024_6[0], addr_1024_6, addr_positional[16387:16384], addr_4096_7);

wire[31:0] addr_4097_7;

Selector_2 s4097_7(wires_1024_6[1], addr_1024_6, addr_positional[16391:16388], addr_4097_7);

wire[31:0] addr_4098_7;

Selector_2 s4098_7(wires_1024_6[2], addr_1024_6, addr_positional[16395:16392], addr_4098_7);

wire[31:0] addr_4099_7;

Selector_2 s4099_7(wires_1024_6[3], addr_1024_6, addr_positional[16399:16396], addr_4099_7);

wire[31:0] addr_4100_7;

Selector_2 s4100_7(wires_1025_6[0], addr_1025_6, addr_positional[16403:16400], addr_4100_7);

wire[31:0] addr_4101_7;

Selector_2 s4101_7(wires_1025_6[1], addr_1025_6, addr_positional[16407:16404], addr_4101_7);

wire[31:0] addr_4102_7;

Selector_2 s4102_7(wires_1025_6[2], addr_1025_6, addr_positional[16411:16408], addr_4102_7);

wire[31:0] addr_4103_7;

Selector_2 s4103_7(wires_1025_6[3], addr_1025_6, addr_positional[16415:16412], addr_4103_7);

wire[31:0] addr_4104_7;

Selector_2 s4104_7(wires_1026_6[0], addr_1026_6, addr_positional[16419:16416], addr_4104_7);

wire[31:0] addr_4105_7;

Selector_2 s4105_7(wires_1026_6[1], addr_1026_6, addr_positional[16423:16420], addr_4105_7);

wire[31:0] addr_4106_7;

Selector_2 s4106_7(wires_1026_6[2], addr_1026_6, addr_positional[16427:16424], addr_4106_7);

wire[31:0] addr_4107_7;

Selector_2 s4107_7(wires_1026_6[3], addr_1026_6, addr_positional[16431:16428], addr_4107_7);

wire[31:0] addr_4108_7;

Selector_2 s4108_7(wires_1027_6[0], addr_1027_6, addr_positional[16435:16432], addr_4108_7);

wire[31:0] addr_4109_7;

Selector_2 s4109_7(wires_1027_6[1], addr_1027_6, addr_positional[16439:16436], addr_4109_7);

wire[31:0] addr_4110_7;

Selector_2 s4110_7(wires_1027_6[2], addr_1027_6, addr_positional[16443:16440], addr_4110_7);

wire[31:0] addr_4111_7;

Selector_2 s4111_7(wires_1027_6[3], addr_1027_6, addr_positional[16447:16444], addr_4111_7);

wire[31:0] addr_4112_7;

Selector_2 s4112_7(wires_1028_6[0], addr_1028_6, addr_positional[16451:16448], addr_4112_7);

wire[31:0] addr_4113_7;

Selector_2 s4113_7(wires_1028_6[1], addr_1028_6, addr_positional[16455:16452], addr_4113_7);

wire[31:0] addr_4114_7;

Selector_2 s4114_7(wires_1028_6[2], addr_1028_6, addr_positional[16459:16456], addr_4114_7);

wire[31:0] addr_4115_7;

Selector_2 s4115_7(wires_1028_6[3], addr_1028_6, addr_positional[16463:16460], addr_4115_7);

wire[31:0] addr_4116_7;

Selector_2 s4116_7(wires_1029_6[0], addr_1029_6, addr_positional[16467:16464], addr_4116_7);

wire[31:0] addr_4117_7;

Selector_2 s4117_7(wires_1029_6[1], addr_1029_6, addr_positional[16471:16468], addr_4117_7);

wire[31:0] addr_4118_7;

Selector_2 s4118_7(wires_1029_6[2], addr_1029_6, addr_positional[16475:16472], addr_4118_7);

wire[31:0] addr_4119_7;

Selector_2 s4119_7(wires_1029_6[3], addr_1029_6, addr_positional[16479:16476], addr_4119_7);

wire[31:0] addr_4120_7;

Selector_2 s4120_7(wires_1030_6[0], addr_1030_6, addr_positional[16483:16480], addr_4120_7);

wire[31:0] addr_4121_7;

Selector_2 s4121_7(wires_1030_6[1], addr_1030_6, addr_positional[16487:16484], addr_4121_7);

wire[31:0] addr_4122_7;

Selector_2 s4122_7(wires_1030_6[2], addr_1030_6, addr_positional[16491:16488], addr_4122_7);

wire[31:0] addr_4123_7;

Selector_2 s4123_7(wires_1030_6[3], addr_1030_6, addr_positional[16495:16492], addr_4123_7);

wire[31:0] addr_4124_7;

Selector_2 s4124_7(wires_1031_6[0], addr_1031_6, addr_positional[16499:16496], addr_4124_7);

wire[31:0] addr_4125_7;

Selector_2 s4125_7(wires_1031_6[1], addr_1031_6, addr_positional[16503:16500], addr_4125_7);

wire[31:0] addr_4126_7;

Selector_2 s4126_7(wires_1031_6[2], addr_1031_6, addr_positional[16507:16504], addr_4126_7);

wire[31:0] addr_4127_7;

Selector_2 s4127_7(wires_1031_6[3], addr_1031_6, addr_positional[16511:16508], addr_4127_7);

wire[31:0] addr_4128_7;

Selector_2 s4128_7(wires_1032_6[0], addr_1032_6, addr_positional[16515:16512], addr_4128_7);

wire[31:0] addr_4129_7;

Selector_2 s4129_7(wires_1032_6[1], addr_1032_6, addr_positional[16519:16516], addr_4129_7);

wire[31:0] addr_4130_7;

Selector_2 s4130_7(wires_1032_6[2], addr_1032_6, addr_positional[16523:16520], addr_4130_7);

wire[31:0] addr_4131_7;

Selector_2 s4131_7(wires_1032_6[3], addr_1032_6, addr_positional[16527:16524], addr_4131_7);

wire[31:0] addr_4132_7;

Selector_2 s4132_7(wires_1033_6[0], addr_1033_6, addr_positional[16531:16528], addr_4132_7);

wire[31:0] addr_4133_7;

Selector_2 s4133_7(wires_1033_6[1], addr_1033_6, addr_positional[16535:16532], addr_4133_7);

wire[31:0] addr_4134_7;

Selector_2 s4134_7(wires_1033_6[2], addr_1033_6, addr_positional[16539:16536], addr_4134_7);

wire[31:0] addr_4135_7;

Selector_2 s4135_7(wires_1033_6[3], addr_1033_6, addr_positional[16543:16540], addr_4135_7);

wire[31:0] addr_4136_7;

Selector_2 s4136_7(wires_1034_6[0], addr_1034_6, addr_positional[16547:16544], addr_4136_7);

wire[31:0] addr_4137_7;

Selector_2 s4137_7(wires_1034_6[1], addr_1034_6, addr_positional[16551:16548], addr_4137_7);

wire[31:0] addr_4138_7;

Selector_2 s4138_7(wires_1034_6[2], addr_1034_6, addr_positional[16555:16552], addr_4138_7);

wire[31:0] addr_4139_7;

Selector_2 s4139_7(wires_1034_6[3], addr_1034_6, addr_positional[16559:16556], addr_4139_7);

wire[31:0] addr_4140_7;

Selector_2 s4140_7(wires_1035_6[0], addr_1035_6, addr_positional[16563:16560], addr_4140_7);

wire[31:0] addr_4141_7;

Selector_2 s4141_7(wires_1035_6[1], addr_1035_6, addr_positional[16567:16564], addr_4141_7);

wire[31:0] addr_4142_7;

Selector_2 s4142_7(wires_1035_6[2], addr_1035_6, addr_positional[16571:16568], addr_4142_7);

wire[31:0] addr_4143_7;

Selector_2 s4143_7(wires_1035_6[3], addr_1035_6, addr_positional[16575:16572], addr_4143_7);

wire[31:0] addr_4144_7;

Selector_2 s4144_7(wires_1036_6[0], addr_1036_6, addr_positional[16579:16576], addr_4144_7);

wire[31:0] addr_4145_7;

Selector_2 s4145_7(wires_1036_6[1], addr_1036_6, addr_positional[16583:16580], addr_4145_7);

wire[31:0] addr_4146_7;

Selector_2 s4146_7(wires_1036_6[2], addr_1036_6, addr_positional[16587:16584], addr_4146_7);

wire[31:0] addr_4147_7;

Selector_2 s4147_7(wires_1036_6[3], addr_1036_6, addr_positional[16591:16588], addr_4147_7);

wire[31:0] addr_4148_7;

Selector_2 s4148_7(wires_1037_6[0], addr_1037_6, addr_positional[16595:16592], addr_4148_7);

wire[31:0] addr_4149_7;

Selector_2 s4149_7(wires_1037_6[1], addr_1037_6, addr_positional[16599:16596], addr_4149_7);

wire[31:0] addr_4150_7;

Selector_2 s4150_7(wires_1037_6[2], addr_1037_6, addr_positional[16603:16600], addr_4150_7);

wire[31:0] addr_4151_7;

Selector_2 s4151_7(wires_1037_6[3], addr_1037_6, addr_positional[16607:16604], addr_4151_7);

wire[31:0] addr_4152_7;

Selector_2 s4152_7(wires_1038_6[0], addr_1038_6, addr_positional[16611:16608], addr_4152_7);

wire[31:0] addr_4153_7;

Selector_2 s4153_7(wires_1038_6[1], addr_1038_6, addr_positional[16615:16612], addr_4153_7);

wire[31:0] addr_4154_7;

Selector_2 s4154_7(wires_1038_6[2], addr_1038_6, addr_positional[16619:16616], addr_4154_7);

wire[31:0] addr_4155_7;

Selector_2 s4155_7(wires_1038_6[3], addr_1038_6, addr_positional[16623:16620], addr_4155_7);

wire[31:0] addr_4156_7;

Selector_2 s4156_7(wires_1039_6[0], addr_1039_6, addr_positional[16627:16624], addr_4156_7);

wire[31:0] addr_4157_7;

Selector_2 s4157_7(wires_1039_6[1], addr_1039_6, addr_positional[16631:16628], addr_4157_7);

wire[31:0] addr_4158_7;

Selector_2 s4158_7(wires_1039_6[2], addr_1039_6, addr_positional[16635:16632], addr_4158_7);

wire[31:0] addr_4159_7;

Selector_2 s4159_7(wires_1039_6[3], addr_1039_6, addr_positional[16639:16636], addr_4159_7);

wire[31:0] addr_4160_7;

Selector_2 s4160_7(wires_1040_6[0], addr_1040_6, addr_positional[16643:16640], addr_4160_7);

wire[31:0] addr_4161_7;

Selector_2 s4161_7(wires_1040_6[1], addr_1040_6, addr_positional[16647:16644], addr_4161_7);

wire[31:0] addr_4162_7;

Selector_2 s4162_7(wires_1040_6[2], addr_1040_6, addr_positional[16651:16648], addr_4162_7);

wire[31:0] addr_4163_7;

Selector_2 s4163_7(wires_1040_6[3], addr_1040_6, addr_positional[16655:16652], addr_4163_7);

wire[31:0] addr_4164_7;

Selector_2 s4164_7(wires_1041_6[0], addr_1041_6, addr_positional[16659:16656], addr_4164_7);

wire[31:0] addr_4165_7;

Selector_2 s4165_7(wires_1041_6[1], addr_1041_6, addr_positional[16663:16660], addr_4165_7);

wire[31:0] addr_4166_7;

Selector_2 s4166_7(wires_1041_6[2], addr_1041_6, addr_positional[16667:16664], addr_4166_7);

wire[31:0] addr_4167_7;

Selector_2 s4167_7(wires_1041_6[3], addr_1041_6, addr_positional[16671:16668], addr_4167_7);

wire[31:0] addr_4168_7;

Selector_2 s4168_7(wires_1042_6[0], addr_1042_6, addr_positional[16675:16672], addr_4168_7);

wire[31:0] addr_4169_7;

Selector_2 s4169_7(wires_1042_6[1], addr_1042_6, addr_positional[16679:16676], addr_4169_7);

wire[31:0] addr_4170_7;

Selector_2 s4170_7(wires_1042_6[2], addr_1042_6, addr_positional[16683:16680], addr_4170_7);

wire[31:0] addr_4171_7;

Selector_2 s4171_7(wires_1042_6[3], addr_1042_6, addr_positional[16687:16684], addr_4171_7);

wire[31:0] addr_4172_7;

Selector_2 s4172_7(wires_1043_6[0], addr_1043_6, addr_positional[16691:16688], addr_4172_7);

wire[31:0] addr_4173_7;

Selector_2 s4173_7(wires_1043_6[1], addr_1043_6, addr_positional[16695:16692], addr_4173_7);

wire[31:0] addr_4174_7;

Selector_2 s4174_7(wires_1043_6[2], addr_1043_6, addr_positional[16699:16696], addr_4174_7);

wire[31:0] addr_4175_7;

Selector_2 s4175_7(wires_1043_6[3], addr_1043_6, addr_positional[16703:16700], addr_4175_7);

wire[31:0] addr_4176_7;

Selector_2 s4176_7(wires_1044_6[0], addr_1044_6, addr_positional[16707:16704], addr_4176_7);

wire[31:0] addr_4177_7;

Selector_2 s4177_7(wires_1044_6[1], addr_1044_6, addr_positional[16711:16708], addr_4177_7);

wire[31:0] addr_4178_7;

Selector_2 s4178_7(wires_1044_6[2], addr_1044_6, addr_positional[16715:16712], addr_4178_7);

wire[31:0] addr_4179_7;

Selector_2 s4179_7(wires_1044_6[3], addr_1044_6, addr_positional[16719:16716], addr_4179_7);

wire[31:0] addr_4180_7;

Selector_2 s4180_7(wires_1045_6[0], addr_1045_6, addr_positional[16723:16720], addr_4180_7);

wire[31:0] addr_4181_7;

Selector_2 s4181_7(wires_1045_6[1], addr_1045_6, addr_positional[16727:16724], addr_4181_7);

wire[31:0] addr_4182_7;

Selector_2 s4182_7(wires_1045_6[2], addr_1045_6, addr_positional[16731:16728], addr_4182_7);

wire[31:0] addr_4183_7;

Selector_2 s4183_7(wires_1045_6[3], addr_1045_6, addr_positional[16735:16732], addr_4183_7);

wire[31:0] addr_4184_7;

Selector_2 s4184_7(wires_1046_6[0], addr_1046_6, addr_positional[16739:16736], addr_4184_7);

wire[31:0] addr_4185_7;

Selector_2 s4185_7(wires_1046_6[1], addr_1046_6, addr_positional[16743:16740], addr_4185_7);

wire[31:0] addr_4186_7;

Selector_2 s4186_7(wires_1046_6[2], addr_1046_6, addr_positional[16747:16744], addr_4186_7);

wire[31:0] addr_4187_7;

Selector_2 s4187_7(wires_1046_6[3], addr_1046_6, addr_positional[16751:16748], addr_4187_7);

wire[31:0] addr_4188_7;

Selector_2 s4188_7(wires_1047_6[0], addr_1047_6, addr_positional[16755:16752], addr_4188_7);

wire[31:0] addr_4189_7;

Selector_2 s4189_7(wires_1047_6[1], addr_1047_6, addr_positional[16759:16756], addr_4189_7);

wire[31:0] addr_4190_7;

Selector_2 s4190_7(wires_1047_6[2], addr_1047_6, addr_positional[16763:16760], addr_4190_7);

wire[31:0] addr_4191_7;

Selector_2 s4191_7(wires_1047_6[3], addr_1047_6, addr_positional[16767:16764], addr_4191_7);

wire[31:0] addr_4192_7;

Selector_2 s4192_7(wires_1048_6[0], addr_1048_6, addr_positional[16771:16768], addr_4192_7);

wire[31:0] addr_4193_7;

Selector_2 s4193_7(wires_1048_6[1], addr_1048_6, addr_positional[16775:16772], addr_4193_7);

wire[31:0] addr_4194_7;

Selector_2 s4194_7(wires_1048_6[2], addr_1048_6, addr_positional[16779:16776], addr_4194_7);

wire[31:0] addr_4195_7;

Selector_2 s4195_7(wires_1048_6[3], addr_1048_6, addr_positional[16783:16780], addr_4195_7);

wire[31:0] addr_4196_7;

Selector_2 s4196_7(wires_1049_6[0], addr_1049_6, addr_positional[16787:16784], addr_4196_7);

wire[31:0] addr_4197_7;

Selector_2 s4197_7(wires_1049_6[1], addr_1049_6, addr_positional[16791:16788], addr_4197_7);

wire[31:0] addr_4198_7;

Selector_2 s4198_7(wires_1049_6[2], addr_1049_6, addr_positional[16795:16792], addr_4198_7);

wire[31:0] addr_4199_7;

Selector_2 s4199_7(wires_1049_6[3], addr_1049_6, addr_positional[16799:16796], addr_4199_7);

wire[31:0] addr_4200_7;

Selector_2 s4200_7(wires_1050_6[0], addr_1050_6, addr_positional[16803:16800], addr_4200_7);

wire[31:0] addr_4201_7;

Selector_2 s4201_7(wires_1050_6[1], addr_1050_6, addr_positional[16807:16804], addr_4201_7);

wire[31:0] addr_4202_7;

Selector_2 s4202_7(wires_1050_6[2], addr_1050_6, addr_positional[16811:16808], addr_4202_7);

wire[31:0] addr_4203_7;

Selector_2 s4203_7(wires_1050_6[3], addr_1050_6, addr_positional[16815:16812], addr_4203_7);

wire[31:0] addr_4204_7;

Selector_2 s4204_7(wires_1051_6[0], addr_1051_6, addr_positional[16819:16816], addr_4204_7);

wire[31:0] addr_4205_7;

Selector_2 s4205_7(wires_1051_6[1], addr_1051_6, addr_positional[16823:16820], addr_4205_7);

wire[31:0] addr_4206_7;

Selector_2 s4206_7(wires_1051_6[2], addr_1051_6, addr_positional[16827:16824], addr_4206_7);

wire[31:0] addr_4207_7;

Selector_2 s4207_7(wires_1051_6[3], addr_1051_6, addr_positional[16831:16828], addr_4207_7);

wire[31:0] addr_4208_7;

Selector_2 s4208_7(wires_1052_6[0], addr_1052_6, addr_positional[16835:16832], addr_4208_7);

wire[31:0] addr_4209_7;

Selector_2 s4209_7(wires_1052_6[1], addr_1052_6, addr_positional[16839:16836], addr_4209_7);

wire[31:0] addr_4210_7;

Selector_2 s4210_7(wires_1052_6[2], addr_1052_6, addr_positional[16843:16840], addr_4210_7);

wire[31:0] addr_4211_7;

Selector_2 s4211_7(wires_1052_6[3], addr_1052_6, addr_positional[16847:16844], addr_4211_7);

wire[31:0] addr_4212_7;

Selector_2 s4212_7(wires_1053_6[0], addr_1053_6, addr_positional[16851:16848], addr_4212_7);

wire[31:0] addr_4213_7;

Selector_2 s4213_7(wires_1053_6[1], addr_1053_6, addr_positional[16855:16852], addr_4213_7);

wire[31:0] addr_4214_7;

Selector_2 s4214_7(wires_1053_6[2], addr_1053_6, addr_positional[16859:16856], addr_4214_7);

wire[31:0] addr_4215_7;

Selector_2 s4215_7(wires_1053_6[3], addr_1053_6, addr_positional[16863:16860], addr_4215_7);

wire[31:0] addr_4216_7;

Selector_2 s4216_7(wires_1054_6[0], addr_1054_6, addr_positional[16867:16864], addr_4216_7);

wire[31:0] addr_4217_7;

Selector_2 s4217_7(wires_1054_6[1], addr_1054_6, addr_positional[16871:16868], addr_4217_7);

wire[31:0] addr_4218_7;

Selector_2 s4218_7(wires_1054_6[2], addr_1054_6, addr_positional[16875:16872], addr_4218_7);

wire[31:0] addr_4219_7;

Selector_2 s4219_7(wires_1054_6[3], addr_1054_6, addr_positional[16879:16876], addr_4219_7);

wire[31:0] addr_4220_7;

Selector_2 s4220_7(wires_1055_6[0], addr_1055_6, addr_positional[16883:16880], addr_4220_7);

wire[31:0] addr_4221_7;

Selector_2 s4221_7(wires_1055_6[1], addr_1055_6, addr_positional[16887:16884], addr_4221_7);

wire[31:0] addr_4222_7;

Selector_2 s4222_7(wires_1055_6[2], addr_1055_6, addr_positional[16891:16888], addr_4222_7);

wire[31:0] addr_4223_7;

Selector_2 s4223_7(wires_1055_6[3], addr_1055_6, addr_positional[16895:16892], addr_4223_7);

wire[31:0] addr_4224_7;

Selector_2 s4224_7(wires_1056_6[0], addr_1056_6, addr_positional[16899:16896], addr_4224_7);

wire[31:0] addr_4225_7;

Selector_2 s4225_7(wires_1056_6[1], addr_1056_6, addr_positional[16903:16900], addr_4225_7);

wire[31:0] addr_4226_7;

Selector_2 s4226_7(wires_1056_6[2], addr_1056_6, addr_positional[16907:16904], addr_4226_7);

wire[31:0] addr_4227_7;

Selector_2 s4227_7(wires_1056_6[3], addr_1056_6, addr_positional[16911:16908], addr_4227_7);

wire[31:0] addr_4228_7;

Selector_2 s4228_7(wires_1057_6[0], addr_1057_6, addr_positional[16915:16912], addr_4228_7);

wire[31:0] addr_4229_7;

Selector_2 s4229_7(wires_1057_6[1], addr_1057_6, addr_positional[16919:16916], addr_4229_7);

wire[31:0] addr_4230_7;

Selector_2 s4230_7(wires_1057_6[2], addr_1057_6, addr_positional[16923:16920], addr_4230_7);

wire[31:0] addr_4231_7;

Selector_2 s4231_7(wires_1057_6[3], addr_1057_6, addr_positional[16927:16924], addr_4231_7);

wire[31:0] addr_4232_7;

Selector_2 s4232_7(wires_1058_6[0], addr_1058_6, addr_positional[16931:16928], addr_4232_7);

wire[31:0] addr_4233_7;

Selector_2 s4233_7(wires_1058_6[1], addr_1058_6, addr_positional[16935:16932], addr_4233_7);

wire[31:0] addr_4234_7;

Selector_2 s4234_7(wires_1058_6[2], addr_1058_6, addr_positional[16939:16936], addr_4234_7);

wire[31:0] addr_4235_7;

Selector_2 s4235_7(wires_1058_6[3], addr_1058_6, addr_positional[16943:16940], addr_4235_7);

wire[31:0] addr_4236_7;

Selector_2 s4236_7(wires_1059_6[0], addr_1059_6, addr_positional[16947:16944], addr_4236_7);

wire[31:0] addr_4237_7;

Selector_2 s4237_7(wires_1059_6[1], addr_1059_6, addr_positional[16951:16948], addr_4237_7);

wire[31:0] addr_4238_7;

Selector_2 s4238_7(wires_1059_6[2], addr_1059_6, addr_positional[16955:16952], addr_4238_7);

wire[31:0] addr_4239_7;

Selector_2 s4239_7(wires_1059_6[3], addr_1059_6, addr_positional[16959:16956], addr_4239_7);

wire[31:0] addr_4240_7;

Selector_2 s4240_7(wires_1060_6[0], addr_1060_6, addr_positional[16963:16960], addr_4240_7);

wire[31:0] addr_4241_7;

Selector_2 s4241_7(wires_1060_6[1], addr_1060_6, addr_positional[16967:16964], addr_4241_7);

wire[31:0] addr_4242_7;

Selector_2 s4242_7(wires_1060_6[2], addr_1060_6, addr_positional[16971:16968], addr_4242_7);

wire[31:0] addr_4243_7;

Selector_2 s4243_7(wires_1060_6[3], addr_1060_6, addr_positional[16975:16972], addr_4243_7);

wire[31:0] addr_4244_7;

Selector_2 s4244_7(wires_1061_6[0], addr_1061_6, addr_positional[16979:16976], addr_4244_7);

wire[31:0] addr_4245_7;

Selector_2 s4245_7(wires_1061_6[1], addr_1061_6, addr_positional[16983:16980], addr_4245_7);

wire[31:0] addr_4246_7;

Selector_2 s4246_7(wires_1061_6[2], addr_1061_6, addr_positional[16987:16984], addr_4246_7);

wire[31:0] addr_4247_7;

Selector_2 s4247_7(wires_1061_6[3], addr_1061_6, addr_positional[16991:16988], addr_4247_7);

wire[31:0] addr_4248_7;

Selector_2 s4248_7(wires_1062_6[0], addr_1062_6, addr_positional[16995:16992], addr_4248_7);

wire[31:0] addr_4249_7;

Selector_2 s4249_7(wires_1062_6[1], addr_1062_6, addr_positional[16999:16996], addr_4249_7);

wire[31:0] addr_4250_7;

Selector_2 s4250_7(wires_1062_6[2], addr_1062_6, addr_positional[17003:17000], addr_4250_7);

wire[31:0] addr_4251_7;

Selector_2 s4251_7(wires_1062_6[3], addr_1062_6, addr_positional[17007:17004], addr_4251_7);

wire[31:0] addr_4252_7;

Selector_2 s4252_7(wires_1063_6[0], addr_1063_6, addr_positional[17011:17008], addr_4252_7);

wire[31:0] addr_4253_7;

Selector_2 s4253_7(wires_1063_6[1], addr_1063_6, addr_positional[17015:17012], addr_4253_7);

wire[31:0] addr_4254_7;

Selector_2 s4254_7(wires_1063_6[2], addr_1063_6, addr_positional[17019:17016], addr_4254_7);

wire[31:0] addr_4255_7;

Selector_2 s4255_7(wires_1063_6[3], addr_1063_6, addr_positional[17023:17020], addr_4255_7);

wire[31:0] addr_4256_7;

Selector_2 s4256_7(wires_1064_6[0], addr_1064_6, addr_positional[17027:17024], addr_4256_7);

wire[31:0] addr_4257_7;

Selector_2 s4257_7(wires_1064_6[1], addr_1064_6, addr_positional[17031:17028], addr_4257_7);

wire[31:0] addr_4258_7;

Selector_2 s4258_7(wires_1064_6[2], addr_1064_6, addr_positional[17035:17032], addr_4258_7);

wire[31:0] addr_4259_7;

Selector_2 s4259_7(wires_1064_6[3], addr_1064_6, addr_positional[17039:17036], addr_4259_7);

wire[31:0] addr_4260_7;

Selector_2 s4260_7(wires_1065_6[0], addr_1065_6, addr_positional[17043:17040], addr_4260_7);

wire[31:0] addr_4261_7;

Selector_2 s4261_7(wires_1065_6[1], addr_1065_6, addr_positional[17047:17044], addr_4261_7);

wire[31:0] addr_4262_7;

Selector_2 s4262_7(wires_1065_6[2], addr_1065_6, addr_positional[17051:17048], addr_4262_7);

wire[31:0] addr_4263_7;

Selector_2 s4263_7(wires_1065_6[3], addr_1065_6, addr_positional[17055:17052], addr_4263_7);

wire[31:0] addr_4264_7;

Selector_2 s4264_7(wires_1066_6[0], addr_1066_6, addr_positional[17059:17056], addr_4264_7);

wire[31:0] addr_4265_7;

Selector_2 s4265_7(wires_1066_6[1], addr_1066_6, addr_positional[17063:17060], addr_4265_7);

wire[31:0] addr_4266_7;

Selector_2 s4266_7(wires_1066_6[2], addr_1066_6, addr_positional[17067:17064], addr_4266_7);

wire[31:0] addr_4267_7;

Selector_2 s4267_7(wires_1066_6[3], addr_1066_6, addr_positional[17071:17068], addr_4267_7);

wire[31:0] addr_4268_7;

Selector_2 s4268_7(wires_1067_6[0], addr_1067_6, addr_positional[17075:17072], addr_4268_7);

wire[31:0] addr_4269_7;

Selector_2 s4269_7(wires_1067_6[1], addr_1067_6, addr_positional[17079:17076], addr_4269_7);

wire[31:0] addr_4270_7;

Selector_2 s4270_7(wires_1067_6[2], addr_1067_6, addr_positional[17083:17080], addr_4270_7);

wire[31:0] addr_4271_7;

Selector_2 s4271_7(wires_1067_6[3], addr_1067_6, addr_positional[17087:17084], addr_4271_7);

wire[31:0] addr_4272_7;

Selector_2 s4272_7(wires_1068_6[0], addr_1068_6, addr_positional[17091:17088], addr_4272_7);

wire[31:0] addr_4273_7;

Selector_2 s4273_7(wires_1068_6[1], addr_1068_6, addr_positional[17095:17092], addr_4273_7);

wire[31:0] addr_4274_7;

Selector_2 s4274_7(wires_1068_6[2], addr_1068_6, addr_positional[17099:17096], addr_4274_7);

wire[31:0] addr_4275_7;

Selector_2 s4275_7(wires_1068_6[3], addr_1068_6, addr_positional[17103:17100], addr_4275_7);

wire[31:0] addr_4276_7;

Selector_2 s4276_7(wires_1069_6[0], addr_1069_6, addr_positional[17107:17104], addr_4276_7);

wire[31:0] addr_4277_7;

Selector_2 s4277_7(wires_1069_6[1], addr_1069_6, addr_positional[17111:17108], addr_4277_7);

wire[31:0] addr_4278_7;

Selector_2 s4278_7(wires_1069_6[2], addr_1069_6, addr_positional[17115:17112], addr_4278_7);

wire[31:0] addr_4279_7;

Selector_2 s4279_7(wires_1069_6[3], addr_1069_6, addr_positional[17119:17116], addr_4279_7);

wire[31:0] addr_4280_7;

Selector_2 s4280_7(wires_1070_6[0], addr_1070_6, addr_positional[17123:17120], addr_4280_7);

wire[31:0] addr_4281_7;

Selector_2 s4281_7(wires_1070_6[1], addr_1070_6, addr_positional[17127:17124], addr_4281_7);

wire[31:0] addr_4282_7;

Selector_2 s4282_7(wires_1070_6[2], addr_1070_6, addr_positional[17131:17128], addr_4282_7);

wire[31:0] addr_4283_7;

Selector_2 s4283_7(wires_1070_6[3], addr_1070_6, addr_positional[17135:17132], addr_4283_7);

wire[31:0] addr_4284_7;

Selector_2 s4284_7(wires_1071_6[0], addr_1071_6, addr_positional[17139:17136], addr_4284_7);

wire[31:0] addr_4285_7;

Selector_2 s4285_7(wires_1071_6[1], addr_1071_6, addr_positional[17143:17140], addr_4285_7);

wire[31:0] addr_4286_7;

Selector_2 s4286_7(wires_1071_6[2], addr_1071_6, addr_positional[17147:17144], addr_4286_7);

wire[31:0] addr_4287_7;

Selector_2 s4287_7(wires_1071_6[3], addr_1071_6, addr_positional[17151:17148], addr_4287_7);

wire[31:0] addr_4288_7;

Selector_2 s4288_7(wires_1072_6[0], addr_1072_6, addr_positional[17155:17152], addr_4288_7);

wire[31:0] addr_4289_7;

Selector_2 s4289_7(wires_1072_6[1], addr_1072_6, addr_positional[17159:17156], addr_4289_7);

wire[31:0] addr_4290_7;

Selector_2 s4290_7(wires_1072_6[2], addr_1072_6, addr_positional[17163:17160], addr_4290_7);

wire[31:0] addr_4291_7;

Selector_2 s4291_7(wires_1072_6[3], addr_1072_6, addr_positional[17167:17164], addr_4291_7);

wire[31:0] addr_4292_7;

Selector_2 s4292_7(wires_1073_6[0], addr_1073_6, addr_positional[17171:17168], addr_4292_7);

wire[31:0] addr_4293_7;

Selector_2 s4293_7(wires_1073_6[1], addr_1073_6, addr_positional[17175:17172], addr_4293_7);

wire[31:0] addr_4294_7;

Selector_2 s4294_7(wires_1073_6[2], addr_1073_6, addr_positional[17179:17176], addr_4294_7);

wire[31:0] addr_4295_7;

Selector_2 s4295_7(wires_1073_6[3], addr_1073_6, addr_positional[17183:17180], addr_4295_7);

wire[31:0] addr_4296_7;

Selector_2 s4296_7(wires_1074_6[0], addr_1074_6, addr_positional[17187:17184], addr_4296_7);

wire[31:0] addr_4297_7;

Selector_2 s4297_7(wires_1074_6[1], addr_1074_6, addr_positional[17191:17188], addr_4297_7);

wire[31:0] addr_4298_7;

Selector_2 s4298_7(wires_1074_6[2], addr_1074_6, addr_positional[17195:17192], addr_4298_7);

wire[31:0] addr_4299_7;

Selector_2 s4299_7(wires_1074_6[3], addr_1074_6, addr_positional[17199:17196], addr_4299_7);

wire[31:0] addr_4300_7;

Selector_2 s4300_7(wires_1075_6[0], addr_1075_6, addr_positional[17203:17200], addr_4300_7);

wire[31:0] addr_4301_7;

Selector_2 s4301_7(wires_1075_6[1], addr_1075_6, addr_positional[17207:17204], addr_4301_7);

wire[31:0] addr_4302_7;

Selector_2 s4302_7(wires_1075_6[2], addr_1075_6, addr_positional[17211:17208], addr_4302_7);

wire[31:0] addr_4303_7;

Selector_2 s4303_7(wires_1075_6[3], addr_1075_6, addr_positional[17215:17212], addr_4303_7);

wire[31:0] addr_4304_7;

Selector_2 s4304_7(wires_1076_6[0], addr_1076_6, addr_positional[17219:17216], addr_4304_7);

wire[31:0] addr_4305_7;

Selector_2 s4305_7(wires_1076_6[1], addr_1076_6, addr_positional[17223:17220], addr_4305_7);

wire[31:0] addr_4306_7;

Selector_2 s4306_7(wires_1076_6[2], addr_1076_6, addr_positional[17227:17224], addr_4306_7);

wire[31:0] addr_4307_7;

Selector_2 s4307_7(wires_1076_6[3], addr_1076_6, addr_positional[17231:17228], addr_4307_7);

wire[31:0] addr_4308_7;

Selector_2 s4308_7(wires_1077_6[0], addr_1077_6, addr_positional[17235:17232], addr_4308_7);

wire[31:0] addr_4309_7;

Selector_2 s4309_7(wires_1077_6[1], addr_1077_6, addr_positional[17239:17236], addr_4309_7);

wire[31:0] addr_4310_7;

Selector_2 s4310_7(wires_1077_6[2], addr_1077_6, addr_positional[17243:17240], addr_4310_7);

wire[31:0] addr_4311_7;

Selector_2 s4311_7(wires_1077_6[3], addr_1077_6, addr_positional[17247:17244], addr_4311_7);

wire[31:0] addr_4312_7;

Selector_2 s4312_7(wires_1078_6[0], addr_1078_6, addr_positional[17251:17248], addr_4312_7);

wire[31:0] addr_4313_7;

Selector_2 s4313_7(wires_1078_6[1], addr_1078_6, addr_positional[17255:17252], addr_4313_7);

wire[31:0] addr_4314_7;

Selector_2 s4314_7(wires_1078_6[2], addr_1078_6, addr_positional[17259:17256], addr_4314_7);

wire[31:0] addr_4315_7;

Selector_2 s4315_7(wires_1078_6[3], addr_1078_6, addr_positional[17263:17260], addr_4315_7);

wire[31:0] addr_4316_7;

Selector_2 s4316_7(wires_1079_6[0], addr_1079_6, addr_positional[17267:17264], addr_4316_7);

wire[31:0] addr_4317_7;

Selector_2 s4317_7(wires_1079_6[1], addr_1079_6, addr_positional[17271:17268], addr_4317_7);

wire[31:0] addr_4318_7;

Selector_2 s4318_7(wires_1079_6[2], addr_1079_6, addr_positional[17275:17272], addr_4318_7);

wire[31:0] addr_4319_7;

Selector_2 s4319_7(wires_1079_6[3], addr_1079_6, addr_positional[17279:17276], addr_4319_7);

wire[31:0] addr_4320_7;

Selector_2 s4320_7(wires_1080_6[0], addr_1080_6, addr_positional[17283:17280], addr_4320_7);

wire[31:0] addr_4321_7;

Selector_2 s4321_7(wires_1080_6[1], addr_1080_6, addr_positional[17287:17284], addr_4321_7);

wire[31:0] addr_4322_7;

Selector_2 s4322_7(wires_1080_6[2], addr_1080_6, addr_positional[17291:17288], addr_4322_7);

wire[31:0] addr_4323_7;

Selector_2 s4323_7(wires_1080_6[3], addr_1080_6, addr_positional[17295:17292], addr_4323_7);

wire[31:0] addr_4324_7;

Selector_2 s4324_7(wires_1081_6[0], addr_1081_6, addr_positional[17299:17296], addr_4324_7);

wire[31:0] addr_4325_7;

Selector_2 s4325_7(wires_1081_6[1], addr_1081_6, addr_positional[17303:17300], addr_4325_7);

wire[31:0] addr_4326_7;

Selector_2 s4326_7(wires_1081_6[2], addr_1081_6, addr_positional[17307:17304], addr_4326_7);

wire[31:0] addr_4327_7;

Selector_2 s4327_7(wires_1081_6[3], addr_1081_6, addr_positional[17311:17308], addr_4327_7);

wire[31:0] addr_4328_7;

Selector_2 s4328_7(wires_1082_6[0], addr_1082_6, addr_positional[17315:17312], addr_4328_7);

wire[31:0] addr_4329_7;

Selector_2 s4329_7(wires_1082_6[1], addr_1082_6, addr_positional[17319:17316], addr_4329_7);

wire[31:0] addr_4330_7;

Selector_2 s4330_7(wires_1082_6[2], addr_1082_6, addr_positional[17323:17320], addr_4330_7);

wire[31:0] addr_4331_7;

Selector_2 s4331_7(wires_1082_6[3], addr_1082_6, addr_positional[17327:17324], addr_4331_7);

wire[31:0] addr_4332_7;

Selector_2 s4332_7(wires_1083_6[0], addr_1083_6, addr_positional[17331:17328], addr_4332_7);

wire[31:0] addr_4333_7;

Selector_2 s4333_7(wires_1083_6[1], addr_1083_6, addr_positional[17335:17332], addr_4333_7);

wire[31:0] addr_4334_7;

Selector_2 s4334_7(wires_1083_6[2], addr_1083_6, addr_positional[17339:17336], addr_4334_7);

wire[31:0] addr_4335_7;

Selector_2 s4335_7(wires_1083_6[3], addr_1083_6, addr_positional[17343:17340], addr_4335_7);

wire[31:0] addr_4336_7;

Selector_2 s4336_7(wires_1084_6[0], addr_1084_6, addr_positional[17347:17344], addr_4336_7);

wire[31:0] addr_4337_7;

Selector_2 s4337_7(wires_1084_6[1], addr_1084_6, addr_positional[17351:17348], addr_4337_7);

wire[31:0] addr_4338_7;

Selector_2 s4338_7(wires_1084_6[2], addr_1084_6, addr_positional[17355:17352], addr_4338_7);

wire[31:0] addr_4339_7;

Selector_2 s4339_7(wires_1084_6[3], addr_1084_6, addr_positional[17359:17356], addr_4339_7);

wire[31:0] addr_4340_7;

Selector_2 s4340_7(wires_1085_6[0], addr_1085_6, addr_positional[17363:17360], addr_4340_7);

wire[31:0] addr_4341_7;

Selector_2 s4341_7(wires_1085_6[1], addr_1085_6, addr_positional[17367:17364], addr_4341_7);

wire[31:0] addr_4342_7;

Selector_2 s4342_7(wires_1085_6[2], addr_1085_6, addr_positional[17371:17368], addr_4342_7);

wire[31:0] addr_4343_7;

Selector_2 s4343_7(wires_1085_6[3], addr_1085_6, addr_positional[17375:17372], addr_4343_7);

wire[31:0] addr_4344_7;

Selector_2 s4344_7(wires_1086_6[0], addr_1086_6, addr_positional[17379:17376], addr_4344_7);

wire[31:0] addr_4345_7;

Selector_2 s4345_7(wires_1086_6[1], addr_1086_6, addr_positional[17383:17380], addr_4345_7);

wire[31:0] addr_4346_7;

Selector_2 s4346_7(wires_1086_6[2], addr_1086_6, addr_positional[17387:17384], addr_4346_7);

wire[31:0] addr_4347_7;

Selector_2 s4347_7(wires_1086_6[3], addr_1086_6, addr_positional[17391:17388], addr_4347_7);

wire[31:0] addr_4348_7;

Selector_2 s4348_7(wires_1087_6[0], addr_1087_6, addr_positional[17395:17392], addr_4348_7);

wire[31:0] addr_4349_7;

Selector_2 s4349_7(wires_1087_6[1], addr_1087_6, addr_positional[17399:17396], addr_4349_7);

wire[31:0] addr_4350_7;

Selector_2 s4350_7(wires_1087_6[2], addr_1087_6, addr_positional[17403:17400], addr_4350_7);

wire[31:0] addr_4351_7;

Selector_2 s4351_7(wires_1087_6[3], addr_1087_6, addr_positional[17407:17404], addr_4351_7);

wire[31:0] addr_4352_7;

Selector_2 s4352_7(wires_1088_6[0], addr_1088_6, addr_positional[17411:17408], addr_4352_7);

wire[31:0] addr_4353_7;

Selector_2 s4353_7(wires_1088_6[1], addr_1088_6, addr_positional[17415:17412], addr_4353_7);

wire[31:0] addr_4354_7;

Selector_2 s4354_7(wires_1088_6[2], addr_1088_6, addr_positional[17419:17416], addr_4354_7);

wire[31:0] addr_4355_7;

Selector_2 s4355_7(wires_1088_6[3], addr_1088_6, addr_positional[17423:17420], addr_4355_7);

wire[31:0] addr_4356_7;

Selector_2 s4356_7(wires_1089_6[0], addr_1089_6, addr_positional[17427:17424], addr_4356_7);

wire[31:0] addr_4357_7;

Selector_2 s4357_7(wires_1089_6[1], addr_1089_6, addr_positional[17431:17428], addr_4357_7);

wire[31:0] addr_4358_7;

Selector_2 s4358_7(wires_1089_6[2], addr_1089_6, addr_positional[17435:17432], addr_4358_7);

wire[31:0] addr_4359_7;

Selector_2 s4359_7(wires_1089_6[3], addr_1089_6, addr_positional[17439:17436], addr_4359_7);

wire[31:0] addr_4360_7;

Selector_2 s4360_7(wires_1090_6[0], addr_1090_6, addr_positional[17443:17440], addr_4360_7);

wire[31:0] addr_4361_7;

Selector_2 s4361_7(wires_1090_6[1], addr_1090_6, addr_positional[17447:17444], addr_4361_7);

wire[31:0] addr_4362_7;

Selector_2 s4362_7(wires_1090_6[2], addr_1090_6, addr_positional[17451:17448], addr_4362_7);

wire[31:0] addr_4363_7;

Selector_2 s4363_7(wires_1090_6[3], addr_1090_6, addr_positional[17455:17452], addr_4363_7);

wire[31:0] addr_4364_7;

Selector_2 s4364_7(wires_1091_6[0], addr_1091_6, addr_positional[17459:17456], addr_4364_7);

wire[31:0] addr_4365_7;

Selector_2 s4365_7(wires_1091_6[1], addr_1091_6, addr_positional[17463:17460], addr_4365_7);

wire[31:0] addr_4366_7;

Selector_2 s4366_7(wires_1091_6[2], addr_1091_6, addr_positional[17467:17464], addr_4366_7);

wire[31:0] addr_4367_7;

Selector_2 s4367_7(wires_1091_6[3], addr_1091_6, addr_positional[17471:17468], addr_4367_7);

wire[31:0] addr_4368_7;

Selector_2 s4368_7(wires_1092_6[0], addr_1092_6, addr_positional[17475:17472], addr_4368_7);

wire[31:0] addr_4369_7;

Selector_2 s4369_7(wires_1092_6[1], addr_1092_6, addr_positional[17479:17476], addr_4369_7);

wire[31:0] addr_4370_7;

Selector_2 s4370_7(wires_1092_6[2], addr_1092_6, addr_positional[17483:17480], addr_4370_7);

wire[31:0] addr_4371_7;

Selector_2 s4371_7(wires_1092_6[3], addr_1092_6, addr_positional[17487:17484], addr_4371_7);

wire[31:0] addr_4372_7;

Selector_2 s4372_7(wires_1093_6[0], addr_1093_6, addr_positional[17491:17488], addr_4372_7);

wire[31:0] addr_4373_7;

Selector_2 s4373_7(wires_1093_6[1], addr_1093_6, addr_positional[17495:17492], addr_4373_7);

wire[31:0] addr_4374_7;

Selector_2 s4374_7(wires_1093_6[2], addr_1093_6, addr_positional[17499:17496], addr_4374_7);

wire[31:0] addr_4375_7;

Selector_2 s4375_7(wires_1093_6[3], addr_1093_6, addr_positional[17503:17500], addr_4375_7);

wire[31:0] addr_4376_7;

Selector_2 s4376_7(wires_1094_6[0], addr_1094_6, addr_positional[17507:17504], addr_4376_7);

wire[31:0] addr_4377_7;

Selector_2 s4377_7(wires_1094_6[1], addr_1094_6, addr_positional[17511:17508], addr_4377_7);

wire[31:0] addr_4378_7;

Selector_2 s4378_7(wires_1094_6[2], addr_1094_6, addr_positional[17515:17512], addr_4378_7);

wire[31:0] addr_4379_7;

Selector_2 s4379_7(wires_1094_6[3], addr_1094_6, addr_positional[17519:17516], addr_4379_7);

wire[31:0] addr_4380_7;

Selector_2 s4380_7(wires_1095_6[0], addr_1095_6, addr_positional[17523:17520], addr_4380_7);

wire[31:0] addr_4381_7;

Selector_2 s4381_7(wires_1095_6[1], addr_1095_6, addr_positional[17527:17524], addr_4381_7);

wire[31:0] addr_4382_7;

Selector_2 s4382_7(wires_1095_6[2], addr_1095_6, addr_positional[17531:17528], addr_4382_7);

wire[31:0] addr_4383_7;

Selector_2 s4383_7(wires_1095_6[3], addr_1095_6, addr_positional[17535:17532], addr_4383_7);

wire[31:0] addr_4384_7;

Selector_2 s4384_7(wires_1096_6[0], addr_1096_6, addr_positional[17539:17536], addr_4384_7);

wire[31:0] addr_4385_7;

Selector_2 s4385_7(wires_1096_6[1], addr_1096_6, addr_positional[17543:17540], addr_4385_7);

wire[31:0] addr_4386_7;

Selector_2 s4386_7(wires_1096_6[2], addr_1096_6, addr_positional[17547:17544], addr_4386_7);

wire[31:0] addr_4387_7;

Selector_2 s4387_7(wires_1096_6[3], addr_1096_6, addr_positional[17551:17548], addr_4387_7);

wire[31:0] addr_4388_7;

Selector_2 s4388_7(wires_1097_6[0], addr_1097_6, addr_positional[17555:17552], addr_4388_7);

wire[31:0] addr_4389_7;

Selector_2 s4389_7(wires_1097_6[1], addr_1097_6, addr_positional[17559:17556], addr_4389_7);

wire[31:0] addr_4390_7;

Selector_2 s4390_7(wires_1097_6[2], addr_1097_6, addr_positional[17563:17560], addr_4390_7);

wire[31:0] addr_4391_7;

Selector_2 s4391_7(wires_1097_6[3], addr_1097_6, addr_positional[17567:17564], addr_4391_7);

wire[31:0] addr_4392_7;

Selector_2 s4392_7(wires_1098_6[0], addr_1098_6, addr_positional[17571:17568], addr_4392_7);

wire[31:0] addr_4393_7;

Selector_2 s4393_7(wires_1098_6[1], addr_1098_6, addr_positional[17575:17572], addr_4393_7);

wire[31:0] addr_4394_7;

Selector_2 s4394_7(wires_1098_6[2], addr_1098_6, addr_positional[17579:17576], addr_4394_7);

wire[31:0] addr_4395_7;

Selector_2 s4395_7(wires_1098_6[3], addr_1098_6, addr_positional[17583:17580], addr_4395_7);

wire[31:0] addr_4396_7;

Selector_2 s4396_7(wires_1099_6[0], addr_1099_6, addr_positional[17587:17584], addr_4396_7);

wire[31:0] addr_4397_7;

Selector_2 s4397_7(wires_1099_6[1], addr_1099_6, addr_positional[17591:17588], addr_4397_7);

wire[31:0] addr_4398_7;

Selector_2 s4398_7(wires_1099_6[2], addr_1099_6, addr_positional[17595:17592], addr_4398_7);

wire[31:0] addr_4399_7;

Selector_2 s4399_7(wires_1099_6[3], addr_1099_6, addr_positional[17599:17596], addr_4399_7);

wire[31:0] addr_4400_7;

Selector_2 s4400_7(wires_1100_6[0], addr_1100_6, addr_positional[17603:17600], addr_4400_7);

wire[31:0] addr_4401_7;

Selector_2 s4401_7(wires_1100_6[1], addr_1100_6, addr_positional[17607:17604], addr_4401_7);

wire[31:0] addr_4402_7;

Selector_2 s4402_7(wires_1100_6[2], addr_1100_6, addr_positional[17611:17608], addr_4402_7);

wire[31:0] addr_4403_7;

Selector_2 s4403_7(wires_1100_6[3], addr_1100_6, addr_positional[17615:17612], addr_4403_7);

wire[31:0] addr_4404_7;

Selector_2 s4404_7(wires_1101_6[0], addr_1101_6, addr_positional[17619:17616], addr_4404_7);

wire[31:0] addr_4405_7;

Selector_2 s4405_7(wires_1101_6[1], addr_1101_6, addr_positional[17623:17620], addr_4405_7);

wire[31:0] addr_4406_7;

Selector_2 s4406_7(wires_1101_6[2], addr_1101_6, addr_positional[17627:17624], addr_4406_7);

wire[31:0] addr_4407_7;

Selector_2 s4407_7(wires_1101_6[3], addr_1101_6, addr_positional[17631:17628], addr_4407_7);

wire[31:0] addr_4408_7;

Selector_2 s4408_7(wires_1102_6[0], addr_1102_6, addr_positional[17635:17632], addr_4408_7);

wire[31:0] addr_4409_7;

Selector_2 s4409_7(wires_1102_6[1], addr_1102_6, addr_positional[17639:17636], addr_4409_7);

wire[31:0] addr_4410_7;

Selector_2 s4410_7(wires_1102_6[2], addr_1102_6, addr_positional[17643:17640], addr_4410_7);

wire[31:0] addr_4411_7;

Selector_2 s4411_7(wires_1102_6[3], addr_1102_6, addr_positional[17647:17644], addr_4411_7);

wire[31:0] addr_4412_7;

Selector_2 s4412_7(wires_1103_6[0], addr_1103_6, addr_positional[17651:17648], addr_4412_7);

wire[31:0] addr_4413_7;

Selector_2 s4413_7(wires_1103_6[1], addr_1103_6, addr_positional[17655:17652], addr_4413_7);

wire[31:0] addr_4414_7;

Selector_2 s4414_7(wires_1103_6[2], addr_1103_6, addr_positional[17659:17656], addr_4414_7);

wire[31:0] addr_4415_7;

Selector_2 s4415_7(wires_1103_6[3], addr_1103_6, addr_positional[17663:17660], addr_4415_7);

wire[31:0] addr_4416_7;

Selector_2 s4416_7(wires_1104_6[0], addr_1104_6, addr_positional[17667:17664], addr_4416_7);

wire[31:0] addr_4417_7;

Selector_2 s4417_7(wires_1104_6[1], addr_1104_6, addr_positional[17671:17668], addr_4417_7);

wire[31:0] addr_4418_7;

Selector_2 s4418_7(wires_1104_6[2], addr_1104_6, addr_positional[17675:17672], addr_4418_7);

wire[31:0] addr_4419_7;

Selector_2 s4419_7(wires_1104_6[3], addr_1104_6, addr_positional[17679:17676], addr_4419_7);

wire[31:0] addr_4420_7;

Selector_2 s4420_7(wires_1105_6[0], addr_1105_6, addr_positional[17683:17680], addr_4420_7);

wire[31:0] addr_4421_7;

Selector_2 s4421_7(wires_1105_6[1], addr_1105_6, addr_positional[17687:17684], addr_4421_7);

wire[31:0] addr_4422_7;

Selector_2 s4422_7(wires_1105_6[2], addr_1105_6, addr_positional[17691:17688], addr_4422_7);

wire[31:0] addr_4423_7;

Selector_2 s4423_7(wires_1105_6[3], addr_1105_6, addr_positional[17695:17692], addr_4423_7);

wire[31:0] addr_4424_7;

Selector_2 s4424_7(wires_1106_6[0], addr_1106_6, addr_positional[17699:17696], addr_4424_7);

wire[31:0] addr_4425_7;

Selector_2 s4425_7(wires_1106_6[1], addr_1106_6, addr_positional[17703:17700], addr_4425_7);

wire[31:0] addr_4426_7;

Selector_2 s4426_7(wires_1106_6[2], addr_1106_6, addr_positional[17707:17704], addr_4426_7);

wire[31:0] addr_4427_7;

Selector_2 s4427_7(wires_1106_6[3], addr_1106_6, addr_positional[17711:17708], addr_4427_7);

wire[31:0] addr_4428_7;

Selector_2 s4428_7(wires_1107_6[0], addr_1107_6, addr_positional[17715:17712], addr_4428_7);

wire[31:0] addr_4429_7;

Selector_2 s4429_7(wires_1107_6[1], addr_1107_6, addr_positional[17719:17716], addr_4429_7);

wire[31:0] addr_4430_7;

Selector_2 s4430_7(wires_1107_6[2], addr_1107_6, addr_positional[17723:17720], addr_4430_7);

wire[31:0] addr_4431_7;

Selector_2 s4431_7(wires_1107_6[3], addr_1107_6, addr_positional[17727:17724], addr_4431_7);

wire[31:0] addr_4432_7;

Selector_2 s4432_7(wires_1108_6[0], addr_1108_6, addr_positional[17731:17728], addr_4432_7);

wire[31:0] addr_4433_7;

Selector_2 s4433_7(wires_1108_6[1], addr_1108_6, addr_positional[17735:17732], addr_4433_7);

wire[31:0] addr_4434_7;

Selector_2 s4434_7(wires_1108_6[2], addr_1108_6, addr_positional[17739:17736], addr_4434_7);

wire[31:0] addr_4435_7;

Selector_2 s4435_7(wires_1108_6[3], addr_1108_6, addr_positional[17743:17740], addr_4435_7);

wire[31:0] addr_4436_7;

Selector_2 s4436_7(wires_1109_6[0], addr_1109_6, addr_positional[17747:17744], addr_4436_7);

wire[31:0] addr_4437_7;

Selector_2 s4437_7(wires_1109_6[1], addr_1109_6, addr_positional[17751:17748], addr_4437_7);

wire[31:0] addr_4438_7;

Selector_2 s4438_7(wires_1109_6[2], addr_1109_6, addr_positional[17755:17752], addr_4438_7);

wire[31:0] addr_4439_7;

Selector_2 s4439_7(wires_1109_6[3], addr_1109_6, addr_positional[17759:17756], addr_4439_7);

wire[31:0] addr_4440_7;

Selector_2 s4440_7(wires_1110_6[0], addr_1110_6, addr_positional[17763:17760], addr_4440_7);

wire[31:0] addr_4441_7;

Selector_2 s4441_7(wires_1110_6[1], addr_1110_6, addr_positional[17767:17764], addr_4441_7);

wire[31:0] addr_4442_7;

Selector_2 s4442_7(wires_1110_6[2], addr_1110_6, addr_positional[17771:17768], addr_4442_7);

wire[31:0] addr_4443_7;

Selector_2 s4443_7(wires_1110_6[3], addr_1110_6, addr_positional[17775:17772], addr_4443_7);

wire[31:0] addr_4444_7;

Selector_2 s4444_7(wires_1111_6[0], addr_1111_6, addr_positional[17779:17776], addr_4444_7);

wire[31:0] addr_4445_7;

Selector_2 s4445_7(wires_1111_6[1], addr_1111_6, addr_positional[17783:17780], addr_4445_7);

wire[31:0] addr_4446_7;

Selector_2 s4446_7(wires_1111_6[2], addr_1111_6, addr_positional[17787:17784], addr_4446_7);

wire[31:0] addr_4447_7;

Selector_2 s4447_7(wires_1111_6[3], addr_1111_6, addr_positional[17791:17788], addr_4447_7);

wire[31:0] addr_4448_7;

Selector_2 s4448_7(wires_1112_6[0], addr_1112_6, addr_positional[17795:17792], addr_4448_7);

wire[31:0] addr_4449_7;

Selector_2 s4449_7(wires_1112_6[1], addr_1112_6, addr_positional[17799:17796], addr_4449_7);

wire[31:0] addr_4450_7;

Selector_2 s4450_7(wires_1112_6[2], addr_1112_6, addr_positional[17803:17800], addr_4450_7);

wire[31:0] addr_4451_7;

Selector_2 s4451_7(wires_1112_6[3], addr_1112_6, addr_positional[17807:17804], addr_4451_7);

wire[31:0] addr_4452_7;

Selector_2 s4452_7(wires_1113_6[0], addr_1113_6, addr_positional[17811:17808], addr_4452_7);

wire[31:0] addr_4453_7;

Selector_2 s4453_7(wires_1113_6[1], addr_1113_6, addr_positional[17815:17812], addr_4453_7);

wire[31:0] addr_4454_7;

Selector_2 s4454_7(wires_1113_6[2], addr_1113_6, addr_positional[17819:17816], addr_4454_7);

wire[31:0] addr_4455_7;

Selector_2 s4455_7(wires_1113_6[3], addr_1113_6, addr_positional[17823:17820], addr_4455_7);

wire[31:0] addr_4456_7;

Selector_2 s4456_7(wires_1114_6[0], addr_1114_6, addr_positional[17827:17824], addr_4456_7);

wire[31:0] addr_4457_7;

Selector_2 s4457_7(wires_1114_6[1], addr_1114_6, addr_positional[17831:17828], addr_4457_7);

wire[31:0] addr_4458_7;

Selector_2 s4458_7(wires_1114_6[2], addr_1114_6, addr_positional[17835:17832], addr_4458_7);

wire[31:0] addr_4459_7;

Selector_2 s4459_7(wires_1114_6[3], addr_1114_6, addr_positional[17839:17836], addr_4459_7);

wire[31:0] addr_4460_7;

Selector_2 s4460_7(wires_1115_6[0], addr_1115_6, addr_positional[17843:17840], addr_4460_7);

wire[31:0] addr_4461_7;

Selector_2 s4461_7(wires_1115_6[1], addr_1115_6, addr_positional[17847:17844], addr_4461_7);

wire[31:0] addr_4462_7;

Selector_2 s4462_7(wires_1115_6[2], addr_1115_6, addr_positional[17851:17848], addr_4462_7);

wire[31:0] addr_4463_7;

Selector_2 s4463_7(wires_1115_6[3], addr_1115_6, addr_positional[17855:17852], addr_4463_7);

wire[31:0] addr_4464_7;

Selector_2 s4464_7(wires_1116_6[0], addr_1116_6, addr_positional[17859:17856], addr_4464_7);

wire[31:0] addr_4465_7;

Selector_2 s4465_7(wires_1116_6[1], addr_1116_6, addr_positional[17863:17860], addr_4465_7);

wire[31:0] addr_4466_7;

Selector_2 s4466_7(wires_1116_6[2], addr_1116_6, addr_positional[17867:17864], addr_4466_7);

wire[31:0] addr_4467_7;

Selector_2 s4467_7(wires_1116_6[3], addr_1116_6, addr_positional[17871:17868], addr_4467_7);

wire[31:0] addr_4468_7;

Selector_2 s4468_7(wires_1117_6[0], addr_1117_6, addr_positional[17875:17872], addr_4468_7);

wire[31:0] addr_4469_7;

Selector_2 s4469_7(wires_1117_6[1], addr_1117_6, addr_positional[17879:17876], addr_4469_7);

wire[31:0] addr_4470_7;

Selector_2 s4470_7(wires_1117_6[2], addr_1117_6, addr_positional[17883:17880], addr_4470_7);

wire[31:0] addr_4471_7;

Selector_2 s4471_7(wires_1117_6[3], addr_1117_6, addr_positional[17887:17884], addr_4471_7);

wire[31:0] addr_4472_7;

Selector_2 s4472_7(wires_1118_6[0], addr_1118_6, addr_positional[17891:17888], addr_4472_7);

wire[31:0] addr_4473_7;

Selector_2 s4473_7(wires_1118_6[1], addr_1118_6, addr_positional[17895:17892], addr_4473_7);

wire[31:0] addr_4474_7;

Selector_2 s4474_7(wires_1118_6[2], addr_1118_6, addr_positional[17899:17896], addr_4474_7);

wire[31:0] addr_4475_7;

Selector_2 s4475_7(wires_1118_6[3], addr_1118_6, addr_positional[17903:17900], addr_4475_7);

wire[31:0] addr_4476_7;

Selector_2 s4476_7(wires_1119_6[0], addr_1119_6, addr_positional[17907:17904], addr_4476_7);

wire[31:0] addr_4477_7;

Selector_2 s4477_7(wires_1119_6[1], addr_1119_6, addr_positional[17911:17908], addr_4477_7);

wire[31:0] addr_4478_7;

Selector_2 s4478_7(wires_1119_6[2], addr_1119_6, addr_positional[17915:17912], addr_4478_7);

wire[31:0] addr_4479_7;

Selector_2 s4479_7(wires_1119_6[3], addr_1119_6, addr_positional[17919:17916], addr_4479_7);

wire[31:0] addr_4480_7;

Selector_2 s4480_7(wires_1120_6[0], addr_1120_6, addr_positional[17923:17920], addr_4480_7);

wire[31:0] addr_4481_7;

Selector_2 s4481_7(wires_1120_6[1], addr_1120_6, addr_positional[17927:17924], addr_4481_7);

wire[31:0] addr_4482_7;

Selector_2 s4482_7(wires_1120_6[2], addr_1120_6, addr_positional[17931:17928], addr_4482_7);

wire[31:0] addr_4483_7;

Selector_2 s4483_7(wires_1120_6[3], addr_1120_6, addr_positional[17935:17932], addr_4483_7);

wire[31:0] addr_4484_7;

Selector_2 s4484_7(wires_1121_6[0], addr_1121_6, addr_positional[17939:17936], addr_4484_7);

wire[31:0] addr_4485_7;

Selector_2 s4485_7(wires_1121_6[1], addr_1121_6, addr_positional[17943:17940], addr_4485_7);

wire[31:0] addr_4486_7;

Selector_2 s4486_7(wires_1121_6[2], addr_1121_6, addr_positional[17947:17944], addr_4486_7);

wire[31:0] addr_4487_7;

Selector_2 s4487_7(wires_1121_6[3], addr_1121_6, addr_positional[17951:17948], addr_4487_7);

wire[31:0] addr_4488_7;

Selector_2 s4488_7(wires_1122_6[0], addr_1122_6, addr_positional[17955:17952], addr_4488_7);

wire[31:0] addr_4489_7;

Selector_2 s4489_7(wires_1122_6[1], addr_1122_6, addr_positional[17959:17956], addr_4489_7);

wire[31:0] addr_4490_7;

Selector_2 s4490_7(wires_1122_6[2], addr_1122_6, addr_positional[17963:17960], addr_4490_7);

wire[31:0] addr_4491_7;

Selector_2 s4491_7(wires_1122_6[3], addr_1122_6, addr_positional[17967:17964], addr_4491_7);

wire[31:0] addr_4492_7;

Selector_2 s4492_7(wires_1123_6[0], addr_1123_6, addr_positional[17971:17968], addr_4492_7);

wire[31:0] addr_4493_7;

Selector_2 s4493_7(wires_1123_6[1], addr_1123_6, addr_positional[17975:17972], addr_4493_7);

wire[31:0] addr_4494_7;

Selector_2 s4494_7(wires_1123_6[2], addr_1123_6, addr_positional[17979:17976], addr_4494_7);

wire[31:0] addr_4495_7;

Selector_2 s4495_7(wires_1123_6[3], addr_1123_6, addr_positional[17983:17980], addr_4495_7);

wire[31:0] addr_4496_7;

Selector_2 s4496_7(wires_1124_6[0], addr_1124_6, addr_positional[17987:17984], addr_4496_7);

wire[31:0] addr_4497_7;

Selector_2 s4497_7(wires_1124_6[1], addr_1124_6, addr_positional[17991:17988], addr_4497_7);

wire[31:0] addr_4498_7;

Selector_2 s4498_7(wires_1124_6[2], addr_1124_6, addr_positional[17995:17992], addr_4498_7);

wire[31:0] addr_4499_7;

Selector_2 s4499_7(wires_1124_6[3], addr_1124_6, addr_positional[17999:17996], addr_4499_7);

wire[31:0] addr_4500_7;

Selector_2 s4500_7(wires_1125_6[0], addr_1125_6, addr_positional[18003:18000], addr_4500_7);

wire[31:0] addr_4501_7;

Selector_2 s4501_7(wires_1125_6[1], addr_1125_6, addr_positional[18007:18004], addr_4501_7);

wire[31:0] addr_4502_7;

Selector_2 s4502_7(wires_1125_6[2], addr_1125_6, addr_positional[18011:18008], addr_4502_7);

wire[31:0] addr_4503_7;

Selector_2 s4503_7(wires_1125_6[3], addr_1125_6, addr_positional[18015:18012], addr_4503_7);

wire[31:0] addr_4504_7;

Selector_2 s4504_7(wires_1126_6[0], addr_1126_6, addr_positional[18019:18016], addr_4504_7);

wire[31:0] addr_4505_7;

Selector_2 s4505_7(wires_1126_6[1], addr_1126_6, addr_positional[18023:18020], addr_4505_7);

wire[31:0] addr_4506_7;

Selector_2 s4506_7(wires_1126_6[2], addr_1126_6, addr_positional[18027:18024], addr_4506_7);

wire[31:0] addr_4507_7;

Selector_2 s4507_7(wires_1126_6[3], addr_1126_6, addr_positional[18031:18028], addr_4507_7);

wire[31:0] addr_4508_7;

Selector_2 s4508_7(wires_1127_6[0], addr_1127_6, addr_positional[18035:18032], addr_4508_7);

wire[31:0] addr_4509_7;

Selector_2 s4509_7(wires_1127_6[1], addr_1127_6, addr_positional[18039:18036], addr_4509_7);

wire[31:0] addr_4510_7;

Selector_2 s4510_7(wires_1127_6[2], addr_1127_6, addr_positional[18043:18040], addr_4510_7);

wire[31:0] addr_4511_7;

Selector_2 s4511_7(wires_1127_6[3], addr_1127_6, addr_positional[18047:18044], addr_4511_7);

wire[31:0] addr_4512_7;

Selector_2 s4512_7(wires_1128_6[0], addr_1128_6, addr_positional[18051:18048], addr_4512_7);

wire[31:0] addr_4513_7;

Selector_2 s4513_7(wires_1128_6[1], addr_1128_6, addr_positional[18055:18052], addr_4513_7);

wire[31:0] addr_4514_7;

Selector_2 s4514_7(wires_1128_6[2], addr_1128_6, addr_positional[18059:18056], addr_4514_7);

wire[31:0] addr_4515_7;

Selector_2 s4515_7(wires_1128_6[3], addr_1128_6, addr_positional[18063:18060], addr_4515_7);

wire[31:0] addr_4516_7;

Selector_2 s4516_7(wires_1129_6[0], addr_1129_6, addr_positional[18067:18064], addr_4516_7);

wire[31:0] addr_4517_7;

Selector_2 s4517_7(wires_1129_6[1], addr_1129_6, addr_positional[18071:18068], addr_4517_7);

wire[31:0] addr_4518_7;

Selector_2 s4518_7(wires_1129_6[2], addr_1129_6, addr_positional[18075:18072], addr_4518_7);

wire[31:0] addr_4519_7;

Selector_2 s4519_7(wires_1129_6[3], addr_1129_6, addr_positional[18079:18076], addr_4519_7);

wire[31:0] addr_4520_7;

Selector_2 s4520_7(wires_1130_6[0], addr_1130_6, addr_positional[18083:18080], addr_4520_7);

wire[31:0] addr_4521_7;

Selector_2 s4521_7(wires_1130_6[1], addr_1130_6, addr_positional[18087:18084], addr_4521_7);

wire[31:0] addr_4522_7;

Selector_2 s4522_7(wires_1130_6[2], addr_1130_6, addr_positional[18091:18088], addr_4522_7);

wire[31:0] addr_4523_7;

Selector_2 s4523_7(wires_1130_6[3], addr_1130_6, addr_positional[18095:18092], addr_4523_7);

wire[31:0] addr_4524_7;

Selector_2 s4524_7(wires_1131_6[0], addr_1131_6, addr_positional[18099:18096], addr_4524_7);

wire[31:0] addr_4525_7;

Selector_2 s4525_7(wires_1131_6[1], addr_1131_6, addr_positional[18103:18100], addr_4525_7);

wire[31:0] addr_4526_7;

Selector_2 s4526_7(wires_1131_6[2], addr_1131_6, addr_positional[18107:18104], addr_4526_7);

wire[31:0] addr_4527_7;

Selector_2 s4527_7(wires_1131_6[3], addr_1131_6, addr_positional[18111:18108], addr_4527_7);

wire[31:0] addr_4528_7;

Selector_2 s4528_7(wires_1132_6[0], addr_1132_6, addr_positional[18115:18112], addr_4528_7);

wire[31:0] addr_4529_7;

Selector_2 s4529_7(wires_1132_6[1], addr_1132_6, addr_positional[18119:18116], addr_4529_7);

wire[31:0] addr_4530_7;

Selector_2 s4530_7(wires_1132_6[2], addr_1132_6, addr_positional[18123:18120], addr_4530_7);

wire[31:0] addr_4531_7;

Selector_2 s4531_7(wires_1132_6[3], addr_1132_6, addr_positional[18127:18124], addr_4531_7);

wire[31:0] addr_4532_7;

Selector_2 s4532_7(wires_1133_6[0], addr_1133_6, addr_positional[18131:18128], addr_4532_7);

wire[31:0] addr_4533_7;

Selector_2 s4533_7(wires_1133_6[1], addr_1133_6, addr_positional[18135:18132], addr_4533_7);

wire[31:0] addr_4534_7;

Selector_2 s4534_7(wires_1133_6[2], addr_1133_6, addr_positional[18139:18136], addr_4534_7);

wire[31:0] addr_4535_7;

Selector_2 s4535_7(wires_1133_6[3], addr_1133_6, addr_positional[18143:18140], addr_4535_7);

wire[31:0] addr_4536_7;

Selector_2 s4536_7(wires_1134_6[0], addr_1134_6, addr_positional[18147:18144], addr_4536_7);

wire[31:0] addr_4537_7;

Selector_2 s4537_7(wires_1134_6[1], addr_1134_6, addr_positional[18151:18148], addr_4537_7);

wire[31:0] addr_4538_7;

Selector_2 s4538_7(wires_1134_6[2], addr_1134_6, addr_positional[18155:18152], addr_4538_7);

wire[31:0] addr_4539_7;

Selector_2 s4539_7(wires_1134_6[3], addr_1134_6, addr_positional[18159:18156], addr_4539_7);

wire[31:0] addr_4540_7;

Selector_2 s4540_7(wires_1135_6[0], addr_1135_6, addr_positional[18163:18160], addr_4540_7);

wire[31:0] addr_4541_7;

Selector_2 s4541_7(wires_1135_6[1], addr_1135_6, addr_positional[18167:18164], addr_4541_7);

wire[31:0] addr_4542_7;

Selector_2 s4542_7(wires_1135_6[2], addr_1135_6, addr_positional[18171:18168], addr_4542_7);

wire[31:0] addr_4543_7;

Selector_2 s4543_7(wires_1135_6[3], addr_1135_6, addr_positional[18175:18172], addr_4543_7);

wire[31:0] addr_4544_7;

Selector_2 s4544_7(wires_1136_6[0], addr_1136_6, addr_positional[18179:18176], addr_4544_7);

wire[31:0] addr_4545_7;

Selector_2 s4545_7(wires_1136_6[1], addr_1136_6, addr_positional[18183:18180], addr_4545_7);

wire[31:0] addr_4546_7;

Selector_2 s4546_7(wires_1136_6[2], addr_1136_6, addr_positional[18187:18184], addr_4546_7);

wire[31:0] addr_4547_7;

Selector_2 s4547_7(wires_1136_6[3], addr_1136_6, addr_positional[18191:18188], addr_4547_7);

wire[31:0] addr_4548_7;

Selector_2 s4548_7(wires_1137_6[0], addr_1137_6, addr_positional[18195:18192], addr_4548_7);

wire[31:0] addr_4549_7;

Selector_2 s4549_7(wires_1137_6[1], addr_1137_6, addr_positional[18199:18196], addr_4549_7);

wire[31:0] addr_4550_7;

Selector_2 s4550_7(wires_1137_6[2], addr_1137_6, addr_positional[18203:18200], addr_4550_7);

wire[31:0] addr_4551_7;

Selector_2 s4551_7(wires_1137_6[3], addr_1137_6, addr_positional[18207:18204], addr_4551_7);

wire[31:0] addr_4552_7;

Selector_2 s4552_7(wires_1138_6[0], addr_1138_6, addr_positional[18211:18208], addr_4552_7);

wire[31:0] addr_4553_7;

Selector_2 s4553_7(wires_1138_6[1], addr_1138_6, addr_positional[18215:18212], addr_4553_7);

wire[31:0] addr_4554_7;

Selector_2 s4554_7(wires_1138_6[2], addr_1138_6, addr_positional[18219:18216], addr_4554_7);

wire[31:0] addr_4555_7;

Selector_2 s4555_7(wires_1138_6[3], addr_1138_6, addr_positional[18223:18220], addr_4555_7);

wire[31:0] addr_4556_7;

Selector_2 s4556_7(wires_1139_6[0], addr_1139_6, addr_positional[18227:18224], addr_4556_7);

wire[31:0] addr_4557_7;

Selector_2 s4557_7(wires_1139_6[1], addr_1139_6, addr_positional[18231:18228], addr_4557_7);

wire[31:0] addr_4558_7;

Selector_2 s4558_7(wires_1139_6[2], addr_1139_6, addr_positional[18235:18232], addr_4558_7);

wire[31:0] addr_4559_7;

Selector_2 s4559_7(wires_1139_6[3], addr_1139_6, addr_positional[18239:18236], addr_4559_7);

wire[31:0] addr_4560_7;

Selector_2 s4560_7(wires_1140_6[0], addr_1140_6, addr_positional[18243:18240], addr_4560_7);

wire[31:0] addr_4561_7;

Selector_2 s4561_7(wires_1140_6[1], addr_1140_6, addr_positional[18247:18244], addr_4561_7);

wire[31:0] addr_4562_7;

Selector_2 s4562_7(wires_1140_6[2], addr_1140_6, addr_positional[18251:18248], addr_4562_7);

wire[31:0] addr_4563_7;

Selector_2 s4563_7(wires_1140_6[3], addr_1140_6, addr_positional[18255:18252], addr_4563_7);

wire[31:0] addr_4564_7;

Selector_2 s4564_7(wires_1141_6[0], addr_1141_6, addr_positional[18259:18256], addr_4564_7);

wire[31:0] addr_4565_7;

Selector_2 s4565_7(wires_1141_6[1], addr_1141_6, addr_positional[18263:18260], addr_4565_7);

wire[31:0] addr_4566_7;

Selector_2 s4566_7(wires_1141_6[2], addr_1141_6, addr_positional[18267:18264], addr_4566_7);

wire[31:0] addr_4567_7;

Selector_2 s4567_7(wires_1141_6[3], addr_1141_6, addr_positional[18271:18268], addr_4567_7);

wire[31:0] addr_4568_7;

Selector_2 s4568_7(wires_1142_6[0], addr_1142_6, addr_positional[18275:18272], addr_4568_7);

wire[31:0] addr_4569_7;

Selector_2 s4569_7(wires_1142_6[1], addr_1142_6, addr_positional[18279:18276], addr_4569_7);

wire[31:0] addr_4570_7;

Selector_2 s4570_7(wires_1142_6[2], addr_1142_6, addr_positional[18283:18280], addr_4570_7);

wire[31:0] addr_4571_7;

Selector_2 s4571_7(wires_1142_6[3], addr_1142_6, addr_positional[18287:18284], addr_4571_7);

wire[31:0] addr_4572_7;

Selector_2 s4572_7(wires_1143_6[0], addr_1143_6, addr_positional[18291:18288], addr_4572_7);

wire[31:0] addr_4573_7;

Selector_2 s4573_7(wires_1143_6[1], addr_1143_6, addr_positional[18295:18292], addr_4573_7);

wire[31:0] addr_4574_7;

Selector_2 s4574_7(wires_1143_6[2], addr_1143_6, addr_positional[18299:18296], addr_4574_7);

wire[31:0] addr_4575_7;

Selector_2 s4575_7(wires_1143_6[3], addr_1143_6, addr_positional[18303:18300], addr_4575_7);

wire[31:0] addr_4576_7;

Selector_2 s4576_7(wires_1144_6[0], addr_1144_6, addr_positional[18307:18304], addr_4576_7);

wire[31:0] addr_4577_7;

Selector_2 s4577_7(wires_1144_6[1], addr_1144_6, addr_positional[18311:18308], addr_4577_7);

wire[31:0] addr_4578_7;

Selector_2 s4578_7(wires_1144_6[2], addr_1144_6, addr_positional[18315:18312], addr_4578_7);

wire[31:0] addr_4579_7;

Selector_2 s4579_7(wires_1144_6[3], addr_1144_6, addr_positional[18319:18316], addr_4579_7);

wire[31:0] addr_4580_7;

Selector_2 s4580_7(wires_1145_6[0], addr_1145_6, addr_positional[18323:18320], addr_4580_7);

wire[31:0] addr_4581_7;

Selector_2 s4581_7(wires_1145_6[1], addr_1145_6, addr_positional[18327:18324], addr_4581_7);

wire[31:0] addr_4582_7;

Selector_2 s4582_7(wires_1145_6[2], addr_1145_6, addr_positional[18331:18328], addr_4582_7);

wire[31:0] addr_4583_7;

Selector_2 s4583_7(wires_1145_6[3], addr_1145_6, addr_positional[18335:18332], addr_4583_7);

wire[31:0] addr_4584_7;

Selector_2 s4584_7(wires_1146_6[0], addr_1146_6, addr_positional[18339:18336], addr_4584_7);

wire[31:0] addr_4585_7;

Selector_2 s4585_7(wires_1146_6[1], addr_1146_6, addr_positional[18343:18340], addr_4585_7);

wire[31:0] addr_4586_7;

Selector_2 s4586_7(wires_1146_6[2], addr_1146_6, addr_positional[18347:18344], addr_4586_7);

wire[31:0] addr_4587_7;

Selector_2 s4587_7(wires_1146_6[3], addr_1146_6, addr_positional[18351:18348], addr_4587_7);

wire[31:0] addr_4588_7;

Selector_2 s4588_7(wires_1147_6[0], addr_1147_6, addr_positional[18355:18352], addr_4588_7);

wire[31:0] addr_4589_7;

Selector_2 s4589_7(wires_1147_6[1], addr_1147_6, addr_positional[18359:18356], addr_4589_7);

wire[31:0] addr_4590_7;

Selector_2 s4590_7(wires_1147_6[2], addr_1147_6, addr_positional[18363:18360], addr_4590_7);

wire[31:0] addr_4591_7;

Selector_2 s4591_7(wires_1147_6[3], addr_1147_6, addr_positional[18367:18364], addr_4591_7);

wire[31:0] addr_4592_7;

Selector_2 s4592_7(wires_1148_6[0], addr_1148_6, addr_positional[18371:18368], addr_4592_7);

wire[31:0] addr_4593_7;

Selector_2 s4593_7(wires_1148_6[1], addr_1148_6, addr_positional[18375:18372], addr_4593_7);

wire[31:0] addr_4594_7;

Selector_2 s4594_7(wires_1148_6[2], addr_1148_6, addr_positional[18379:18376], addr_4594_7);

wire[31:0] addr_4595_7;

Selector_2 s4595_7(wires_1148_6[3], addr_1148_6, addr_positional[18383:18380], addr_4595_7);

wire[31:0] addr_4596_7;

Selector_2 s4596_7(wires_1149_6[0], addr_1149_6, addr_positional[18387:18384], addr_4596_7);

wire[31:0] addr_4597_7;

Selector_2 s4597_7(wires_1149_6[1], addr_1149_6, addr_positional[18391:18388], addr_4597_7);

wire[31:0] addr_4598_7;

Selector_2 s4598_7(wires_1149_6[2], addr_1149_6, addr_positional[18395:18392], addr_4598_7);

wire[31:0] addr_4599_7;

Selector_2 s4599_7(wires_1149_6[3], addr_1149_6, addr_positional[18399:18396], addr_4599_7);

wire[31:0] addr_4600_7;

Selector_2 s4600_7(wires_1150_6[0], addr_1150_6, addr_positional[18403:18400], addr_4600_7);

wire[31:0] addr_4601_7;

Selector_2 s4601_7(wires_1150_6[1], addr_1150_6, addr_positional[18407:18404], addr_4601_7);

wire[31:0] addr_4602_7;

Selector_2 s4602_7(wires_1150_6[2], addr_1150_6, addr_positional[18411:18408], addr_4602_7);

wire[31:0] addr_4603_7;

Selector_2 s4603_7(wires_1150_6[3], addr_1150_6, addr_positional[18415:18412], addr_4603_7);

wire[31:0] addr_4604_7;

Selector_2 s4604_7(wires_1151_6[0], addr_1151_6, addr_positional[18419:18416], addr_4604_7);

wire[31:0] addr_4605_7;

Selector_2 s4605_7(wires_1151_6[1], addr_1151_6, addr_positional[18423:18420], addr_4605_7);

wire[31:0] addr_4606_7;

Selector_2 s4606_7(wires_1151_6[2], addr_1151_6, addr_positional[18427:18424], addr_4606_7);

wire[31:0] addr_4607_7;

Selector_2 s4607_7(wires_1151_6[3], addr_1151_6, addr_positional[18431:18428], addr_4607_7);

wire[31:0] addr_4608_7;

Selector_2 s4608_7(wires_1152_6[0], addr_1152_6, addr_positional[18435:18432], addr_4608_7);

wire[31:0] addr_4609_7;

Selector_2 s4609_7(wires_1152_6[1], addr_1152_6, addr_positional[18439:18436], addr_4609_7);

wire[31:0] addr_4610_7;

Selector_2 s4610_7(wires_1152_6[2], addr_1152_6, addr_positional[18443:18440], addr_4610_7);

wire[31:0] addr_4611_7;

Selector_2 s4611_7(wires_1152_6[3], addr_1152_6, addr_positional[18447:18444], addr_4611_7);

wire[31:0] addr_4612_7;

Selector_2 s4612_7(wires_1153_6[0], addr_1153_6, addr_positional[18451:18448], addr_4612_7);

wire[31:0] addr_4613_7;

Selector_2 s4613_7(wires_1153_6[1], addr_1153_6, addr_positional[18455:18452], addr_4613_7);

wire[31:0] addr_4614_7;

Selector_2 s4614_7(wires_1153_6[2], addr_1153_6, addr_positional[18459:18456], addr_4614_7);

wire[31:0] addr_4615_7;

Selector_2 s4615_7(wires_1153_6[3], addr_1153_6, addr_positional[18463:18460], addr_4615_7);

wire[31:0] addr_4616_7;

Selector_2 s4616_7(wires_1154_6[0], addr_1154_6, addr_positional[18467:18464], addr_4616_7);

wire[31:0] addr_4617_7;

Selector_2 s4617_7(wires_1154_6[1], addr_1154_6, addr_positional[18471:18468], addr_4617_7);

wire[31:0] addr_4618_7;

Selector_2 s4618_7(wires_1154_6[2], addr_1154_6, addr_positional[18475:18472], addr_4618_7);

wire[31:0] addr_4619_7;

Selector_2 s4619_7(wires_1154_6[3], addr_1154_6, addr_positional[18479:18476], addr_4619_7);

wire[31:0] addr_4620_7;

Selector_2 s4620_7(wires_1155_6[0], addr_1155_6, addr_positional[18483:18480], addr_4620_7);

wire[31:0] addr_4621_7;

Selector_2 s4621_7(wires_1155_6[1], addr_1155_6, addr_positional[18487:18484], addr_4621_7);

wire[31:0] addr_4622_7;

Selector_2 s4622_7(wires_1155_6[2], addr_1155_6, addr_positional[18491:18488], addr_4622_7);

wire[31:0] addr_4623_7;

Selector_2 s4623_7(wires_1155_6[3], addr_1155_6, addr_positional[18495:18492], addr_4623_7);

wire[31:0] addr_4624_7;

Selector_2 s4624_7(wires_1156_6[0], addr_1156_6, addr_positional[18499:18496], addr_4624_7);

wire[31:0] addr_4625_7;

Selector_2 s4625_7(wires_1156_6[1], addr_1156_6, addr_positional[18503:18500], addr_4625_7);

wire[31:0] addr_4626_7;

Selector_2 s4626_7(wires_1156_6[2], addr_1156_6, addr_positional[18507:18504], addr_4626_7);

wire[31:0] addr_4627_7;

Selector_2 s4627_7(wires_1156_6[3], addr_1156_6, addr_positional[18511:18508], addr_4627_7);

wire[31:0] addr_4628_7;

Selector_2 s4628_7(wires_1157_6[0], addr_1157_6, addr_positional[18515:18512], addr_4628_7);

wire[31:0] addr_4629_7;

Selector_2 s4629_7(wires_1157_6[1], addr_1157_6, addr_positional[18519:18516], addr_4629_7);

wire[31:0] addr_4630_7;

Selector_2 s4630_7(wires_1157_6[2], addr_1157_6, addr_positional[18523:18520], addr_4630_7);

wire[31:0] addr_4631_7;

Selector_2 s4631_7(wires_1157_6[3], addr_1157_6, addr_positional[18527:18524], addr_4631_7);

wire[31:0] addr_4632_7;

Selector_2 s4632_7(wires_1158_6[0], addr_1158_6, addr_positional[18531:18528], addr_4632_7);

wire[31:0] addr_4633_7;

Selector_2 s4633_7(wires_1158_6[1], addr_1158_6, addr_positional[18535:18532], addr_4633_7);

wire[31:0] addr_4634_7;

Selector_2 s4634_7(wires_1158_6[2], addr_1158_6, addr_positional[18539:18536], addr_4634_7);

wire[31:0] addr_4635_7;

Selector_2 s4635_7(wires_1158_6[3], addr_1158_6, addr_positional[18543:18540], addr_4635_7);

wire[31:0] addr_4636_7;

Selector_2 s4636_7(wires_1159_6[0], addr_1159_6, addr_positional[18547:18544], addr_4636_7);

wire[31:0] addr_4637_7;

Selector_2 s4637_7(wires_1159_6[1], addr_1159_6, addr_positional[18551:18548], addr_4637_7);

wire[31:0] addr_4638_7;

Selector_2 s4638_7(wires_1159_6[2], addr_1159_6, addr_positional[18555:18552], addr_4638_7);

wire[31:0] addr_4639_7;

Selector_2 s4639_7(wires_1159_6[3], addr_1159_6, addr_positional[18559:18556], addr_4639_7);

wire[31:0] addr_4640_7;

Selector_2 s4640_7(wires_1160_6[0], addr_1160_6, addr_positional[18563:18560], addr_4640_7);

wire[31:0] addr_4641_7;

Selector_2 s4641_7(wires_1160_6[1], addr_1160_6, addr_positional[18567:18564], addr_4641_7);

wire[31:0] addr_4642_7;

Selector_2 s4642_7(wires_1160_6[2], addr_1160_6, addr_positional[18571:18568], addr_4642_7);

wire[31:0] addr_4643_7;

Selector_2 s4643_7(wires_1160_6[3], addr_1160_6, addr_positional[18575:18572], addr_4643_7);

wire[31:0] addr_4644_7;

Selector_2 s4644_7(wires_1161_6[0], addr_1161_6, addr_positional[18579:18576], addr_4644_7);

wire[31:0] addr_4645_7;

Selector_2 s4645_7(wires_1161_6[1], addr_1161_6, addr_positional[18583:18580], addr_4645_7);

wire[31:0] addr_4646_7;

Selector_2 s4646_7(wires_1161_6[2], addr_1161_6, addr_positional[18587:18584], addr_4646_7);

wire[31:0] addr_4647_7;

Selector_2 s4647_7(wires_1161_6[3], addr_1161_6, addr_positional[18591:18588], addr_4647_7);

wire[31:0] addr_4648_7;

Selector_2 s4648_7(wires_1162_6[0], addr_1162_6, addr_positional[18595:18592], addr_4648_7);

wire[31:0] addr_4649_7;

Selector_2 s4649_7(wires_1162_6[1], addr_1162_6, addr_positional[18599:18596], addr_4649_7);

wire[31:0] addr_4650_7;

Selector_2 s4650_7(wires_1162_6[2], addr_1162_6, addr_positional[18603:18600], addr_4650_7);

wire[31:0] addr_4651_7;

Selector_2 s4651_7(wires_1162_6[3], addr_1162_6, addr_positional[18607:18604], addr_4651_7);

wire[31:0] addr_4652_7;

Selector_2 s4652_7(wires_1163_6[0], addr_1163_6, addr_positional[18611:18608], addr_4652_7);

wire[31:0] addr_4653_7;

Selector_2 s4653_7(wires_1163_6[1], addr_1163_6, addr_positional[18615:18612], addr_4653_7);

wire[31:0] addr_4654_7;

Selector_2 s4654_7(wires_1163_6[2], addr_1163_6, addr_positional[18619:18616], addr_4654_7);

wire[31:0] addr_4655_7;

Selector_2 s4655_7(wires_1163_6[3], addr_1163_6, addr_positional[18623:18620], addr_4655_7);

wire[31:0] addr_4656_7;

Selector_2 s4656_7(wires_1164_6[0], addr_1164_6, addr_positional[18627:18624], addr_4656_7);

wire[31:0] addr_4657_7;

Selector_2 s4657_7(wires_1164_6[1], addr_1164_6, addr_positional[18631:18628], addr_4657_7);

wire[31:0] addr_4658_7;

Selector_2 s4658_7(wires_1164_6[2], addr_1164_6, addr_positional[18635:18632], addr_4658_7);

wire[31:0] addr_4659_7;

Selector_2 s4659_7(wires_1164_6[3], addr_1164_6, addr_positional[18639:18636], addr_4659_7);

wire[31:0] addr_4660_7;

Selector_2 s4660_7(wires_1165_6[0], addr_1165_6, addr_positional[18643:18640], addr_4660_7);

wire[31:0] addr_4661_7;

Selector_2 s4661_7(wires_1165_6[1], addr_1165_6, addr_positional[18647:18644], addr_4661_7);

wire[31:0] addr_4662_7;

Selector_2 s4662_7(wires_1165_6[2], addr_1165_6, addr_positional[18651:18648], addr_4662_7);

wire[31:0] addr_4663_7;

Selector_2 s4663_7(wires_1165_6[3], addr_1165_6, addr_positional[18655:18652], addr_4663_7);

wire[31:0] addr_4664_7;

Selector_2 s4664_7(wires_1166_6[0], addr_1166_6, addr_positional[18659:18656], addr_4664_7);

wire[31:0] addr_4665_7;

Selector_2 s4665_7(wires_1166_6[1], addr_1166_6, addr_positional[18663:18660], addr_4665_7);

wire[31:0] addr_4666_7;

Selector_2 s4666_7(wires_1166_6[2], addr_1166_6, addr_positional[18667:18664], addr_4666_7);

wire[31:0] addr_4667_7;

Selector_2 s4667_7(wires_1166_6[3], addr_1166_6, addr_positional[18671:18668], addr_4667_7);

wire[31:0] addr_4668_7;

Selector_2 s4668_7(wires_1167_6[0], addr_1167_6, addr_positional[18675:18672], addr_4668_7);

wire[31:0] addr_4669_7;

Selector_2 s4669_7(wires_1167_6[1], addr_1167_6, addr_positional[18679:18676], addr_4669_7);

wire[31:0] addr_4670_7;

Selector_2 s4670_7(wires_1167_6[2], addr_1167_6, addr_positional[18683:18680], addr_4670_7);

wire[31:0] addr_4671_7;

Selector_2 s4671_7(wires_1167_6[3], addr_1167_6, addr_positional[18687:18684], addr_4671_7);

wire[31:0] addr_4672_7;

Selector_2 s4672_7(wires_1168_6[0], addr_1168_6, addr_positional[18691:18688], addr_4672_7);

wire[31:0] addr_4673_7;

Selector_2 s4673_7(wires_1168_6[1], addr_1168_6, addr_positional[18695:18692], addr_4673_7);

wire[31:0] addr_4674_7;

Selector_2 s4674_7(wires_1168_6[2], addr_1168_6, addr_positional[18699:18696], addr_4674_7);

wire[31:0] addr_4675_7;

Selector_2 s4675_7(wires_1168_6[3], addr_1168_6, addr_positional[18703:18700], addr_4675_7);

wire[31:0] addr_4676_7;

Selector_2 s4676_7(wires_1169_6[0], addr_1169_6, addr_positional[18707:18704], addr_4676_7);

wire[31:0] addr_4677_7;

Selector_2 s4677_7(wires_1169_6[1], addr_1169_6, addr_positional[18711:18708], addr_4677_7);

wire[31:0] addr_4678_7;

Selector_2 s4678_7(wires_1169_6[2], addr_1169_6, addr_positional[18715:18712], addr_4678_7);

wire[31:0] addr_4679_7;

Selector_2 s4679_7(wires_1169_6[3], addr_1169_6, addr_positional[18719:18716], addr_4679_7);

wire[31:0] addr_4680_7;

Selector_2 s4680_7(wires_1170_6[0], addr_1170_6, addr_positional[18723:18720], addr_4680_7);

wire[31:0] addr_4681_7;

Selector_2 s4681_7(wires_1170_6[1], addr_1170_6, addr_positional[18727:18724], addr_4681_7);

wire[31:0] addr_4682_7;

Selector_2 s4682_7(wires_1170_6[2], addr_1170_6, addr_positional[18731:18728], addr_4682_7);

wire[31:0] addr_4683_7;

Selector_2 s4683_7(wires_1170_6[3], addr_1170_6, addr_positional[18735:18732], addr_4683_7);

wire[31:0] addr_4684_7;

Selector_2 s4684_7(wires_1171_6[0], addr_1171_6, addr_positional[18739:18736], addr_4684_7);

wire[31:0] addr_4685_7;

Selector_2 s4685_7(wires_1171_6[1], addr_1171_6, addr_positional[18743:18740], addr_4685_7);

wire[31:0] addr_4686_7;

Selector_2 s4686_7(wires_1171_6[2], addr_1171_6, addr_positional[18747:18744], addr_4686_7);

wire[31:0] addr_4687_7;

Selector_2 s4687_7(wires_1171_6[3], addr_1171_6, addr_positional[18751:18748], addr_4687_7);

wire[31:0] addr_4688_7;

Selector_2 s4688_7(wires_1172_6[0], addr_1172_6, addr_positional[18755:18752], addr_4688_7);

wire[31:0] addr_4689_7;

Selector_2 s4689_7(wires_1172_6[1], addr_1172_6, addr_positional[18759:18756], addr_4689_7);

wire[31:0] addr_4690_7;

Selector_2 s4690_7(wires_1172_6[2], addr_1172_6, addr_positional[18763:18760], addr_4690_7);

wire[31:0] addr_4691_7;

Selector_2 s4691_7(wires_1172_6[3], addr_1172_6, addr_positional[18767:18764], addr_4691_7);

wire[31:0] addr_4692_7;

Selector_2 s4692_7(wires_1173_6[0], addr_1173_6, addr_positional[18771:18768], addr_4692_7);

wire[31:0] addr_4693_7;

Selector_2 s4693_7(wires_1173_6[1], addr_1173_6, addr_positional[18775:18772], addr_4693_7);

wire[31:0] addr_4694_7;

Selector_2 s4694_7(wires_1173_6[2], addr_1173_6, addr_positional[18779:18776], addr_4694_7);

wire[31:0] addr_4695_7;

Selector_2 s4695_7(wires_1173_6[3], addr_1173_6, addr_positional[18783:18780], addr_4695_7);

wire[31:0] addr_4696_7;

Selector_2 s4696_7(wires_1174_6[0], addr_1174_6, addr_positional[18787:18784], addr_4696_7);

wire[31:0] addr_4697_7;

Selector_2 s4697_7(wires_1174_6[1], addr_1174_6, addr_positional[18791:18788], addr_4697_7);

wire[31:0] addr_4698_7;

Selector_2 s4698_7(wires_1174_6[2], addr_1174_6, addr_positional[18795:18792], addr_4698_7);

wire[31:0] addr_4699_7;

Selector_2 s4699_7(wires_1174_6[3], addr_1174_6, addr_positional[18799:18796], addr_4699_7);

wire[31:0] addr_4700_7;

Selector_2 s4700_7(wires_1175_6[0], addr_1175_6, addr_positional[18803:18800], addr_4700_7);

wire[31:0] addr_4701_7;

Selector_2 s4701_7(wires_1175_6[1], addr_1175_6, addr_positional[18807:18804], addr_4701_7);

wire[31:0] addr_4702_7;

Selector_2 s4702_7(wires_1175_6[2], addr_1175_6, addr_positional[18811:18808], addr_4702_7);

wire[31:0] addr_4703_7;

Selector_2 s4703_7(wires_1175_6[3], addr_1175_6, addr_positional[18815:18812], addr_4703_7);

wire[31:0] addr_4704_7;

Selector_2 s4704_7(wires_1176_6[0], addr_1176_6, addr_positional[18819:18816], addr_4704_7);

wire[31:0] addr_4705_7;

Selector_2 s4705_7(wires_1176_6[1], addr_1176_6, addr_positional[18823:18820], addr_4705_7);

wire[31:0] addr_4706_7;

Selector_2 s4706_7(wires_1176_6[2], addr_1176_6, addr_positional[18827:18824], addr_4706_7);

wire[31:0] addr_4707_7;

Selector_2 s4707_7(wires_1176_6[3], addr_1176_6, addr_positional[18831:18828], addr_4707_7);

wire[31:0] addr_4708_7;

Selector_2 s4708_7(wires_1177_6[0], addr_1177_6, addr_positional[18835:18832], addr_4708_7);

wire[31:0] addr_4709_7;

Selector_2 s4709_7(wires_1177_6[1], addr_1177_6, addr_positional[18839:18836], addr_4709_7);

wire[31:0] addr_4710_7;

Selector_2 s4710_7(wires_1177_6[2], addr_1177_6, addr_positional[18843:18840], addr_4710_7);

wire[31:0] addr_4711_7;

Selector_2 s4711_7(wires_1177_6[3], addr_1177_6, addr_positional[18847:18844], addr_4711_7);

wire[31:0] addr_4712_7;

Selector_2 s4712_7(wires_1178_6[0], addr_1178_6, addr_positional[18851:18848], addr_4712_7);

wire[31:0] addr_4713_7;

Selector_2 s4713_7(wires_1178_6[1], addr_1178_6, addr_positional[18855:18852], addr_4713_7);

wire[31:0] addr_4714_7;

Selector_2 s4714_7(wires_1178_6[2], addr_1178_6, addr_positional[18859:18856], addr_4714_7);

wire[31:0] addr_4715_7;

Selector_2 s4715_7(wires_1178_6[3], addr_1178_6, addr_positional[18863:18860], addr_4715_7);

wire[31:0] addr_4716_7;

Selector_2 s4716_7(wires_1179_6[0], addr_1179_6, addr_positional[18867:18864], addr_4716_7);

wire[31:0] addr_4717_7;

Selector_2 s4717_7(wires_1179_6[1], addr_1179_6, addr_positional[18871:18868], addr_4717_7);

wire[31:0] addr_4718_7;

Selector_2 s4718_7(wires_1179_6[2], addr_1179_6, addr_positional[18875:18872], addr_4718_7);

wire[31:0] addr_4719_7;

Selector_2 s4719_7(wires_1179_6[3], addr_1179_6, addr_positional[18879:18876], addr_4719_7);

wire[31:0] addr_4720_7;

Selector_2 s4720_7(wires_1180_6[0], addr_1180_6, addr_positional[18883:18880], addr_4720_7);

wire[31:0] addr_4721_7;

Selector_2 s4721_7(wires_1180_6[1], addr_1180_6, addr_positional[18887:18884], addr_4721_7);

wire[31:0] addr_4722_7;

Selector_2 s4722_7(wires_1180_6[2], addr_1180_6, addr_positional[18891:18888], addr_4722_7);

wire[31:0] addr_4723_7;

Selector_2 s4723_7(wires_1180_6[3], addr_1180_6, addr_positional[18895:18892], addr_4723_7);

wire[31:0] addr_4724_7;

Selector_2 s4724_7(wires_1181_6[0], addr_1181_6, addr_positional[18899:18896], addr_4724_7);

wire[31:0] addr_4725_7;

Selector_2 s4725_7(wires_1181_6[1], addr_1181_6, addr_positional[18903:18900], addr_4725_7);

wire[31:0] addr_4726_7;

Selector_2 s4726_7(wires_1181_6[2], addr_1181_6, addr_positional[18907:18904], addr_4726_7);

wire[31:0] addr_4727_7;

Selector_2 s4727_7(wires_1181_6[3], addr_1181_6, addr_positional[18911:18908], addr_4727_7);

wire[31:0] addr_4728_7;

Selector_2 s4728_7(wires_1182_6[0], addr_1182_6, addr_positional[18915:18912], addr_4728_7);

wire[31:0] addr_4729_7;

Selector_2 s4729_7(wires_1182_6[1], addr_1182_6, addr_positional[18919:18916], addr_4729_7);

wire[31:0] addr_4730_7;

Selector_2 s4730_7(wires_1182_6[2], addr_1182_6, addr_positional[18923:18920], addr_4730_7);

wire[31:0] addr_4731_7;

Selector_2 s4731_7(wires_1182_6[3], addr_1182_6, addr_positional[18927:18924], addr_4731_7);

wire[31:0] addr_4732_7;

Selector_2 s4732_7(wires_1183_6[0], addr_1183_6, addr_positional[18931:18928], addr_4732_7);

wire[31:0] addr_4733_7;

Selector_2 s4733_7(wires_1183_6[1], addr_1183_6, addr_positional[18935:18932], addr_4733_7);

wire[31:0] addr_4734_7;

Selector_2 s4734_7(wires_1183_6[2], addr_1183_6, addr_positional[18939:18936], addr_4734_7);

wire[31:0] addr_4735_7;

Selector_2 s4735_7(wires_1183_6[3], addr_1183_6, addr_positional[18943:18940], addr_4735_7);

wire[31:0] addr_4736_7;

Selector_2 s4736_7(wires_1184_6[0], addr_1184_6, addr_positional[18947:18944], addr_4736_7);

wire[31:0] addr_4737_7;

Selector_2 s4737_7(wires_1184_6[1], addr_1184_6, addr_positional[18951:18948], addr_4737_7);

wire[31:0] addr_4738_7;

Selector_2 s4738_7(wires_1184_6[2], addr_1184_6, addr_positional[18955:18952], addr_4738_7);

wire[31:0] addr_4739_7;

Selector_2 s4739_7(wires_1184_6[3], addr_1184_6, addr_positional[18959:18956], addr_4739_7);

wire[31:0] addr_4740_7;

Selector_2 s4740_7(wires_1185_6[0], addr_1185_6, addr_positional[18963:18960], addr_4740_7);

wire[31:0] addr_4741_7;

Selector_2 s4741_7(wires_1185_6[1], addr_1185_6, addr_positional[18967:18964], addr_4741_7);

wire[31:0] addr_4742_7;

Selector_2 s4742_7(wires_1185_6[2], addr_1185_6, addr_positional[18971:18968], addr_4742_7);

wire[31:0] addr_4743_7;

Selector_2 s4743_7(wires_1185_6[3], addr_1185_6, addr_positional[18975:18972], addr_4743_7);

wire[31:0] addr_4744_7;

Selector_2 s4744_7(wires_1186_6[0], addr_1186_6, addr_positional[18979:18976], addr_4744_7);

wire[31:0] addr_4745_7;

Selector_2 s4745_7(wires_1186_6[1], addr_1186_6, addr_positional[18983:18980], addr_4745_7);

wire[31:0] addr_4746_7;

Selector_2 s4746_7(wires_1186_6[2], addr_1186_6, addr_positional[18987:18984], addr_4746_7);

wire[31:0] addr_4747_7;

Selector_2 s4747_7(wires_1186_6[3], addr_1186_6, addr_positional[18991:18988], addr_4747_7);

wire[31:0] addr_4748_7;

Selector_2 s4748_7(wires_1187_6[0], addr_1187_6, addr_positional[18995:18992], addr_4748_7);

wire[31:0] addr_4749_7;

Selector_2 s4749_7(wires_1187_6[1], addr_1187_6, addr_positional[18999:18996], addr_4749_7);

wire[31:0] addr_4750_7;

Selector_2 s4750_7(wires_1187_6[2], addr_1187_6, addr_positional[19003:19000], addr_4750_7);

wire[31:0] addr_4751_7;

Selector_2 s4751_7(wires_1187_6[3], addr_1187_6, addr_positional[19007:19004], addr_4751_7);

wire[31:0] addr_4752_7;

Selector_2 s4752_7(wires_1188_6[0], addr_1188_6, addr_positional[19011:19008], addr_4752_7);

wire[31:0] addr_4753_7;

Selector_2 s4753_7(wires_1188_6[1], addr_1188_6, addr_positional[19015:19012], addr_4753_7);

wire[31:0] addr_4754_7;

Selector_2 s4754_7(wires_1188_6[2], addr_1188_6, addr_positional[19019:19016], addr_4754_7);

wire[31:0] addr_4755_7;

Selector_2 s4755_7(wires_1188_6[3], addr_1188_6, addr_positional[19023:19020], addr_4755_7);

wire[31:0] addr_4756_7;

Selector_2 s4756_7(wires_1189_6[0], addr_1189_6, addr_positional[19027:19024], addr_4756_7);

wire[31:0] addr_4757_7;

Selector_2 s4757_7(wires_1189_6[1], addr_1189_6, addr_positional[19031:19028], addr_4757_7);

wire[31:0] addr_4758_7;

Selector_2 s4758_7(wires_1189_6[2], addr_1189_6, addr_positional[19035:19032], addr_4758_7);

wire[31:0] addr_4759_7;

Selector_2 s4759_7(wires_1189_6[3], addr_1189_6, addr_positional[19039:19036], addr_4759_7);

wire[31:0] addr_4760_7;

Selector_2 s4760_7(wires_1190_6[0], addr_1190_6, addr_positional[19043:19040], addr_4760_7);

wire[31:0] addr_4761_7;

Selector_2 s4761_7(wires_1190_6[1], addr_1190_6, addr_positional[19047:19044], addr_4761_7);

wire[31:0] addr_4762_7;

Selector_2 s4762_7(wires_1190_6[2], addr_1190_6, addr_positional[19051:19048], addr_4762_7);

wire[31:0] addr_4763_7;

Selector_2 s4763_7(wires_1190_6[3], addr_1190_6, addr_positional[19055:19052], addr_4763_7);

wire[31:0] addr_4764_7;

Selector_2 s4764_7(wires_1191_6[0], addr_1191_6, addr_positional[19059:19056], addr_4764_7);

wire[31:0] addr_4765_7;

Selector_2 s4765_7(wires_1191_6[1], addr_1191_6, addr_positional[19063:19060], addr_4765_7);

wire[31:0] addr_4766_7;

Selector_2 s4766_7(wires_1191_6[2], addr_1191_6, addr_positional[19067:19064], addr_4766_7);

wire[31:0] addr_4767_7;

Selector_2 s4767_7(wires_1191_6[3], addr_1191_6, addr_positional[19071:19068], addr_4767_7);

wire[31:0] addr_4768_7;

Selector_2 s4768_7(wires_1192_6[0], addr_1192_6, addr_positional[19075:19072], addr_4768_7);

wire[31:0] addr_4769_7;

Selector_2 s4769_7(wires_1192_6[1], addr_1192_6, addr_positional[19079:19076], addr_4769_7);

wire[31:0] addr_4770_7;

Selector_2 s4770_7(wires_1192_6[2], addr_1192_6, addr_positional[19083:19080], addr_4770_7);

wire[31:0] addr_4771_7;

Selector_2 s4771_7(wires_1192_6[3], addr_1192_6, addr_positional[19087:19084], addr_4771_7);

wire[31:0] addr_4772_7;

Selector_2 s4772_7(wires_1193_6[0], addr_1193_6, addr_positional[19091:19088], addr_4772_7);

wire[31:0] addr_4773_7;

Selector_2 s4773_7(wires_1193_6[1], addr_1193_6, addr_positional[19095:19092], addr_4773_7);

wire[31:0] addr_4774_7;

Selector_2 s4774_7(wires_1193_6[2], addr_1193_6, addr_positional[19099:19096], addr_4774_7);

wire[31:0] addr_4775_7;

Selector_2 s4775_7(wires_1193_6[3], addr_1193_6, addr_positional[19103:19100], addr_4775_7);

wire[31:0] addr_4776_7;

Selector_2 s4776_7(wires_1194_6[0], addr_1194_6, addr_positional[19107:19104], addr_4776_7);

wire[31:0] addr_4777_7;

Selector_2 s4777_7(wires_1194_6[1], addr_1194_6, addr_positional[19111:19108], addr_4777_7);

wire[31:0] addr_4778_7;

Selector_2 s4778_7(wires_1194_6[2], addr_1194_6, addr_positional[19115:19112], addr_4778_7);

wire[31:0] addr_4779_7;

Selector_2 s4779_7(wires_1194_6[3], addr_1194_6, addr_positional[19119:19116], addr_4779_7);

wire[31:0] addr_4780_7;

Selector_2 s4780_7(wires_1195_6[0], addr_1195_6, addr_positional[19123:19120], addr_4780_7);

wire[31:0] addr_4781_7;

Selector_2 s4781_7(wires_1195_6[1], addr_1195_6, addr_positional[19127:19124], addr_4781_7);

wire[31:0] addr_4782_7;

Selector_2 s4782_7(wires_1195_6[2], addr_1195_6, addr_positional[19131:19128], addr_4782_7);

wire[31:0] addr_4783_7;

Selector_2 s4783_7(wires_1195_6[3], addr_1195_6, addr_positional[19135:19132], addr_4783_7);

wire[31:0] addr_4784_7;

Selector_2 s4784_7(wires_1196_6[0], addr_1196_6, addr_positional[19139:19136], addr_4784_7);

wire[31:0] addr_4785_7;

Selector_2 s4785_7(wires_1196_6[1], addr_1196_6, addr_positional[19143:19140], addr_4785_7);

wire[31:0] addr_4786_7;

Selector_2 s4786_7(wires_1196_6[2], addr_1196_6, addr_positional[19147:19144], addr_4786_7);

wire[31:0] addr_4787_7;

Selector_2 s4787_7(wires_1196_6[3], addr_1196_6, addr_positional[19151:19148], addr_4787_7);

wire[31:0] addr_4788_7;

Selector_2 s4788_7(wires_1197_6[0], addr_1197_6, addr_positional[19155:19152], addr_4788_7);

wire[31:0] addr_4789_7;

Selector_2 s4789_7(wires_1197_6[1], addr_1197_6, addr_positional[19159:19156], addr_4789_7);

wire[31:0] addr_4790_7;

Selector_2 s4790_7(wires_1197_6[2], addr_1197_6, addr_positional[19163:19160], addr_4790_7);

wire[31:0] addr_4791_7;

Selector_2 s4791_7(wires_1197_6[3], addr_1197_6, addr_positional[19167:19164], addr_4791_7);

wire[31:0] addr_4792_7;

Selector_2 s4792_7(wires_1198_6[0], addr_1198_6, addr_positional[19171:19168], addr_4792_7);

wire[31:0] addr_4793_7;

Selector_2 s4793_7(wires_1198_6[1], addr_1198_6, addr_positional[19175:19172], addr_4793_7);

wire[31:0] addr_4794_7;

Selector_2 s4794_7(wires_1198_6[2], addr_1198_6, addr_positional[19179:19176], addr_4794_7);

wire[31:0] addr_4795_7;

Selector_2 s4795_7(wires_1198_6[3], addr_1198_6, addr_positional[19183:19180], addr_4795_7);

wire[31:0] addr_4796_7;

Selector_2 s4796_7(wires_1199_6[0], addr_1199_6, addr_positional[19187:19184], addr_4796_7);

wire[31:0] addr_4797_7;

Selector_2 s4797_7(wires_1199_6[1], addr_1199_6, addr_positional[19191:19188], addr_4797_7);

wire[31:0] addr_4798_7;

Selector_2 s4798_7(wires_1199_6[2], addr_1199_6, addr_positional[19195:19192], addr_4798_7);

wire[31:0] addr_4799_7;

Selector_2 s4799_7(wires_1199_6[3], addr_1199_6, addr_positional[19199:19196], addr_4799_7);

wire[31:0] addr_4800_7;

Selector_2 s4800_7(wires_1200_6[0], addr_1200_6, addr_positional[19203:19200], addr_4800_7);

wire[31:0] addr_4801_7;

Selector_2 s4801_7(wires_1200_6[1], addr_1200_6, addr_positional[19207:19204], addr_4801_7);

wire[31:0] addr_4802_7;

Selector_2 s4802_7(wires_1200_6[2], addr_1200_6, addr_positional[19211:19208], addr_4802_7);

wire[31:0] addr_4803_7;

Selector_2 s4803_7(wires_1200_6[3], addr_1200_6, addr_positional[19215:19212], addr_4803_7);

wire[31:0] addr_4804_7;

Selector_2 s4804_7(wires_1201_6[0], addr_1201_6, addr_positional[19219:19216], addr_4804_7);

wire[31:0] addr_4805_7;

Selector_2 s4805_7(wires_1201_6[1], addr_1201_6, addr_positional[19223:19220], addr_4805_7);

wire[31:0] addr_4806_7;

Selector_2 s4806_7(wires_1201_6[2], addr_1201_6, addr_positional[19227:19224], addr_4806_7);

wire[31:0] addr_4807_7;

Selector_2 s4807_7(wires_1201_6[3], addr_1201_6, addr_positional[19231:19228], addr_4807_7);

wire[31:0] addr_4808_7;

Selector_2 s4808_7(wires_1202_6[0], addr_1202_6, addr_positional[19235:19232], addr_4808_7);

wire[31:0] addr_4809_7;

Selector_2 s4809_7(wires_1202_6[1], addr_1202_6, addr_positional[19239:19236], addr_4809_7);

wire[31:0] addr_4810_7;

Selector_2 s4810_7(wires_1202_6[2], addr_1202_6, addr_positional[19243:19240], addr_4810_7);

wire[31:0] addr_4811_7;

Selector_2 s4811_7(wires_1202_6[3], addr_1202_6, addr_positional[19247:19244], addr_4811_7);

wire[31:0] addr_4812_7;

Selector_2 s4812_7(wires_1203_6[0], addr_1203_6, addr_positional[19251:19248], addr_4812_7);

wire[31:0] addr_4813_7;

Selector_2 s4813_7(wires_1203_6[1], addr_1203_6, addr_positional[19255:19252], addr_4813_7);

wire[31:0] addr_4814_7;

Selector_2 s4814_7(wires_1203_6[2], addr_1203_6, addr_positional[19259:19256], addr_4814_7);

wire[31:0] addr_4815_7;

Selector_2 s4815_7(wires_1203_6[3], addr_1203_6, addr_positional[19263:19260], addr_4815_7);

wire[31:0] addr_4816_7;

Selector_2 s4816_7(wires_1204_6[0], addr_1204_6, addr_positional[19267:19264], addr_4816_7);

wire[31:0] addr_4817_7;

Selector_2 s4817_7(wires_1204_6[1], addr_1204_6, addr_positional[19271:19268], addr_4817_7);

wire[31:0] addr_4818_7;

Selector_2 s4818_7(wires_1204_6[2], addr_1204_6, addr_positional[19275:19272], addr_4818_7);

wire[31:0] addr_4819_7;

Selector_2 s4819_7(wires_1204_6[3], addr_1204_6, addr_positional[19279:19276], addr_4819_7);

wire[31:0] addr_4820_7;

Selector_2 s4820_7(wires_1205_6[0], addr_1205_6, addr_positional[19283:19280], addr_4820_7);

wire[31:0] addr_4821_7;

Selector_2 s4821_7(wires_1205_6[1], addr_1205_6, addr_positional[19287:19284], addr_4821_7);

wire[31:0] addr_4822_7;

Selector_2 s4822_7(wires_1205_6[2], addr_1205_6, addr_positional[19291:19288], addr_4822_7);

wire[31:0] addr_4823_7;

Selector_2 s4823_7(wires_1205_6[3], addr_1205_6, addr_positional[19295:19292], addr_4823_7);

wire[31:0] addr_4824_7;

Selector_2 s4824_7(wires_1206_6[0], addr_1206_6, addr_positional[19299:19296], addr_4824_7);

wire[31:0] addr_4825_7;

Selector_2 s4825_7(wires_1206_6[1], addr_1206_6, addr_positional[19303:19300], addr_4825_7);

wire[31:0] addr_4826_7;

Selector_2 s4826_7(wires_1206_6[2], addr_1206_6, addr_positional[19307:19304], addr_4826_7);

wire[31:0] addr_4827_7;

Selector_2 s4827_7(wires_1206_6[3], addr_1206_6, addr_positional[19311:19308], addr_4827_7);

wire[31:0] addr_4828_7;

Selector_2 s4828_7(wires_1207_6[0], addr_1207_6, addr_positional[19315:19312], addr_4828_7);

wire[31:0] addr_4829_7;

Selector_2 s4829_7(wires_1207_6[1], addr_1207_6, addr_positional[19319:19316], addr_4829_7);

wire[31:0] addr_4830_7;

Selector_2 s4830_7(wires_1207_6[2], addr_1207_6, addr_positional[19323:19320], addr_4830_7);

wire[31:0] addr_4831_7;

Selector_2 s4831_7(wires_1207_6[3], addr_1207_6, addr_positional[19327:19324], addr_4831_7);

wire[31:0] addr_4832_7;

Selector_2 s4832_7(wires_1208_6[0], addr_1208_6, addr_positional[19331:19328], addr_4832_7);

wire[31:0] addr_4833_7;

Selector_2 s4833_7(wires_1208_6[1], addr_1208_6, addr_positional[19335:19332], addr_4833_7);

wire[31:0] addr_4834_7;

Selector_2 s4834_7(wires_1208_6[2], addr_1208_6, addr_positional[19339:19336], addr_4834_7);

wire[31:0] addr_4835_7;

Selector_2 s4835_7(wires_1208_6[3], addr_1208_6, addr_positional[19343:19340], addr_4835_7);

wire[31:0] addr_4836_7;

Selector_2 s4836_7(wires_1209_6[0], addr_1209_6, addr_positional[19347:19344], addr_4836_7);

wire[31:0] addr_4837_7;

Selector_2 s4837_7(wires_1209_6[1], addr_1209_6, addr_positional[19351:19348], addr_4837_7);

wire[31:0] addr_4838_7;

Selector_2 s4838_7(wires_1209_6[2], addr_1209_6, addr_positional[19355:19352], addr_4838_7);

wire[31:0] addr_4839_7;

Selector_2 s4839_7(wires_1209_6[3], addr_1209_6, addr_positional[19359:19356], addr_4839_7);

wire[31:0] addr_4840_7;

Selector_2 s4840_7(wires_1210_6[0], addr_1210_6, addr_positional[19363:19360], addr_4840_7);

wire[31:0] addr_4841_7;

Selector_2 s4841_7(wires_1210_6[1], addr_1210_6, addr_positional[19367:19364], addr_4841_7);

wire[31:0] addr_4842_7;

Selector_2 s4842_7(wires_1210_6[2], addr_1210_6, addr_positional[19371:19368], addr_4842_7);

wire[31:0] addr_4843_7;

Selector_2 s4843_7(wires_1210_6[3], addr_1210_6, addr_positional[19375:19372], addr_4843_7);

wire[31:0] addr_4844_7;

Selector_2 s4844_7(wires_1211_6[0], addr_1211_6, addr_positional[19379:19376], addr_4844_7);

wire[31:0] addr_4845_7;

Selector_2 s4845_7(wires_1211_6[1], addr_1211_6, addr_positional[19383:19380], addr_4845_7);

wire[31:0] addr_4846_7;

Selector_2 s4846_7(wires_1211_6[2], addr_1211_6, addr_positional[19387:19384], addr_4846_7);

wire[31:0] addr_4847_7;

Selector_2 s4847_7(wires_1211_6[3], addr_1211_6, addr_positional[19391:19388], addr_4847_7);

wire[31:0] addr_4848_7;

Selector_2 s4848_7(wires_1212_6[0], addr_1212_6, addr_positional[19395:19392], addr_4848_7);

wire[31:0] addr_4849_7;

Selector_2 s4849_7(wires_1212_6[1], addr_1212_6, addr_positional[19399:19396], addr_4849_7);

wire[31:0] addr_4850_7;

Selector_2 s4850_7(wires_1212_6[2], addr_1212_6, addr_positional[19403:19400], addr_4850_7);

wire[31:0] addr_4851_7;

Selector_2 s4851_7(wires_1212_6[3], addr_1212_6, addr_positional[19407:19404], addr_4851_7);

wire[31:0] addr_4852_7;

Selector_2 s4852_7(wires_1213_6[0], addr_1213_6, addr_positional[19411:19408], addr_4852_7);

wire[31:0] addr_4853_7;

Selector_2 s4853_7(wires_1213_6[1], addr_1213_6, addr_positional[19415:19412], addr_4853_7);

wire[31:0] addr_4854_7;

Selector_2 s4854_7(wires_1213_6[2], addr_1213_6, addr_positional[19419:19416], addr_4854_7);

wire[31:0] addr_4855_7;

Selector_2 s4855_7(wires_1213_6[3], addr_1213_6, addr_positional[19423:19420], addr_4855_7);

wire[31:0] addr_4856_7;

Selector_2 s4856_7(wires_1214_6[0], addr_1214_6, addr_positional[19427:19424], addr_4856_7);

wire[31:0] addr_4857_7;

Selector_2 s4857_7(wires_1214_6[1], addr_1214_6, addr_positional[19431:19428], addr_4857_7);

wire[31:0] addr_4858_7;

Selector_2 s4858_7(wires_1214_6[2], addr_1214_6, addr_positional[19435:19432], addr_4858_7);

wire[31:0] addr_4859_7;

Selector_2 s4859_7(wires_1214_6[3], addr_1214_6, addr_positional[19439:19436], addr_4859_7);

wire[31:0] addr_4860_7;

Selector_2 s4860_7(wires_1215_6[0], addr_1215_6, addr_positional[19443:19440], addr_4860_7);

wire[31:0] addr_4861_7;

Selector_2 s4861_7(wires_1215_6[1], addr_1215_6, addr_positional[19447:19444], addr_4861_7);

wire[31:0] addr_4862_7;

Selector_2 s4862_7(wires_1215_6[2], addr_1215_6, addr_positional[19451:19448], addr_4862_7);

wire[31:0] addr_4863_7;

Selector_2 s4863_7(wires_1215_6[3], addr_1215_6, addr_positional[19455:19452], addr_4863_7);

wire[31:0] addr_4864_7;

Selector_2 s4864_7(wires_1216_6[0], addr_1216_6, addr_positional[19459:19456], addr_4864_7);

wire[31:0] addr_4865_7;

Selector_2 s4865_7(wires_1216_6[1], addr_1216_6, addr_positional[19463:19460], addr_4865_7);

wire[31:0] addr_4866_7;

Selector_2 s4866_7(wires_1216_6[2], addr_1216_6, addr_positional[19467:19464], addr_4866_7);

wire[31:0] addr_4867_7;

Selector_2 s4867_7(wires_1216_6[3], addr_1216_6, addr_positional[19471:19468], addr_4867_7);

wire[31:0] addr_4868_7;

Selector_2 s4868_7(wires_1217_6[0], addr_1217_6, addr_positional[19475:19472], addr_4868_7);

wire[31:0] addr_4869_7;

Selector_2 s4869_7(wires_1217_6[1], addr_1217_6, addr_positional[19479:19476], addr_4869_7);

wire[31:0] addr_4870_7;

Selector_2 s4870_7(wires_1217_6[2], addr_1217_6, addr_positional[19483:19480], addr_4870_7);

wire[31:0] addr_4871_7;

Selector_2 s4871_7(wires_1217_6[3], addr_1217_6, addr_positional[19487:19484], addr_4871_7);

wire[31:0] addr_4872_7;

Selector_2 s4872_7(wires_1218_6[0], addr_1218_6, addr_positional[19491:19488], addr_4872_7);

wire[31:0] addr_4873_7;

Selector_2 s4873_7(wires_1218_6[1], addr_1218_6, addr_positional[19495:19492], addr_4873_7);

wire[31:0] addr_4874_7;

Selector_2 s4874_7(wires_1218_6[2], addr_1218_6, addr_positional[19499:19496], addr_4874_7);

wire[31:0] addr_4875_7;

Selector_2 s4875_7(wires_1218_6[3], addr_1218_6, addr_positional[19503:19500], addr_4875_7);

wire[31:0] addr_4876_7;

Selector_2 s4876_7(wires_1219_6[0], addr_1219_6, addr_positional[19507:19504], addr_4876_7);

wire[31:0] addr_4877_7;

Selector_2 s4877_7(wires_1219_6[1], addr_1219_6, addr_positional[19511:19508], addr_4877_7);

wire[31:0] addr_4878_7;

Selector_2 s4878_7(wires_1219_6[2], addr_1219_6, addr_positional[19515:19512], addr_4878_7);

wire[31:0] addr_4879_7;

Selector_2 s4879_7(wires_1219_6[3], addr_1219_6, addr_positional[19519:19516], addr_4879_7);

wire[31:0] addr_4880_7;

Selector_2 s4880_7(wires_1220_6[0], addr_1220_6, addr_positional[19523:19520], addr_4880_7);

wire[31:0] addr_4881_7;

Selector_2 s4881_7(wires_1220_6[1], addr_1220_6, addr_positional[19527:19524], addr_4881_7);

wire[31:0] addr_4882_7;

Selector_2 s4882_7(wires_1220_6[2], addr_1220_6, addr_positional[19531:19528], addr_4882_7);

wire[31:0] addr_4883_7;

Selector_2 s4883_7(wires_1220_6[3], addr_1220_6, addr_positional[19535:19532], addr_4883_7);

wire[31:0] addr_4884_7;

Selector_2 s4884_7(wires_1221_6[0], addr_1221_6, addr_positional[19539:19536], addr_4884_7);

wire[31:0] addr_4885_7;

Selector_2 s4885_7(wires_1221_6[1], addr_1221_6, addr_positional[19543:19540], addr_4885_7);

wire[31:0] addr_4886_7;

Selector_2 s4886_7(wires_1221_6[2], addr_1221_6, addr_positional[19547:19544], addr_4886_7);

wire[31:0] addr_4887_7;

Selector_2 s4887_7(wires_1221_6[3], addr_1221_6, addr_positional[19551:19548], addr_4887_7);

wire[31:0] addr_4888_7;

Selector_2 s4888_7(wires_1222_6[0], addr_1222_6, addr_positional[19555:19552], addr_4888_7);

wire[31:0] addr_4889_7;

Selector_2 s4889_7(wires_1222_6[1], addr_1222_6, addr_positional[19559:19556], addr_4889_7);

wire[31:0] addr_4890_7;

Selector_2 s4890_7(wires_1222_6[2], addr_1222_6, addr_positional[19563:19560], addr_4890_7);

wire[31:0] addr_4891_7;

Selector_2 s4891_7(wires_1222_6[3], addr_1222_6, addr_positional[19567:19564], addr_4891_7);

wire[31:0] addr_4892_7;

Selector_2 s4892_7(wires_1223_6[0], addr_1223_6, addr_positional[19571:19568], addr_4892_7);

wire[31:0] addr_4893_7;

Selector_2 s4893_7(wires_1223_6[1], addr_1223_6, addr_positional[19575:19572], addr_4893_7);

wire[31:0] addr_4894_7;

Selector_2 s4894_7(wires_1223_6[2], addr_1223_6, addr_positional[19579:19576], addr_4894_7);

wire[31:0] addr_4895_7;

Selector_2 s4895_7(wires_1223_6[3], addr_1223_6, addr_positional[19583:19580], addr_4895_7);

wire[31:0] addr_4896_7;

Selector_2 s4896_7(wires_1224_6[0], addr_1224_6, addr_positional[19587:19584], addr_4896_7);

wire[31:0] addr_4897_7;

Selector_2 s4897_7(wires_1224_6[1], addr_1224_6, addr_positional[19591:19588], addr_4897_7);

wire[31:0] addr_4898_7;

Selector_2 s4898_7(wires_1224_6[2], addr_1224_6, addr_positional[19595:19592], addr_4898_7);

wire[31:0] addr_4899_7;

Selector_2 s4899_7(wires_1224_6[3], addr_1224_6, addr_positional[19599:19596], addr_4899_7);

wire[31:0] addr_4900_7;

Selector_2 s4900_7(wires_1225_6[0], addr_1225_6, addr_positional[19603:19600], addr_4900_7);

wire[31:0] addr_4901_7;

Selector_2 s4901_7(wires_1225_6[1], addr_1225_6, addr_positional[19607:19604], addr_4901_7);

wire[31:0] addr_4902_7;

Selector_2 s4902_7(wires_1225_6[2], addr_1225_6, addr_positional[19611:19608], addr_4902_7);

wire[31:0] addr_4903_7;

Selector_2 s4903_7(wires_1225_6[3], addr_1225_6, addr_positional[19615:19612], addr_4903_7);

wire[31:0] addr_4904_7;

Selector_2 s4904_7(wires_1226_6[0], addr_1226_6, addr_positional[19619:19616], addr_4904_7);

wire[31:0] addr_4905_7;

Selector_2 s4905_7(wires_1226_6[1], addr_1226_6, addr_positional[19623:19620], addr_4905_7);

wire[31:0] addr_4906_7;

Selector_2 s4906_7(wires_1226_6[2], addr_1226_6, addr_positional[19627:19624], addr_4906_7);

wire[31:0] addr_4907_7;

Selector_2 s4907_7(wires_1226_6[3], addr_1226_6, addr_positional[19631:19628], addr_4907_7);

wire[31:0] addr_4908_7;

Selector_2 s4908_7(wires_1227_6[0], addr_1227_6, addr_positional[19635:19632], addr_4908_7);

wire[31:0] addr_4909_7;

Selector_2 s4909_7(wires_1227_6[1], addr_1227_6, addr_positional[19639:19636], addr_4909_7);

wire[31:0] addr_4910_7;

Selector_2 s4910_7(wires_1227_6[2], addr_1227_6, addr_positional[19643:19640], addr_4910_7);

wire[31:0] addr_4911_7;

Selector_2 s4911_7(wires_1227_6[3], addr_1227_6, addr_positional[19647:19644], addr_4911_7);

wire[31:0] addr_4912_7;

Selector_2 s4912_7(wires_1228_6[0], addr_1228_6, addr_positional[19651:19648], addr_4912_7);

wire[31:0] addr_4913_7;

Selector_2 s4913_7(wires_1228_6[1], addr_1228_6, addr_positional[19655:19652], addr_4913_7);

wire[31:0] addr_4914_7;

Selector_2 s4914_7(wires_1228_6[2], addr_1228_6, addr_positional[19659:19656], addr_4914_7);

wire[31:0] addr_4915_7;

Selector_2 s4915_7(wires_1228_6[3], addr_1228_6, addr_positional[19663:19660], addr_4915_7);

wire[31:0] addr_4916_7;

Selector_2 s4916_7(wires_1229_6[0], addr_1229_6, addr_positional[19667:19664], addr_4916_7);

wire[31:0] addr_4917_7;

Selector_2 s4917_7(wires_1229_6[1], addr_1229_6, addr_positional[19671:19668], addr_4917_7);

wire[31:0] addr_4918_7;

Selector_2 s4918_7(wires_1229_6[2], addr_1229_6, addr_positional[19675:19672], addr_4918_7);

wire[31:0] addr_4919_7;

Selector_2 s4919_7(wires_1229_6[3], addr_1229_6, addr_positional[19679:19676], addr_4919_7);

wire[31:0] addr_4920_7;

Selector_2 s4920_7(wires_1230_6[0], addr_1230_6, addr_positional[19683:19680], addr_4920_7);

wire[31:0] addr_4921_7;

Selector_2 s4921_7(wires_1230_6[1], addr_1230_6, addr_positional[19687:19684], addr_4921_7);

wire[31:0] addr_4922_7;

Selector_2 s4922_7(wires_1230_6[2], addr_1230_6, addr_positional[19691:19688], addr_4922_7);

wire[31:0] addr_4923_7;

Selector_2 s4923_7(wires_1230_6[3], addr_1230_6, addr_positional[19695:19692], addr_4923_7);

wire[31:0] addr_4924_7;

Selector_2 s4924_7(wires_1231_6[0], addr_1231_6, addr_positional[19699:19696], addr_4924_7);

wire[31:0] addr_4925_7;

Selector_2 s4925_7(wires_1231_6[1], addr_1231_6, addr_positional[19703:19700], addr_4925_7);

wire[31:0] addr_4926_7;

Selector_2 s4926_7(wires_1231_6[2], addr_1231_6, addr_positional[19707:19704], addr_4926_7);

wire[31:0] addr_4927_7;

Selector_2 s4927_7(wires_1231_6[3], addr_1231_6, addr_positional[19711:19708], addr_4927_7);

wire[31:0] addr_4928_7;

Selector_2 s4928_7(wires_1232_6[0], addr_1232_6, addr_positional[19715:19712], addr_4928_7);

wire[31:0] addr_4929_7;

Selector_2 s4929_7(wires_1232_6[1], addr_1232_6, addr_positional[19719:19716], addr_4929_7);

wire[31:0] addr_4930_7;

Selector_2 s4930_7(wires_1232_6[2], addr_1232_6, addr_positional[19723:19720], addr_4930_7);

wire[31:0] addr_4931_7;

Selector_2 s4931_7(wires_1232_6[3], addr_1232_6, addr_positional[19727:19724], addr_4931_7);

wire[31:0] addr_4932_7;

Selector_2 s4932_7(wires_1233_6[0], addr_1233_6, addr_positional[19731:19728], addr_4932_7);

wire[31:0] addr_4933_7;

Selector_2 s4933_7(wires_1233_6[1], addr_1233_6, addr_positional[19735:19732], addr_4933_7);

wire[31:0] addr_4934_7;

Selector_2 s4934_7(wires_1233_6[2], addr_1233_6, addr_positional[19739:19736], addr_4934_7);

wire[31:0] addr_4935_7;

Selector_2 s4935_7(wires_1233_6[3], addr_1233_6, addr_positional[19743:19740], addr_4935_7);

wire[31:0] addr_4936_7;

Selector_2 s4936_7(wires_1234_6[0], addr_1234_6, addr_positional[19747:19744], addr_4936_7);

wire[31:0] addr_4937_7;

Selector_2 s4937_7(wires_1234_6[1], addr_1234_6, addr_positional[19751:19748], addr_4937_7);

wire[31:0] addr_4938_7;

Selector_2 s4938_7(wires_1234_6[2], addr_1234_6, addr_positional[19755:19752], addr_4938_7);

wire[31:0] addr_4939_7;

Selector_2 s4939_7(wires_1234_6[3], addr_1234_6, addr_positional[19759:19756], addr_4939_7);

wire[31:0] addr_4940_7;

Selector_2 s4940_7(wires_1235_6[0], addr_1235_6, addr_positional[19763:19760], addr_4940_7);

wire[31:0] addr_4941_7;

Selector_2 s4941_7(wires_1235_6[1], addr_1235_6, addr_positional[19767:19764], addr_4941_7);

wire[31:0] addr_4942_7;

Selector_2 s4942_7(wires_1235_6[2], addr_1235_6, addr_positional[19771:19768], addr_4942_7);

wire[31:0] addr_4943_7;

Selector_2 s4943_7(wires_1235_6[3], addr_1235_6, addr_positional[19775:19772], addr_4943_7);

wire[31:0] addr_4944_7;

Selector_2 s4944_7(wires_1236_6[0], addr_1236_6, addr_positional[19779:19776], addr_4944_7);

wire[31:0] addr_4945_7;

Selector_2 s4945_7(wires_1236_6[1], addr_1236_6, addr_positional[19783:19780], addr_4945_7);

wire[31:0] addr_4946_7;

Selector_2 s4946_7(wires_1236_6[2], addr_1236_6, addr_positional[19787:19784], addr_4946_7);

wire[31:0] addr_4947_7;

Selector_2 s4947_7(wires_1236_6[3], addr_1236_6, addr_positional[19791:19788], addr_4947_7);

wire[31:0] addr_4948_7;

Selector_2 s4948_7(wires_1237_6[0], addr_1237_6, addr_positional[19795:19792], addr_4948_7);

wire[31:0] addr_4949_7;

Selector_2 s4949_7(wires_1237_6[1], addr_1237_6, addr_positional[19799:19796], addr_4949_7);

wire[31:0] addr_4950_7;

Selector_2 s4950_7(wires_1237_6[2], addr_1237_6, addr_positional[19803:19800], addr_4950_7);

wire[31:0] addr_4951_7;

Selector_2 s4951_7(wires_1237_6[3], addr_1237_6, addr_positional[19807:19804], addr_4951_7);

wire[31:0] addr_4952_7;

Selector_2 s4952_7(wires_1238_6[0], addr_1238_6, addr_positional[19811:19808], addr_4952_7);

wire[31:0] addr_4953_7;

Selector_2 s4953_7(wires_1238_6[1], addr_1238_6, addr_positional[19815:19812], addr_4953_7);

wire[31:0] addr_4954_7;

Selector_2 s4954_7(wires_1238_6[2], addr_1238_6, addr_positional[19819:19816], addr_4954_7);

wire[31:0] addr_4955_7;

Selector_2 s4955_7(wires_1238_6[3], addr_1238_6, addr_positional[19823:19820], addr_4955_7);

wire[31:0] addr_4956_7;

Selector_2 s4956_7(wires_1239_6[0], addr_1239_6, addr_positional[19827:19824], addr_4956_7);

wire[31:0] addr_4957_7;

Selector_2 s4957_7(wires_1239_6[1], addr_1239_6, addr_positional[19831:19828], addr_4957_7);

wire[31:0] addr_4958_7;

Selector_2 s4958_7(wires_1239_6[2], addr_1239_6, addr_positional[19835:19832], addr_4958_7);

wire[31:0] addr_4959_7;

Selector_2 s4959_7(wires_1239_6[3], addr_1239_6, addr_positional[19839:19836], addr_4959_7);

wire[31:0] addr_4960_7;

Selector_2 s4960_7(wires_1240_6[0], addr_1240_6, addr_positional[19843:19840], addr_4960_7);

wire[31:0] addr_4961_7;

Selector_2 s4961_7(wires_1240_6[1], addr_1240_6, addr_positional[19847:19844], addr_4961_7);

wire[31:0] addr_4962_7;

Selector_2 s4962_7(wires_1240_6[2], addr_1240_6, addr_positional[19851:19848], addr_4962_7);

wire[31:0] addr_4963_7;

Selector_2 s4963_7(wires_1240_6[3], addr_1240_6, addr_positional[19855:19852], addr_4963_7);

wire[31:0] addr_4964_7;

Selector_2 s4964_7(wires_1241_6[0], addr_1241_6, addr_positional[19859:19856], addr_4964_7);

wire[31:0] addr_4965_7;

Selector_2 s4965_7(wires_1241_6[1], addr_1241_6, addr_positional[19863:19860], addr_4965_7);

wire[31:0] addr_4966_7;

Selector_2 s4966_7(wires_1241_6[2], addr_1241_6, addr_positional[19867:19864], addr_4966_7);

wire[31:0] addr_4967_7;

Selector_2 s4967_7(wires_1241_6[3], addr_1241_6, addr_positional[19871:19868], addr_4967_7);

wire[31:0] addr_4968_7;

Selector_2 s4968_7(wires_1242_6[0], addr_1242_6, addr_positional[19875:19872], addr_4968_7);

wire[31:0] addr_4969_7;

Selector_2 s4969_7(wires_1242_6[1], addr_1242_6, addr_positional[19879:19876], addr_4969_7);

wire[31:0] addr_4970_7;

Selector_2 s4970_7(wires_1242_6[2], addr_1242_6, addr_positional[19883:19880], addr_4970_7);

wire[31:0] addr_4971_7;

Selector_2 s4971_7(wires_1242_6[3], addr_1242_6, addr_positional[19887:19884], addr_4971_7);

wire[31:0] addr_4972_7;

Selector_2 s4972_7(wires_1243_6[0], addr_1243_6, addr_positional[19891:19888], addr_4972_7);

wire[31:0] addr_4973_7;

Selector_2 s4973_7(wires_1243_6[1], addr_1243_6, addr_positional[19895:19892], addr_4973_7);

wire[31:0] addr_4974_7;

Selector_2 s4974_7(wires_1243_6[2], addr_1243_6, addr_positional[19899:19896], addr_4974_7);

wire[31:0] addr_4975_7;

Selector_2 s4975_7(wires_1243_6[3], addr_1243_6, addr_positional[19903:19900], addr_4975_7);

wire[31:0] addr_4976_7;

Selector_2 s4976_7(wires_1244_6[0], addr_1244_6, addr_positional[19907:19904], addr_4976_7);

wire[31:0] addr_4977_7;

Selector_2 s4977_7(wires_1244_6[1], addr_1244_6, addr_positional[19911:19908], addr_4977_7);

wire[31:0] addr_4978_7;

Selector_2 s4978_7(wires_1244_6[2], addr_1244_6, addr_positional[19915:19912], addr_4978_7);

wire[31:0] addr_4979_7;

Selector_2 s4979_7(wires_1244_6[3], addr_1244_6, addr_positional[19919:19916], addr_4979_7);

wire[31:0] addr_4980_7;

Selector_2 s4980_7(wires_1245_6[0], addr_1245_6, addr_positional[19923:19920], addr_4980_7);

wire[31:0] addr_4981_7;

Selector_2 s4981_7(wires_1245_6[1], addr_1245_6, addr_positional[19927:19924], addr_4981_7);

wire[31:0] addr_4982_7;

Selector_2 s4982_7(wires_1245_6[2], addr_1245_6, addr_positional[19931:19928], addr_4982_7);

wire[31:0] addr_4983_7;

Selector_2 s4983_7(wires_1245_6[3], addr_1245_6, addr_positional[19935:19932], addr_4983_7);

wire[31:0] addr_4984_7;

Selector_2 s4984_7(wires_1246_6[0], addr_1246_6, addr_positional[19939:19936], addr_4984_7);

wire[31:0] addr_4985_7;

Selector_2 s4985_7(wires_1246_6[1], addr_1246_6, addr_positional[19943:19940], addr_4985_7);

wire[31:0] addr_4986_7;

Selector_2 s4986_7(wires_1246_6[2], addr_1246_6, addr_positional[19947:19944], addr_4986_7);

wire[31:0] addr_4987_7;

Selector_2 s4987_7(wires_1246_6[3], addr_1246_6, addr_positional[19951:19948], addr_4987_7);

wire[31:0] addr_4988_7;

Selector_2 s4988_7(wires_1247_6[0], addr_1247_6, addr_positional[19955:19952], addr_4988_7);

wire[31:0] addr_4989_7;

Selector_2 s4989_7(wires_1247_6[1], addr_1247_6, addr_positional[19959:19956], addr_4989_7);

wire[31:0] addr_4990_7;

Selector_2 s4990_7(wires_1247_6[2], addr_1247_6, addr_positional[19963:19960], addr_4990_7);

wire[31:0] addr_4991_7;

Selector_2 s4991_7(wires_1247_6[3], addr_1247_6, addr_positional[19967:19964], addr_4991_7);

wire[31:0] addr_4992_7;

Selector_2 s4992_7(wires_1248_6[0], addr_1248_6, addr_positional[19971:19968], addr_4992_7);

wire[31:0] addr_4993_7;

Selector_2 s4993_7(wires_1248_6[1], addr_1248_6, addr_positional[19975:19972], addr_4993_7);

wire[31:0] addr_4994_7;

Selector_2 s4994_7(wires_1248_6[2], addr_1248_6, addr_positional[19979:19976], addr_4994_7);

wire[31:0] addr_4995_7;

Selector_2 s4995_7(wires_1248_6[3], addr_1248_6, addr_positional[19983:19980], addr_4995_7);

wire[31:0] addr_4996_7;

Selector_2 s4996_7(wires_1249_6[0], addr_1249_6, addr_positional[19987:19984], addr_4996_7);

wire[31:0] addr_4997_7;

Selector_2 s4997_7(wires_1249_6[1], addr_1249_6, addr_positional[19991:19988], addr_4997_7);

wire[31:0] addr_4998_7;

Selector_2 s4998_7(wires_1249_6[2], addr_1249_6, addr_positional[19995:19992], addr_4998_7);

wire[31:0] addr_4999_7;

Selector_2 s4999_7(wires_1249_6[3], addr_1249_6, addr_positional[19999:19996], addr_4999_7);

wire[31:0] addr_5000_7;

Selector_2 s5000_7(wires_1250_6[0], addr_1250_6, addr_positional[20003:20000], addr_5000_7);

wire[31:0] addr_5001_7;

Selector_2 s5001_7(wires_1250_6[1], addr_1250_6, addr_positional[20007:20004], addr_5001_7);

wire[31:0] addr_5002_7;

Selector_2 s5002_7(wires_1250_6[2], addr_1250_6, addr_positional[20011:20008], addr_5002_7);

wire[31:0] addr_5003_7;

Selector_2 s5003_7(wires_1250_6[3], addr_1250_6, addr_positional[20015:20012], addr_5003_7);

wire[31:0] addr_5004_7;

Selector_2 s5004_7(wires_1251_6[0], addr_1251_6, addr_positional[20019:20016], addr_5004_7);

wire[31:0] addr_5005_7;

Selector_2 s5005_7(wires_1251_6[1], addr_1251_6, addr_positional[20023:20020], addr_5005_7);

wire[31:0] addr_5006_7;

Selector_2 s5006_7(wires_1251_6[2], addr_1251_6, addr_positional[20027:20024], addr_5006_7);

wire[31:0] addr_5007_7;

Selector_2 s5007_7(wires_1251_6[3], addr_1251_6, addr_positional[20031:20028], addr_5007_7);

wire[31:0] addr_5008_7;

Selector_2 s5008_7(wires_1252_6[0], addr_1252_6, addr_positional[20035:20032], addr_5008_7);

wire[31:0] addr_5009_7;

Selector_2 s5009_7(wires_1252_6[1], addr_1252_6, addr_positional[20039:20036], addr_5009_7);

wire[31:0] addr_5010_7;

Selector_2 s5010_7(wires_1252_6[2], addr_1252_6, addr_positional[20043:20040], addr_5010_7);

wire[31:0] addr_5011_7;

Selector_2 s5011_7(wires_1252_6[3], addr_1252_6, addr_positional[20047:20044], addr_5011_7);

wire[31:0] addr_5012_7;

Selector_2 s5012_7(wires_1253_6[0], addr_1253_6, addr_positional[20051:20048], addr_5012_7);

wire[31:0] addr_5013_7;

Selector_2 s5013_7(wires_1253_6[1], addr_1253_6, addr_positional[20055:20052], addr_5013_7);

wire[31:0] addr_5014_7;

Selector_2 s5014_7(wires_1253_6[2], addr_1253_6, addr_positional[20059:20056], addr_5014_7);

wire[31:0] addr_5015_7;

Selector_2 s5015_7(wires_1253_6[3], addr_1253_6, addr_positional[20063:20060], addr_5015_7);

wire[31:0] addr_5016_7;

Selector_2 s5016_7(wires_1254_6[0], addr_1254_6, addr_positional[20067:20064], addr_5016_7);

wire[31:0] addr_5017_7;

Selector_2 s5017_7(wires_1254_6[1], addr_1254_6, addr_positional[20071:20068], addr_5017_7);

wire[31:0] addr_5018_7;

Selector_2 s5018_7(wires_1254_6[2], addr_1254_6, addr_positional[20075:20072], addr_5018_7);

wire[31:0] addr_5019_7;

Selector_2 s5019_7(wires_1254_6[3], addr_1254_6, addr_positional[20079:20076], addr_5019_7);

wire[31:0] addr_5020_7;

Selector_2 s5020_7(wires_1255_6[0], addr_1255_6, addr_positional[20083:20080], addr_5020_7);

wire[31:0] addr_5021_7;

Selector_2 s5021_7(wires_1255_6[1], addr_1255_6, addr_positional[20087:20084], addr_5021_7);

wire[31:0] addr_5022_7;

Selector_2 s5022_7(wires_1255_6[2], addr_1255_6, addr_positional[20091:20088], addr_5022_7);

wire[31:0] addr_5023_7;

Selector_2 s5023_7(wires_1255_6[3], addr_1255_6, addr_positional[20095:20092], addr_5023_7);

wire[31:0] addr_5024_7;

Selector_2 s5024_7(wires_1256_6[0], addr_1256_6, addr_positional[20099:20096], addr_5024_7);

wire[31:0] addr_5025_7;

Selector_2 s5025_7(wires_1256_6[1], addr_1256_6, addr_positional[20103:20100], addr_5025_7);

wire[31:0] addr_5026_7;

Selector_2 s5026_7(wires_1256_6[2], addr_1256_6, addr_positional[20107:20104], addr_5026_7);

wire[31:0] addr_5027_7;

Selector_2 s5027_7(wires_1256_6[3], addr_1256_6, addr_positional[20111:20108], addr_5027_7);

wire[31:0] addr_5028_7;

Selector_2 s5028_7(wires_1257_6[0], addr_1257_6, addr_positional[20115:20112], addr_5028_7);

wire[31:0] addr_5029_7;

Selector_2 s5029_7(wires_1257_6[1], addr_1257_6, addr_positional[20119:20116], addr_5029_7);

wire[31:0] addr_5030_7;

Selector_2 s5030_7(wires_1257_6[2], addr_1257_6, addr_positional[20123:20120], addr_5030_7);

wire[31:0] addr_5031_7;

Selector_2 s5031_7(wires_1257_6[3], addr_1257_6, addr_positional[20127:20124], addr_5031_7);

wire[31:0] addr_5032_7;

Selector_2 s5032_7(wires_1258_6[0], addr_1258_6, addr_positional[20131:20128], addr_5032_7);

wire[31:0] addr_5033_7;

Selector_2 s5033_7(wires_1258_6[1], addr_1258_6, addr_positional[20135:20132], addr_5033_7);

wire[31:0] addr_5034_7;

Selector_2 s5034_7(wires_1258_6[2], addr_1258_6, addr_positional[20139:20136], addr_5034_7);

wire[31:0] addr_5035_7;

Selector_2 s5035_7(wires_1258_6[3], addr_1258_6, addr_positional[20143:20140], addr_5035_7);

wire[31:0] addr_5036_7;

Selector_2 s5036_7(wires_1259_6[0], addr_1259_6, addr_positional[20147:20144], addr_5036_7);

wire[31:0] addr_5037_7;

Selector_2 s5037_7(wires_1259_6[1], addr_1259_6, addr_positional[20151:20148], addr_5037_7);

wire[31:0] addr_5038_7;

Selector_2 s5038_7(wires_1259_6[2], addr_1259_6, addr_positional[20155:20152], addr_5038_7);

wire[31:0] addr_5039_7;

Selector_2 s5039_7(wires_1259_6[3], addr_1259_6, addr_positional[20159:20156], addr_5039_7);

wire[31:0] addr_5040_7;

Selector_2 s5040_7(wires_1260_6[0], addr_1260_6, addr_positional[20163:20160], addr_5040_7);

wire[31:0] addr_5041_7;

Selector_2 s5041_7(wires_1260_6[1], addr_1260_6, addr_positional[20167:20164], addr_5041_7);

wire[31:0] addr_5042_7;

Selector_2 s5042_7(wires_1260_6[2], addr_1260_6, addr_positional[20171:20168], addr_5042_7);

wire[31:0] addr_5043_7;

Selector_2 s5043_7(wires_1260_6[3], addr_1260_6, addr_positional[20175:20172], addr_5043_7);

wire[31:0] addr_5044_7;

Selector_2 s5044_7(wires_1261_6[0], addr_1261_6, addr_positional[20179:20176], addr_5044_7);

wire[31:0] addr_5045_7;

Selector_2 s5045_7(wires_1261_6[1], addr_1261_6, addr_positional[20183:20180], addr_5045_7);

wire[31:0] addr_5046_7;

Selector_2 s5046_7(wires_1261_6[2], addr_1261_6, addr_positional[20187:20184], addr_5046_7);

wire[31:0] addr_5047_7;

Selector_2 s5047_7(wires_1261_6[3], addr_1261_6, addr_positional[20191:20188], addr_5047_7);

wire[31:0] addr_5048_7;

Selector_2 s5048_7(wires_1262_6[0], addr_1262_6, addr_positional[20195:20192], addr_5048_7);

wire[31:0] addr_5049_7;

Selector_2 s5049_7(wires_1262_6[1], addr_1262_6, addr_positional[20199:20196], addr_5049_7);

wire[31:0] addr_5050_7;

Selector_2 s5050_7(wires_1262_6[2], addr_1262_6, addr_positional[20203:20200], addr_5050_7);

wire[31:0] addr_5051_7;

Selector_2 s5051_7(wires_1262_6[3], addr_1262_6, addr_positional[20207:20204], addr_5051_7);

wire[31:0] addr_5052_7;

Selector_2 s5052_7(wires_1263_6[0], addr_1263_6, addr_positional[20211:20208], addr_5052_7);

wire[31:0] addr_5053_7;

Selector_2 s5053_7(wires_1263_6[1], addr_1263_6, addr_positional[20215:20212], addr_5053_7);

wire[31:0] addr_5054_7;

Selector_2 s5054_7(wires_1263_6[2], addr_1263_6, addr_positional[20219:20216], addr_5054_7);

wire[31:0] addr_5055_7;

Selector_2 s5055_7(wires_1263_6[3], addr_1263_6, addr_positional[20223:20220], addr_5055_7);

wire[31:0] addr_5056_7;

Selector_2 s5056_7(wires_1264_6[0], addr_1264_6, addr_positional[20227:20224], addr_5056_7);

wire[31:0] addr_5057_7;

Selector_2 s5057_7(wires_1264_6[1], addr_1264_6, addr_positional[20231:20228], addr_5057_7);

wire[31:0] addr_5058_7;

Selector_2 s5058_7(wires_1264_6[2], addr_1264_6, addr_positional[20235:20232], addr_5058_7);

wire[31:0] addr_5059_7;

Selector_2 s5059_7(wires_1264_6[3], addr_1264_6, addr_positional[20239:20236], addr_5059_7);

wire[31:0] addr_5060_7;

Selector_2 s5060_7(wires_1265_6[0], addr_1265_6, addr_positional[20243:20240], addr_5060_7);

wire[31:0] addr_5061_7;

Selector_2 s5061_7(wires_1265_6[1], addr_1265_6, addr_positional[20247:20244], addr_5061_7);

wire[31:0] addr_5062_7;

Selector_2 s5062_7(wires_1265_6[2], addr_1265_6, addr_positional[20251:20248], addr_5062_7);

wire[31:0] addr_5063_7;

Selector_2 s5063_7(wires_1265_6[3], addr_1265_6, addr_positional[20255:20252], addr_5063_7);

wire[31:0] addr_5064_7;

Selector_2 s5064_7(wires_1266_6[0], addr_1266_6, addr_positional[20259:20256], addr_5064_7);

wire[31:0] addr_5065_7;

Selector_2 s5065_7(wires_1266_6[1], addr_1266_6, addr_positional[20263:20260], addr_5065_7);

wire[31:0] addr_5066_7;

Selector_2 s5066_7(wires_1266_6[2], addr_1266_6, addr_positional[20267:20264], addr_5066_7);

wire[31:0] addr_5067_7;

Selector_2 s5067_7(wires_1266_6[3], addr_1266_6, addr_positional[20271:20268], addr_5067_7);

wire[31:0] addr_5068_7;

Selector_2 s5068_7(wires_1267_6[0], addr_1267_6, addr_positional[20275:20272], addr_5068_7);

wire[31:0] addr_5069_7;

Selector_2 s5069_7(wires_1267_6[1], addr_1267_6, addr_positional[20279:20276], addr_5069_7);

wire[31:0] addr_5070_7;

Selector_2 s5070_7(wires_1267_6[2], addr_1267_6, addr_positional[20283:20280], addr_5070_7);

wire[31:0] addr_5071_7;

Selector_2 s5071_7(wires_1267_6[3], addr_1267_6, addr_positional[20287:20284], addr_5071_7);

wire[31:0] addr_5072_7;

Selector_2 s5072_7(wires_1268_6[0], addr_1268_6, addr_positional[20291:20288], addr_5072_7);

wire[31:0] addr_5073_7;

Selector_2 s5073_7(wires_1268_6[1], addr_1268_6, addr_positional[20295:20292], addr_5073_7);

wire[31:0] addr_5074_7;

Selector_2 s5074_7(wires_1268_6[2], addr_1268_6, addr_positional[20299:20296], addr_5074_7);

wire[31:0] addr_5075_7;

Selector_2 s5075_7(wires_1268_6[3], addr_1268_6, addr_positional[20303:20300], addr_5075_7);

wire[31:0] addr_5076_7;

Selector_2 s5076_7(wires_1269_6[0], addr_1269_6, addr_positional[20307:20304], addr_5076_7);

wire[31:0] addr_5077_7;

Selector_2 s5077_7(wires_1269_6[1], addr_1269_6, addr_positional[20311:20308], addr_5077_7);

wire[31:0] addr_5078_7;

Selector_2 s5078_7(wires_1269_6[2], addr_1269_6, addr_positional[20315:20312], addr_5078_7);

wire[31:0] addr_5079_7;

Selector_2 s5079_7(wires_1269_6[3], addr_1269_6, addr_positional[20319:20316], addr_5079_7);

wire[31:0] addr_5080_7;

Selector_2 s5080_7(wires_1270_6[0], addr_1270_6, addr_positional[20323:20320], addr_5080_7);

wire[31:0] addr_5081_7;

Selector_2 s5081_7(wires_1270_6[1], addr_1270_6, addr_positional[20327:20324], addr_5081_7);

wire[31:0] addr_5082_7;

Selector_2 s5082_7(wires_1270_6[2], addr_1270_6, addr_positional[20331:20328], addr_5082_7);

wire[31:0] addr_5083_7;

Selector_2 s5083_7(wires_1270_6[3], addr_1270_6, addr_positional[20335:20332], addr_5083_7);

wire[31:0] addr_5084_7;

Selector_2 s5084_7(wires_1271_6[0], addr_1271_6, addr_positional[20339:20336], addr_5084_7);

wire[31:0] addr_5085_7;

Selector_2 s5085_7(wires_1271_6[1], addr_1271_6, addr_positional[20343:20340], addr_5085_7);

wire[31:0] addr_5086_7;

Selector_2 s5086_7(wires_1271_6[2], addr_1271_6, addr_positional[20347:20344], addr_5086_7);

wire[31:0] addr_5087_7;

Selector_2 s5087_7(wires_1271_6[3], addr_1271_6, addr_positional[20351:20348], addr_5087_7);

wire[31:0] addr_5088_7;

Selector_2 s5088_7(wires_1272_6[0], addr_1272_6, addr_positional[20355:20352], addr_5088_7);

wire[31:0] addr_5089_7;

Selector_2 s5089_7(wires_1272_6[1], addr_1272_6, addr_positional[20359:20356], addr_5089_7);

wire[31:0] addr_5090_7;

Selector_2 s5090_7(wires_1272_6[2], addr_1272_6, addr_positional[20363:20360], addr_5090_7);

wire[31:0] addr_5091_7;

Selector_2 s5091_7(wires_1272_6[3], addr_1272_6, addr_positional[20367:20364], addr_5091_7);

wire[31:0] addr_5092_7;

Selector_2 s5092_7(wires_1273_6[0], addr_1273_6, addr_positional[20371:20368], addr_5092_7);

wire[31:0] addr_5093_7;

Selector_2 s5093_7(wires_1273_6[1], addr_1273_6, addr_positional[20375:20372], addr_5093_7);

wire[31:0] addr_5094_7;

Selector_2 s5094_7(wires_1273_6[2], addr_1273_6, addr_positional[20379:20376], addr_5094_7);

wire[31:0] addr_5095_7;

Selector_2 s5095_7(wires_1273_6[3], addr_1273_6, addr_positional[20383:20380], addr_5095_7);

wire[31:0] addr_5096_7;

Selector_2 s5096_7(wires_1274_6[0], addr_1274_6, addr_positional[20387:20384], addr_5096_7);

wire[31:0] addr_5097_7;

Selector_2 s5097_7(wires_1274_6[1], addr_1274_6, addr_positional[20391:20388], addr_5097_7);

wire[31:0] addr_5098_7;

Selector_2 s5098_7(wires_1274_6[2], addr_1274_6, addr_positional[20395:20392], addr_5098_7);

wire[31:0] addr_5099_7;

Selector_2 s5099_7(wires_1274_6[3], addr_1274_6, addr_positional[20399:20396], addr_5099_7);

wire[31:0] addr_5100_7;

Selector_2 s5100_7(wires_1275_6[0], addr_1275_6, addr_positional[20403:20400], addr_5100_7);

wire[31:0] addr_5101_7;

Selector_2 s5101_7(wires_1275_6[1], addr_1275_6, addr_positional[20407:20404], addr_5101_7);

wire[31:0] addr_5102_7;

Selector_2 s5102_7(wires_1275_6[2], addr_1275_6, addr_positional[20411:20408], addr_5102_7);

wire[31:0] addr_5103_7;

Selector_2 s5103_7(wires_1275_6[3], addr_1275_6, addr_positional[20415:20412], addr_5103_7);

wire[31:0] addr_5104_7;

Selector_2 s5104_7(wires_1276_6[0], addr_1276_6, addr_positional[20419:20416], addr_5104_7);

wire[31:0] addr_5105_7;

Selector_2 s5105_7(wires_1276_6[1], addr_1276_6, addr_positional[20423:20420], addr_5105_7);

wire[31:0] addr_5106_7;

Selector_2 s5106_7(wires_1276_6[2], addr_1276_6, addr_positional[20427:20424], addr_5106_7);

wire[31:0] addr_5107_7;

Selector_2 s5107_7(wires_1276_6[3], addr_1276_6, addr_positional[20431:20428], addr_5107_7);

wire[31:0] addr_5108_7;

Selector_2 s5108_7(wires_1277_6[0], addr_1277_6, addr_positional[20435:20432], addr_5108_7);

wire[31:0] addr_5109_7;

Selector_2 s5109_7(wires_1277_6[1], addr_1277_6, addr_positional[20439:20436], addr_5109_7);

wire[31:0] addr_5110_7;

Selector_2 s5110_7(wires_1277_6[2], addr_1277_6, addr_positional[20443:20440], addr_5110_7);

wire[31:0] addr_5111_7;

Selector_2 s5111_7(wires_1277_6[3], addr_1277_6, addr_positional[20447:20444], addr_5111_7);

wire[31:0] addr_5112_7;

Selector_2 s5112_7(wires_1278_6[0], addr_1278_6, addr_positional[20451:20448], addr_5112_7);

wire[31:0] addr_5113_7;

Selector_2 s5113_7(wires_1278_6[1], addr_1278_6, addr_positional[20455:20452], addr_5113_7);

wire[31:0] addr_5114_7;

Selector_2 s5114_7(wires_1278_6[2], addr_1278_6, addr_positional[20459:20456], addr_5114_7);

wire[31:0] addr_5115_7;

Selector_2 s5115_7(wires_1278_6[3], addr_1278_6, addr_positional[20463:20460], addr_5115_7);

wire[31:0] addr_5116_7;

Selector_2 s5116_7(wires_1279_6[0], addr_1279_6, addr_positional[20467:20464], addr_5116_7);

wire[31:0] addr_5117_7;

Selector_2 s5117_7(wires_1279_6[1], addr_1279_6, addr_positional[20471:20468], addr_5117_7);

wire[31:0] addr_5118_7;

Selector_2 s5118_7(wires_1279_6[2], addr_1279_6, addr_positional[20475:20472], addr_5118_7);

wire[31:0] addr_5119_7;

Selector_2 s5119_7(wires_1279_6[3], addr_1279_6, addr_positional[20479:20476], addr_5119_7);

wire[31:0] addr_5120_7;

Selector_2 s5120_7(wires_1280_6[0], addr_1280_6, addr_positional[20483:20480], addr_5120_7);

wire[31:0] addr_5121_7;

Selector_2 s5121_7(wires_1280_6[1], addr_1280_6, addr_positional[20487:20484], addr_5121_7);

wire[31:0] addr_5122_7;

Selector_2 s5122_7(wires_1280_6[2], addr_1280_6, addr_positional[20491:20488], addr_5122_7);

wire[31:0] addr_5123_7;

Selector_2 s5123_7(wires_1280_6[3], addr_1280_6, addr_positional[20495:20492], addr_5123_7);

wire[31:0] addr_5124_7;

Selector_2 s5124_7(wires_1281_6[0], addr_1281_6, addr_positional[20499:20496], addr_5124_7);

wire[31:0] addr_5125_7;

Selector_2 s5125_7(wires_1281_6[1], addr_1281_6, addr_positional[20503:20500], addr_5125_7);

wire[31:0] addr_5126_7;

Selector_2 s5126_7(wires_1281_6[2], addr_1281_6, addr_positional[20507:20504], addr_5126_7);

wire[31:0] addr_5127_7;

Selector_2 s5127_7(wires_1281_6[3], addr_1281_6, addr_positional[20511:20508], addr_5127_7);

wire[31:0] addr_5128_7;

Selector_2 s5128_7(wires_1282_6[0], addr_1282_6, addr_positional[20515:20512], addr_5128_7);

wire[31:0] addr_5129_7;

Selector_2 s5129_7(wires_1282_6[1], addr_1282_6, addr_positional[20519:20516], addr_5129_7);

wire[31:0] addr_5130_7;

Selector_2 s5130_7(wires_1282_6[2], addr_1282_6, addr_positional[20523:20520], addr_5130_7);

wire[31:0] addr_5131_7;

Selector_2 s5131_7(wires_1282_6[3], addr_1282_6, addr_positional[20527:20524], addr_5131_7);

wire[31:0] addr_5132_7;

Selector_2 s5132_7(wires_1283_6[0], addr_1283_6, addr_positional[20531:20528], addr_5132_7);

wire[31:0] addr_5133_7;

Selector_2 s5133_7(wires_1283_6[1], addr_1283_6, addr_positional[20535:20532], addr_5133_7);

wire[31:0] addr_5134_7;

Selector_2 s5134_7(wires_1283_6[2], addr_1283_6, addr_positional[20539:20536], addr_5134_7);

wire[31:0] addr_5135_7;

Selector_2 s5135_7(wires_1283_6[3], addr_1283_6, addr_positional[20543:20540], addr_5135_7);

wire[31:0] addr_5136_7;

Selector_2 s5136_7(wires_1284_6[0], addr_1284_6, addr_positional[20547:20544], addr_5136_7);

wire[31:0] addr_5137_7;

Selector_2 s5137_7(wires_1284_6[1], addr_1284_6, addr_positional[20551:20548], addr_5137_7);

wire[31:0] addr_5138_7;

Selector_2 s5138_7(wires_1284_6[2], addr_1284_6, addr_positional[20555:20552], addr_5138_7);

wire[31:0] addr_5139_7;

Selector_2 s5139_7(wires_1284_6[3], addr_1284_6, addr_positional[20559:20556], addr_5139_7);

wire[31:0] addr_5140_7;

Selector_2 s5140_7(wires_1285_6[0], addr_1285_6, addr_positional[20563:20560], addr_5140_7);

wire[31:0] addr_5141_7;

Selector_2 s5141_7(wires_1285_6[1], addr_1285_6, addr_positional[20567:20564], addr_5141_7);

wire[31:0] addr_5142_7;

Selector_2 s5142_7(wires_1285_6[2], addr_1285_6, addr_positional[20571:20568], addr_5142_7);

wire[31:0] addr_5143_7;

Selector_2 s5143_7(wires_1285_6[3], addr_1285_6, addr_positional[20575:20572], addr_5143_7);

wire[31:0] addr_5144_7;

Selector_2 s5144_7(wires_1286_6[0], addr_1286_6, addr_positional[20579:20576], addr_5144_7);

wire[31:0] addr_5145_7;

Selector_2 s5145_7(wires_1286_6[1], addr_1286_6, addr_positional[20583:20580], addr_5145_7);

wire[31:0] addr_5146_7;

Selector_2 s5146_7(wires_1286_6[2], addr_1286_6, addr_positional[20587:20584], addr_5146_7);

wire[31:0] addr_5147_7;

Selector_2 s5147_7(wires_1286_6[3], addr_1286_6, addr_positional[20591:20588], addr_5147_7);

wire[31:0] addr_5148_7;

Selector_2 s5148_7(wires_1287_6[0], addr_1287_6, addr_positional[20595:20592], addr_5148_7);

wire[31:0] addr_5149_7;

Selector_2 s5149_7(wires_1287_6[1], addr_1287_6, addr_positional[20599:20596], addr_5149_7);

wire[31:0] addr_5150_7;

Selector_2 s5150_7(wires_1287_6[2], addr_1287_6, addr_positional[20603:20600], addr_5150_7);

wire[31:0] addr_5151_7;

Selector_2 s5151_7(wires_1287_6[3], addr_1287_6, addr_positional[20607:20604], addr_5151_7);

wire[31:0] addr_5152_7;

Selector_2 s5152_7(wires_1288_6[0], addr_1288_6, addr_positional[20611:20608], addr_5152_7);

wire[31:0] addr_5153_7;

Selector_2 s5153_7(wires_1288_6[1], addr_1288_6, addr_positional[20615:20612], addr_5153_7);

wire[31:0] addr_5154_7;

Selector_2 s5154_7(wires_1288_6[2], addr_1288_6, addr_positional[20619:20616], addr_5154_7);

wire[31:0] addr_5155_7;

Selector_2 s5155_7(wires_1288_6[3], addr_1288_6, addr_positional[20623:20620], addr_5155_7);

wire[31:0] addr_5156_7;

Selector_2 s5156_7(wires_1289_6[0], addr_1289_6, addr_positional[20627:20624], addr_5156_7);

wire[31:0] addr_5157_7;

Selector_2 s5157_7(wires_1289_6[1], addr_1289_6, addr_positional[20631:20628], addr_5157_7);

wire[31:0] addr_5158_7;

Selector_2 s5158_7(wires_1289_6[2], addr_1289_6, addr_positional[20635:20632], addr_5158_7);

wire[31:0] addr_5159_7;

Selector_2 s5159_7(wires_1289_6[3], addr_1289_6, addr_positional[20639:20636], addr_5159_7);

wire[31:0] addr_5160_7;

Selector_2 s5160_7(wires_1290_6[0], addr_1290_6, addr_positional[20643:20640], addr_5160_7);

wire[31:0] addr_5161_7;

Selector_2 s5161_7(wires_1290_6[1], addr_1290_6, addr_positional[20647:20644], addr_5161_7);

wire[31:0] addr_5162_7;

Selector_2 s5162_7(wires_1290_6[2], addr_1290_6, addr_positional[20651:20648], addr_5162_7);

wire[31:0] addr_5163_7;

Selector_2 s5163_7(wires_1290_6[3], addr_1290_6, addr_positional[20655:20652], addr_5163_7);

wire[31:0] addr_5164_7;

Selector_2 s5164_7(wires_1291_6[0], addr_1291_6, addr_positional[20659:20656], addr_5164_7);

wire[31:0] addr_5165_7;

Selector_2 s5165_7(wires_1291_6[1], addr_1291_6, addr_positional[20663:20660], addr_5165_7);

wire[31:0] addr_5166_7;

Selector_2 s5166_7(wires_1291_6[2], addr_1291_6, addr_positional[20667:20664], addr_5166_7);

wire[31:0] addr_5167_7;

Selector_2 s5167_7(wires_1291_6[3], addr_1291_6, addr_positional[20671:20668], addr_5167_7);

wire[31:0] addr_5168_7;

Selector_2 s5168_7(wires_1292_6[0], addr_1292_6, addr_positional[20675:20672], addr_5168_7);

wire[31:0] addr_5169_7;

Selector_2 s5169_7(wires_1292_6[1], addr_1292_6, addr_positional[20679:20676], addr_5169_7);

wire[31:0] addr_5170_7;

Selector_2 s5170_7(wires_1292_6[2], addr_1292_6, addr_positional[20683:20680], addr_5170_7);

wire[31:0] addr_5171_7;

Selector_2 s5171_7(wires_1292_6[3], addr_1292_6, addr_positional[20687:20684], addr_5171_7);

wire[31:0] addr_5172_7;

Selector_2 s5172_7(wires_1293_6[0], addr_1293_6, addr_positional[20691:20688], addr_5172_7);

wire[31:0] addr_5173_7;

Selector_2 s5173_7(wires_1293_6[1], addr_1293_6, addr_positional[20695:20692], addr_5173_7);

wire[31:0] addr_5174_7;

Selector_2 s5174_7(wires_1293_6[2], addr_1293_6, addr_positional[20699:20696], addr_5174_7);

wire[31:0] addr_5175_7;

Selector_2 s5175_7(wires_1293_6[3], addr_1293_6, addr_positional[20703:20700], addr_5175_7);

wire[31:0] addr_5176_7;

Selector_2 s5176_7(wires_1294_6[0], addr_1294_6, addr_positional[20707:20704], addr_5176_7);

wire[31:0] addr_5177_7;

Selector_2 s5177_7(wires_1294_6[1], addr_1294_6, addr_positional[20711:20708], addr_5177_7);

wire[31:0] addr_5178_7;

Selector_2 s5178_7(wires_1294_6[2], addr_1294_6, addr_positional[20715:20712], addr_5178_7);

wire[31:0] addr_5179_7;

Selector_2 s5179_7(wires_1294_6[3], addr_1294_6, addr_positional[20719:20716], addr_5179_7);

wire[31:0] addr_5180_7;

Selector_2 s5180_7(wires_1295_6[0], addr_1295_6, addr_positional[20723:20720], addr_5180_7);

wire[31:0] addr_5181_7;

Selector_2 s5181_7(wires_1295_6[1], addr_1295_6, addr_positional[20727:20724], addr_5181_7);

wire[31:0] addr_5182_7;

Selector_2 s5182_7(wires_1295_6[2], addr_1295_6, addr_positional[20731:20728], addr_5182_7);

wire[31:0] addr_5183_7;

Selector_2 s5183_7(wires_1295_6[3], addr_1295_6, addr_positional[20735:20732], addr_5183_7);

wire[31:0] addr_5184_7;

Selector_2 s5184_7(wires_1296_6[0], addr_1296_6, addr_positional[20739:20736], addr_5184_7);

wire[31:0] addr_5185_7;

Selector_2 s5185_7(wires_1296_6[1], addr_1296_6, addr_positional[20743:20740], addr_5185_7);

wire[31:0] addr_5186_7;

Selector_2 s5186_7(wires_1296_6[2], addr_1296_6, addr_positional[20747:20744], addr_5186_7);

wire[31:0] addr_5187_7;

Selector_2 s5187_7(wires_1296_6[3], addr_1296_6, addr_positional[20751:20748], addr_5187_7);

wire[31:0] addr_5188_7;

Selector_2 s5188_7(wires_1297_6[0], addr_1297_6, addr_positional[20755:20752], addr_5188_7);

wire[31:0] addr_5189_7;

Selector_2 s5189_7(wires_1297_6[1], addr_1297_6, addr_positional[20759:20756], addr_5189_7);

wire[31:0] addr_5190_7;

Selector_2 s5190_7(wires_1297_6[2], addr_1297_6, addr_positional[20763:20760], addr_5190_7);

wire[31:0] addr_5191_7;

Selector_2 s5191_7(wires_1297_6[3], addr_1297_6, addr_positional[20767:20764], addr_5191_7);

wire[31:0] addr_5192_7;

Selector_2 s5192_7(wires_1298_6[0], addr_1298_6, addr_positional[20771:20768], addr_5192_7);

wire[31:0] addr_5193_7;

Selector_2 s5193_7(wires_1298_6[1], addr_1298_6, addr_positional[20775:20772], addr_5193_7);

wire[31:0] addr_5194_7;

Selector_2 s5194_7(wires_1298_6[2], addr_1298_6, addr_positional[20779:20776], addr_5194_7);

wire[31:0] addr_5195_7;

Selector_2 s5195_7(wires_1298_6[3], addr_1298_6, addr_positional[20783:20780], addr_5195_7);

wire[31:0] addr_5196_7;

Selector_2 s5196_7(wires_1299_6[0], addr_1299_6, addr_positional[20787:20784], addr_5196_7);

wire[31:0] addr_5197_7;

Selector_2 s5197_7(wires_1299_6[1], addr_1299_6, addr_positional[20791:20788], addr_5197_7);

wire[31:0] addr_5198_7;

Selector_2 s5198_7(wires_1299_6[2], addr_1299_6, addr_positional[20795:20792], addr_5198_7);

wire[31:0] addr_5199_7;

Selector_2 s5199_7(wires_1299_6[3], addr_1299_6, addr_positional[20799:20796], addr_5199_7);

wire[31:0] addr_5200_7;

Selector_2 s5200_7(wires_1300_6[0], addr_1300_6, addr_positional[20803:20800], addr_5200_7);

wire[31:0] addr_5201_7;

Selector_2 s5201_7(wires_1300_6[1], addr_1300_6, addr_positional[20807:20804], addr_5201_7);

wire[31:0] addr_5202_7;

Selector_2 s5202_7(wires_1300_6[2], addr_1300_6, addr_positional[20811:20808], addr_5202_7);

wire[31:0] addr_5203_7;

Selector_2 s5203_7(wires_1300_6[3], addr_1300_6, addr_positional[20815:20812], addr_5203_7);

wire[31:0] addr_5204_7;

Selector_2 s5204_7(wires_1301_6[0], addr_1301_6, addr_positional[20819:20816], addr_5204_7);

wire[31:0] addr_5205_7;

Selector_2 s5205_7(wires_1301_6[1], addr_1301_6, addr_positional[20823:20820], addr_5205_7);

wire[31:0] addr_5206_7;

Selector_2 s5206_7(wires_1301_6[2], addr_1301_6, addr_positional[20827:20824], addr_5206_7);

wire[31:0] addr_5207_7;

Selector_2 s5207_7(wires_1301_6[3], addr_1301_6, addr_positional[20831:20828], addr_5207_7);

wire[31:0] addr_5208_7;

Selector_2 s5208_7(wires_1302_6[0], addr_1302_6, addr_positional[20835:20832], addr_5208_7);

wire[31:0] addr_5209_7;

Selector_2 s5209_7(wires_1302_6[1], addr_1302_6, addr_positional[20839:20836], addr_5209_7);

wire[31:0] addr_5210_7;

Selector_2 s5210_7(wires_1302_6[2], addr_1302_6, addr_positional[20843:20840], addr_5210_7);

wire[31:0] addr_5211_7;

Selector_2 s5211_7(wires_1302_6[3], addr_1302_6, addr_positional[20847:20844], addr_5211_7);

wire[31:0] addr_5212_7;

Selector_2 s5212_7(wires_1303_6[0], addr_1303_6, addr_positional[20851:20848], addr_5212_7);

wire[31:0] addr_5213_7;

Selector_2 s5213_7(wires_1303_6[1], addr_1303_6, addr_positional[20855:20852], addr_5213_7);

wire[31:0] addr_5214_7;

Selector_2 s5214_7(wires_1303_6[2], addr_1303_6, addr_positional[20859:20856], addr_5214_7);

wire[31:0] addr_5215_7;

Selector_2 s5215_7(wires_1303_6[3], addr_1303_6, addr_positional[20863:20860], addr_5215_7);

wire[31:0] addr_5216_7;

Selector_2 s5216_7(wires_1304_6[0], addr_1304_6, addr_positional[20867:20864], addr_5216_7);

wire[31:0] addr_5217_7;

Selector_2 s5217_7(wires_1304_6[1], addr_1304_6, addr_positional[20871:20868], addr_5217_7);

wire[31:0] addr_5218_7;

Selector_2 s5218_7(wires_1304_6[2], addr_1304_6, addr_positional[20875:20872], addr_5218_7);

wire[31:0] addr_5219_7;

Selector_2 s5219_7(wires_1304_6[3], addr_1304_6, addr_positional[20879:20876], addr_5219_7);

wire[31:0] addr_5220_7;

Selector_2 s5220_7(wires_1305_6[0], addr_1305_6, addr_positional[20883:20880], addr_5220_7);

wire[31:0] addr_5221_7;

Selector_2 s5221_7(wires_1305_6[1], addr_1305_6, addr_positional[20887:20884], addr_5221_7);

wire[31:0] addr_5222_7;

Selector_2 s5222_7(wires_1305_6[2], addr_1305_6, addr_positional[20891:20888], addr_5222_7);

wire[31:0] addr_5223_7;

Selector_2 s5223_7(wires_1305_6[3], addr_1305_6, addr_positional[20895:20892], addr_5223_7);

wire[31:0] addr_5224_7;

Selector_2 s5224_7(wires_1306_6[0], addr_1306_6, addr_positional[20899:20896], addr_5224_7);

wire[31:0] addr_5225_7;

Selector_2 s5225_7(wires_1306_6[1], addr_1306_6, addr_positional[20903:20900], addr_5225_7);

wire[31:0] addr_5226_7;

Selector_2 s5226_7(wires_1306_6[2], addr_1306_6, addr_positional[20907:20904], addr_5226_7);

wire[31:0] addr_5227_7;

Selector_2 s5227_7(wires_1306_6[3], addr_1306_6, addr_positional[20911:20908], addr_5227_7);

wire[31:0] addr_5228_7;

Selector_2 s5228_7(wires_1307_6[0], addr_1307_6, addr_positional[20915:20912], addr_5228_7);

wire[31:0] addr_5229_7;

Selector_2 s5229_7(wires_1307_6[1], addr_1307_6, addr_positional[20919:20916], addr_5229_7);

wire[31:0] addr_5230_7;

Selector_2 s5230_7(wires_1307_6[2], addr_1307_6, addr_positional[20923:20920], addr_5230_7);

wire[31:0] addr_5231_7;

Selector_2 s5231_7(wires_1307_6[3], addr_1307_6, addr_positional[20927:20924], addr_5231_7);

wire[31:0] addr_5232_7;

Selector_2 s5232_7(wires_1308_6[0], addr_1308_6, addr_positional[20931:20928], addr_5232_7);

wire[31:0] addr_5233_7;

Selector_2 s5233_7(wires_1308_6[1], addr_1308_6, addr_positional[20935:20932], addr_5233_7);

wire[31:0] addr_5234_7;

Selector_2 s5234_7(wires_1308_6[2], addr_1308_6, addr_positional[20939:20936], addr_5234_7);

wire[31:0] addr_5235_7;

Selector_2 s5235_7(wires_1308_6[3], addr_1308_6, addr_positional[20943:20940], addr_5235_7);

wire[31:0] addr_5236_7;

Selector_2 s5236_7(wires_1309_6[0], addr_1309_6, addr_positional[20947:20944], addr_5236_7);

wire[31:0] addr_5237_7;

Selector_2 s5237_7(wires_1309_6[1], addr_1309_6, addr_positional[20951:20948], addr_5237_7);

wire[31:0] addr_5238_7;

Selector_2 s5238_7(wires_1309_6[2], addr_1309_6, addr_positional[20955:20952], addr_5238_7);

wire[31:0] addr_5239_7;

Selector_2 s5239_7(wires_1309_6[3], addr_1309_6, addr_positional[20959:20956], addr_5239_7);

wire[31:0] addr_5240_7;

Selector_2 s5240_7(wires_1310_6[0], addr_1310_6, addr_positional[20963:20960], addr_5240_7);

wire[31:0] addr_5241_7;

Selector_2 s5241_7(wires_1310_6[1], addr_1310_6, addr_positional[20967:20964], addr_5241_7);

wire[31:0] addr_5242_7;

Selector_2 s5242_7(wires_1310_6[2], addr_1310_6, addr_positional[20971:20968], addr_5242_7);

wire[31:0] addr_5243_7;

Selector_2 s5243_7(wires_1310_6[3], addr_1310_6, addr_positional[20975:20972], addr_5243_7);

wire[31:0] addr_5244_7;

Selector_2 s5244_7(wires_1311_6[0], addr_1311_6, addr_positional[20979:20976], addr_5244_7);

wire[31:0] addr_5245_7;

Selector_2 s5245_7(wires_1311_6[1], addr_1311_6, addr_positional[20983:20980], addr_5245_7);

wire[31:0] addr_5246_7;

Selector_2 s5246_7(wires_1311_6[2], addr_1311_6, addr_positional[20987:20984], addr_5246_7);

wire[31:0] addr_5247_7;

Selector_2 s5247_7(wires_1311_6[3], addr_1311_6, addr_positional[20991:20988], addr_5247_7);

wire[31:0] addr_5248_7;

Selector_2 s5248_7(wires_1312_6[0], addr_1312_6, addr_positional[20995:20992], addr_5248_7);

wire[31:0] addr_5249_7;

Selector_2 s5249_7(wires_1312_6[1], addr_1312_6, addr_positional[20999:20996], addr_5249_7);

wire[31:0] addr_5250_7;

Selector_2 s5250_7(wires_1312_6[2], addr_1312_6, addr_positional[21003:21000], addr_5250_7);

wire[31:0] addr_5251_7;

Selector_2 s5251_7(wires_1312_6[3], addr_1312_6, addr_positional[21007:21004], addr_5251_7);

wire[31:0] addr_5252_7;

Selector_2 s5252_7(wires_1313_6[0], addr_1313_6, addr_positional[21011:21008], addr_5252_7);

wire[31:0] addr_5253_7;

Selector_2 s5253_7(wires_1313_6[1], addr_1313_6, addr_positional[21015:21012], addr_5253_7);

wire[31:0] addr_5254_7;

Selector_2 s5254_7(wires_1313_6[2], addr_1313_6, addr_positional[21019:21016], addr_5254_7);

wire[31:0] addr_5255_7;

Selector_2 s5255_7(wires_1313_6[3], addr_1313_6, addr_positional[21023:21020], addr_5255_7);

wire[31:0] addr_5256_7;

Selector_2 s5256_7(wires_1314_6[0], addr_1314_6, addr_positional[21027:21024], addr_5256_7);

wire[31:0] addr_5257_7;

Selector_2 s5257_7(wires_1314_6[1], addr_1314_6, addr_positional[21031:21028], addr_5257_7);

wire[31:0] addr_5258_7;

Selector_2 s5258_7(wires_1314_6[2], addr_1314_6, addr_positional[21035:21032], addr_5258_7);

wire[31:0] addr_5259_7;

Selector_2 s5259_7(wires_1314_6[3], addr_1314_6, addr_positional[21039:21036], addr_5259_7);

wire[31:0] addr_5260_7;

Selector_2 s5260_7(wires_1315_6[0], addr_1315_6, addr_positional[21043:21040], addr_5260_7);

wire[31:0] addr_5261_7;

Selector_2 s5261_7(wires_1315_6[1], addr_1315_6, addr_positional[21047:21044], addr_5261_7);

wire[31:0] addr_5262_7;

Selector_2 s5262_7(wires_1315_6[2], addr_1315_6, addr_positional[21051:21048], addr_5262_7);

wire[31:0] addr_5263_7;

Selector_2 s5263_7(wires_1315_6[3], addr_1315_6, addr_positional[21055:21052], addr_5263_7);

wire[31:0] addr_5264_7;

Selector_2 s5264_7(wires_1316_6[0], addr_1316_6, addr_positional[21059:21056], addr_5264_7);

wire[31:0] addr_5265_7;

Selector_2 s5265_7(wires_1316_6[1], addr_1316_6, addr_positional[21063:21060], addr_5265_7);

wire[31:0] addr_5266_7;

Selector_2 s5266_7(wires_1316_6[2], addr_1316_6, addr_positional[21067:21064], addr_5266_7);

wire[31:0] addr_5267_7;

Selector_2 s5267_7(wires_1316_6[3], addr_1316_6, addr_positional[21071:21068], addr_5267_7);

wire[31:0] addr_5268_7;

Selector_2 s5268_7(wires_1317_6[0], addr_1317_6, addr_positional[21075:21072], addr_5268_7);

wire[31:0] addr_5269_7;

Selector_2 s5269_7(wires_1317_6[1], addr_1317_6, addr_positional[21079:21076], addr_5269_7);

wire[31:0] addr_5270_7;

Selector_2 s5270_7(wires_1317_6[2], addr_1317_6, addr_positional[21083:21080], addr_5270_7);

wire[31:0] addr_5271_7;

Selector_2 s5271_7(wires_1317_6[3], addr_1317_6, addr_positional[21087:21084], addr_5271_7);

wire[31:0] addr_5272_7;

Selector_2 s5272_7(wires_1318_6[0], addr_1318_6, addr_positional[21091:21088], addr_5272_7);

wire[31:0] addr_5273_7;

Selector_2 s5273_7(wires_1318_6[1], addr_1318_6, addr_positional[21095:21092], addr_5273_7);

wire[31:0] addr_5274_7;

Selector_2 s5274_7(wires_1318_6[2], addr_1318_6, addr_positional[21099:21096], addr_5274_7);

wire[31:0] addr_5275_7;

Selector_2 s5275_7(wires_1318_6[3], addr_1318_6, addr_positional[21103:21100], addr_5275_7);

wire[31:0] addr_5276_7;

Selector_2 s5276_7(wires_1319_6[0], addr_1319_6, addr_positional[21107:21104], addr_5276_7);

wire[31:0] addr_5277_7;

Selector_2 s5277_7(wires_1319_6[1], addr_1319_6, addr_positional[21111:21108], addr_5277_7);

wire[31:0] addr_5278_7;

Selector_2 s5278_7(wires_1319_6[2], addr_1319_6, addr_positional[21115:21112], addr_5278_7);

wire[31:0] addr_5279_7;

Selector_2 s5279_7(wires_1319_6[3], addr_1319_6, addr_positional[21119:21116], addr_5279_7);

wire[31:0] addr_5280_7;

Selector_2 s5280_7(wires_1320_6[0], addr_1320_6, addr_positional[21123:21120], addr_5280_7);

wire[31:0] addr_5281_7;

Selector_2 s5281_7(wires_1320_6[1], addr_1320_6, addr_positional[21127:21124], addr_5281_7);

wire[31:0] addr_5282_7;

Selector_2 s5282_7(wires_1320_6[2], addr_1320_6, addr_positional[21131:21128], addr_5282_7);

wire[31:0] addr_5283_7;

Selector_2 s5283_7(wires_1320_6[3], addr_1320_6, addr_positional[21135:21132], addr_5283_7);

wire[31:0] addr_5284_7;

Selector_2 s5284_7(wires_1321_6[0], addr_1321_6, addr_positional[21139:21136], addr_5284_7);

wire[31:0] addr_5285_7;

Selector_2 s5285_7(wires_1321_6[1], addr_1321_6, addr_positional[21143:21140], addr_5285_7);

wire[31:0] addr_5286_7;

Selector_2 s5286_7(wires_1321_6[2], addr_1321_6, addr_positional[21147:21144], addr_5286_7);

wire[31:0] addr_5287_7;

Selector_2 s5287_7(wires_1321_6[3], addr_1321_6, addr_positional[21151:21148], addr_5287_7);

wire[31:0] addr_5288_7;

Selector_2 s5288_7(wires_1322_6[0], addr_1322_6, addr_positional[21155:21152], addr_5288_7);

wire[31:0] addr_5289_7;

Selector_2 s5289_7(wires_1322_6[1], addr_1322_6, addr_positional[21159:21156], addr_5289_7);

wire[31:0] addr_5290_7;

Selector_2 s5290_7(wires_1322_6[2], addr_1322_6, addr_positional[21163:21160], addr_5290_7);

wire[31:0] addr_5291_7;

Selector_2 s5291_7(wires_1322_6[3], addr_1322_6, addr_positional[21167:21164], addr_5291_7);

wire[31:0] addr_5292_7;

Selector_2 s5292_7(wires_1323_6[0], addr_1323_6, addr_positional[21171:21168], addr_5292_7);

wire[31:0] addr_5293_7;

Selector_2 s5293_7(wires_1323_6[1], addr_1323_6, addr_positional[21175:21172], addr_5293_7);

wire[31:0] addr_5294_7;

Selector_2 s5294_7(wires_1323_6[2], addr_1323_6, addr_positional[21179:21176], addr_5294_7);

wire[31:0] addr_5295_7;

Selector_2 s5295_7(wires_1323_6[3], addr_1323_6, addr_positional[21183:21180], addr_5295_7);

wire[31:0] addr_5296_7;

Selector_2 s5296_7(wires_1324_6[0], addr_1324_6, addr_positional[21187:21184], addr_5296_7);

wire[31:0] addr_5297_7;

Selector_2 s5297_7(wires_1324_6[1], addr_1324_6, addr_positional[21191:21188], addr_5297_7);

wire[31:0] addr_5298_7;

Selector_2 s5298_7(wires_1324_6[2], addr_1324_6, addr_positional[21195:21192], addr_5298_7);

wire[31:0] addr_5299_7;

Selector_2 s5299_7(wires_1324_6[3], addr_1324_6, addr_positional[21199:21196], addr_5299_7);

wire[31:0] addr_5300_7;

Selector_2 s5300_7(wires_1325_6[0], addr_1325_6, addr_positional[21203:21200], addr_5300_7);

wire[31:0] addr_5301_7;

Selector_2 s5301_7(wires_1325_6[1], addr_1325_6, addr_positional[21207:21204], addr_5301_7);

wire[31:0] addr_5302_7;

Selector_2 s5302_7(wires_1325_6[2], addr_1325_6, addr_positional[21211:21208], addr_5302_7);

wire[31:0] addr_5303_7;

Selector_2 s5303_7(wires_1325_6[3], addr_1325_6, addr_positional[21215:21212], addr_5303_7);

wire[31:0] addr_5304_7;

Selector_2 s5304_7(wires_1326_6[0], addr_1326_6, addr_positional[21219:21216], addr_5304_7);

wire[31:0] addr_5305_7;

Selector_2 s5305_7(wires_1326_6[1], addr_1326_6, addr_positional[21223:21220], addr_5305_7);

wire[31:0] addr_5306_7;

Selector_2 s5306_7(wires_1326_6[2], addr_1326_6, addr_positional[21227:21224], addr_5306_7);

wire[31:0] addr_5307_7;

Selector_2 s5307_7(wires_1326_6[3], addr_1326_6, addr_positional[21231:21228], addr_5307_7);

wire[31:0] addr_5308_7;

Selector_2 s5308_7(wires_1327_6[0], addr_1327_6, addr_positional[21235:21232], addr_5308_7);

wire[31:0] addr_5309_7;

Selector_2 s5309_7(wires_1327_6[1], addr_1327_6, addr_positional[21239:21236], addr_5309_7);

wire[31:0] addr_5310_7;

Selector_2 s5310_7(wires_1327_6[2], addr_1327_6, addr_positional[21243:21240], addr_5310_7);

wire[31:0] addr_5311_7;

Selector_2 s5311_7(wires_1327_6[3], addr_1327_6, addr_positional[21247:21244], addr_5311_7);

wire[31:0] addr_5312_7;

Selector_2 s5312_7(wires_1328_6[0], addr_1328_6, addr_positional[21251:21248], addr_5312_7);

wire[31:0] addr_5313_7;

Selector_2 s5313_7(wires_1328_6[1], addr_1328_6, addr_positional[21255:21252], addr_5313_7);

wire[31:0] addr_5314_7;

Selector_2 s5314_7(wires_1328_6[2], addr_1328_6, addr_positional[21259:21256], addr_5314_7);

wire[31:0] addr_5315_7;

Selector_2 s5315_7(wires_1328_6[3], addr_1328_6, addr_positional[21263:21260], addr_5315_7);

wire[31:0] addr_5316_7;

Selector_2 s5316_7(wires_1329_6[0], addr_1329_6, addr_positional[21267:21264], addr_5316_7);

wire[31:0] addr_5317_7;

Selector_2 s5317_7(wires_1329_6[1], addr_1329_6, addr_positional[21271:21268], addr_5317_7);

wire[31:0] addr_5318_7;

Selector_2 s5318_7(wires_1329_6[2], addr_1329_6, addr_positional[21275:21272], addr_5318_7);

wire[31:0] addr_5319_7;

Selector_2 s5319_7(wires_1329_6[3], addr_1329_6, addr_positional[21279:21276], addr_5319_7);

wire[31:0] addr_5320_7;

Selector_2 s5320_7(wires_1330_6[0], addr_1330_6, addr_positional[21283:21280], addr_5320_7);

wire[31:0] addr_5321_7;

Selector_2 s5321_7(wires_1330_6[1], addr_1330_6, addr_positional[21287:21284], addr_5321_7);

wire[31:0] addr_5322_7;

Selector_2 s5322_7(wires_1330_6[2], addr_1330_6, addr_positional[21291:21288], addr_5322_7);

wire[31:0] addr_5323_7;

Selector_2 s5323_7(wires_1330_6[3], addr_1330_6, addr_positional[21295:21292], addr_5323_7);

wire[31:0] addr_5324_7;

Selector_2 s5324_7(wires_1331_6[0], addr_1331_6, addr_positional[21299:21296], addr_5324_7);

wire[31:0] addr_5325_7;

Selector_2 s5325_7(wires_1331_6[1], addr_1331_6, addr_positional[21303:21300], addr_5325_7);

wire[31:0] addr_5326_7;

Selector_2 s5326_7(wires_1331_6[2], addr_1331_6, addr_positional[21307:21304], addr_5326_7);

wire[31:0] addr_5327_7;

Selector_2 s5327_7(wires_1331_6[3], addr_1331_6, addr_positional[21311:21308], addr_5327_7);

wire[31:0] addr_5328_7;

Selector_2 s5328_7(wires_1332_6[0], addr_1332_6, addr_positional[21315:21312], addr_5328_7);

wire[31:0] addr_5329_7;

Selector_2 s5329_7(wires_1332_6[1], addr_1332_6, addr_positional[21319:21316], addr_5329_7);

wire[31:0] addr_5330_7;

Selector_2 s5330_7(wires_1332_6[2], addr_1332_6, addr_positional[21323:21320], addr_5330_7);

wire[31:0] addr_5331_7;

Selector_2 s5331_7(wires_1332_6[3], addr_1332_6, addr_positional[21327:21324], addr_5331_7);

wire[31:0] addr_5332_7;

Selector_2 s5332_7(wires_1333_6[0], addr_1333_6, addr_positional[21331:21328], addr_5332_7);

wire[31:0] addr_5333_7;

Selector_2 s5333_7(wires_1333_6[1], addr_1333_6, addr_positional[21335:21332], addr_5333_7);

wire[31:0] addr_5334_7;

Selector_2 s5334_7(wires_1333_6[2], addr_1333_6, addr_positional[21339:21336], addr_5334_7);

wire[31:0] addr_5335_7;

Selector_2 s5335_7(wires_1333_6[3], addr_1333_6, addr_positional[21343:21340], addr_5335_7);

wire[31:0] addr_5336_7;

Selector_2 s5336_7(wires_1334_6[0], addr_1334_6, addr_positional[21347:21344], addr_5336_7);

wire[31:0] addr_5337_7;

Selector_2 s5337_7(wires_1334_6[1], addr_1334_6, addr_positional[21351:21348], addr_5337_7);

wire[31:0] addr_5338_7;

Selector_2 s5338_7(wires_1334_6[2], addr_1334_6, addr_positional[21355:21352], addr_5338_7);

wire[31:0] addr_5339_7;

Selector_2 s5339_7(wires_1334_6[3], addr_1334_6, addr_positional[21359:21356], addr_5339_7);

wire[31:0] addr_5340_7;

Selector_2 s5340_7(wires_1335_6[0], addr_1335_6, addr_positional[21363:21360], addr_5340_7);

wire[31:0] addr_5341_7;

Selector_2 s5341_7(wires_1335_6[1], addr_1335_6, addr_positional[21367:21364], addr_5341_7);

wire[31:0] addr_5342_7;

Selector_2 s5342_7(wires_1335_6[2], addr_1335_6, addr_positional[21371:21368], addr_5342_7);

wire[31:0] addr_5343_7;

Selector_2 s5343_7(wires_1335_6[3], addr_1335_6, addr_positional[21375:21372], addr_5343_7);

wire[31:0] addr_5344_7;

Selector_2 s5344_7(wires_1336_6[0], addr_1336_6, addr_positional[21379:21376], addr_5344_7);

wire[31:0] addr_5345_7;

Selector_2 s5345_7(wires_1336_6[1], addr_1336_6, addr_positional[21383:21380], addr_5345_7);

wire[31:0] addr_5346_7;

Selector_2 s5346_7(wires_1336_6[2], addr_1336_6, addr_positional[21387:21384], addr_5346_7);

wire[31:0] addr_5347_7;

Selector_2 s5347_7(wires_1336_6[3], addr_1336_6, addr_positional[21391:21388], addr_5347_7);

wire[31:0] addr_5348_7;

Selector_2 s5348_7(wires_1337_6[0], addr_1337_6, addr_positional[21395:21392], addr_5348_7);

wire[31:0] addr_5349_7;

Selector_2 s5349_7(wires_1337_6[1], addr_1337_6, addr_positional[21399:21396], addr_5349_7);

wire[31:0] addr_5350_7;

Selector_2 s5350_7(wires_1337_6[2], addr_1337_6, addr_positional[21403:21400], addr_5350_7);

wire[31:0] addr_5351_7;

Selector_2 s5351_7(wires_1337_6[3], addr_1337_6, addr_positional[21407:21404], addr_5351_7);

wire[31:0] addr_5352_7;

Selector_2 s5352_7(wires_1338_6[0], addr_1338_6, addr_positional[21411:21408], addr_5352_7);

wire[31:0] addr_5353_7;

Selector_2 s5353_7(wires_1338_6[1], addr_1338_6, addr_positional[21415:21412], addr_5353_7);

wire[31:0] addr_5354_7;

Selector_2 s5354_7(wires_1338_6[2], addr_1338_6, addr_positional[21419:21416], addr_5354_7);

wire[31:0] addr_5355_7;

Selector_2 s5355_7(wires_1338_6[3], addr_1338_6, addr_positional[21423:21420], addr_5355_7);

wire[31:0] addr_5356_7;

Selector_2 s5356_7(wires_1339_6[0], addr_1339_6, addr_positional[21427:21424], addr_5356_7);

wire[31:0] addr_5357_7;

Selector_2 s5357_7(wires_1339_6[1], addr_1339_6, addr_positional[21431:21428], addr_5357_7);

wire[31:0] addr_5358_7;

Selector_2 s5358_7(wires_1339_6[2], addr_1339_6, addr_positional[21435:21432], addr_5358_7);

wire[31:0] addr_5359_7;

Selector_2 s5359_7(wires_1339_6[3], addr_1339_6, addr_positional[21439:21436], addr_5359_7);

wire[31:0] addr_5360_7;

Selector_2 s5360_7(wires_1340_6[0], addr_1340_6, addr_positional[21443:21440], addr_5360_7);

wire[31:0] addr_5361_7;

Selector_2 s5361_7(wires_1340_6[1], addr_1340_6, addr_positional[21447:21444], addr_5361_7);

wire[31:0] addr_5362_7;

Selector_2 s5362_7(wires_1340_6[2], addr_1340_6, addr_positional[21451:21448], addr_5362_7);

wire[31:0] addr_5363_7;

Selector_2 s5363_7(wires_1340_6[3], addr_1340_6, addr_positional[21455:21452], addr_5363_7);

wire[31:0] addr_5364_7;

Selector_2 s5364_7(wires_1341_6[0], addr_1341_6, addr_positional[21459:21456], addr_5364_7);

wire[31:0] addr_5365_7;

Selector_2 s5365_7(wires_1341_6[1], addr_1341_6, addr_positional[21463:21460], addr_5365_7);

wire[31:0] addr_5366_7;

Selector_2 s5366_7(wires_1341_6[2], addr_1341_6, addr_positional[21467:21464], addr_5366_7);

wire[31:0] addr_5367_7;

Selector_2 s5367_7(wires_1341_6[3], addr_1341_6, addr_positional[21471:21468], addr_5367_7);

wire[31:0] addr_5368_7;

Selector_2 s5368_7(wires_1342_6[0], addr_1342_6, addr_positional[21475:21472], addr_5368_7);

wire[31:0] addr_5369_7;

Selector_2 s5369_7(wires_1342_6[1], addr_1342_6, addr_positional[21479:21476], addr_5369_7);

wire[31:0] addr_5370_7;

Selector_2 s5370_7(wires_1342_6[2], addr_1342_6, addr_positional[21483:21480], addr_5370_7);

wire[31:0] addr_5371_7;

Selector_2 s5371_7(wires_1342_6[3], addr_1342_6, addr_positional[21487:21484], addr_5371_7);

wire[31:0] addr_5372_7;

Selector_2 s5372_7(wires_1343_6[0], addr_1343_6, addr_positional[21491:21488], addr_5372_7);

wire[31:0] addr_5373_7;

Selector_2 s5373_7(wires_1343_6[1], addr_1343_6, addr_positional[21495:21492], addr_5373_7);

wire[31:0] addr_5374_7;

Selector_2 s5374_7(wires_1343_6[2], addr_1343_6, addr_positional[21499:21496], addr_5374_7);

wire[31:0] addr_5375_7;

Selector_2 s5375_7(wires_1343_6[3], addr_1343_6, addr_positional[21503:21500], addr_5375_7);

wire[31:0] addr_5376_7;

Selector_2 s5376_7(wires_1344_6[0], addr_1344_6, addr_positional[21507:21504], addr_5376_7);

wire[31:0] addr_5377_7;

Selector_2 s5377_7(wires_1344_6[1], addr_1344_6, addr_positional[21511:21508], addr_5377_7);

wire[31:0] addr_5378_7;

Selector_2 s5378_7(wires_1344_6[2], addr_1344_6, addr_positional[21515:21512], addr_5378_7);

wire[31:0] addr_5379_7;

Selector_2 s5379_7(wires_1344_6[3], addr_1344_6, addr_positional[21519:21516], addr_5379_7);

wire[31:0] addr_5380_7;

Selector_2 s5380_7(wires_1345_6[0], addr_1345_6, addr_positional[21523:21520], addr_5380_7);

wire[31:0] addr_5381_7;

Selector_2 s5381_7(wires_1345_6[1], addr_1345_6, addr_positional[21527:21524], addr_5381_7);

wire[31:0] addr_5382_7;

Selector_2 s5382_7(wires_1345_6[2], addr_1345_6, addr_positional[21531:21528], addr_5382_7);

wire[31:0] addr_5383_7;

Selector_2 s5383_7(wires_1345_6[3], addr_1345_6, addr_positional[21535:21532], addr_5383_7);

wire[31:0] addr_5384_7;

Selector_2 s5384_7(wires_1346_6[0], addr_1346_6, addr_positional[21539:21536], addr_5384_7);

wire[31:0] addr_5385_7;

Selector_2 s5385_7(wires_1346_6[1], addr_1346_6, addr_positional[21543:21540], addr_5385_7);

wire[31:0] addr_5386_7;

Selector_2 s5386_7(wires_1346_6[2], addr_1346_6, addr_positional[21547:21544], addr_5386_7);

wire[31:0] addr_5387_7;

Selector_2 s5387_7(wires_1346_6[3], addr_1346_6, addr_positional[21551:21548], addr_5387_7);

wire[31:0] addr_5388_7;

Selector_2 s5388_7(wires_1347_6[0], addr_1347_6, addr_positional[21555:21552], addr_5388_7);

wire[31:0] addr_5389_7;

Selector_2 s5389_7(wires_1347_6[1], addr_1347_6, addr_positional[21559:21556], addr_5389_7);

wire[31:0] addr_5390_7;

Selector_2 s5390_7(wires_1347_6[2], addr_1347_6, addr_positional[21563:21560], addr_5390_7);

wire[31:0] addr_5391_7;

Selector_2 s5391_7(wires_1347_6[3], addr_1347_6, addr_positional[21567:21564], addr_5391_7);

wire[31:0] addr_5392_7;

Selector_2 s5392_7(wires_1348_6[0], addr_1348_6, addr_positional[21571:21568], addr_5392_7);

wire[31:0] addr_5393_7;

Selector_2 s5393_7(wires_1348_6[1], addr_1348_6, addr_positional[21575:21572], addr_5393_7);

wire[31:0] addr_5394_7;

Selector_2 s5394_7(wires_1348_6[2], addr_1348_6, addr_positional[21579:21576], addr_5394_7);

wire[31:0] addr_5395_7;

Selector_2 s5395_7(wires_1348_6[3], addr_1348_6, addr_positional[21583:21580], addr_5395_7);

wire[31:0] addr_5396_7;

Selector_2 s5396_7(wires_1349_6[0], addr_1349_6, addr_positional[21587:21584], addr_5396_7);

wire[31:0] addr_5397_7;

Selector_2 s5397_7(wires_1349_6[1], addr_1349_6, addr_positional[21591:21588], addr_5397_7);

wire[31:0] addr_5398_7;

Selector_2 s5398_7(wires_1349_6[2], addr_1349_6, addr_positional[21595:21592], addr_5398_7);

wire[31:0] addr_5399_7;

Selector_2 s5399_7(wires_1349_6[3], addr_1349_6, addr_positional[21599:21596], addr_5399_7);

wire[31:0] addr_5400_7;

Selector_2 s5400_7(wires_1350_6[0], addr_1350_6, addr_positional[21603:21600], addr_5400_7);

wire[31:0] addr_5401_7;

Selector_2 s5401_7(wires_1350_6[1], addr_1350_6, addr_positional[21607:21604], addr_5401_7);

wire[31:0] addr_5402_7;

Selector_2 s5402_7(wires_1350_6[2], addr_1350_6, addr_positional[21611:21608], addr_5402_7);

wire[31:0] addr_5403_7;

Selector_2 s5403_7(wires_1350_6[3], addr_1350_6, addr_positional[21615:21612], addr_5403_7);

wire[31:0] addr_5404_7;

Selector_2 s5404_7(wires_1351_6[0], addr_1351_6, addr_positional[21619:21616], addr_5404_7);

wire[31:0] addr_5405_7;

Selector_2 s5405_7(wires_1351_6[1], addr_1351_6, addr_positional[21623:21620], addr_5405_7);

wire[31:0] addr_5406_7;

Selector_2 s5406_7(wires_1351_6[2], addr_1351_6, addr_positional[21627:21624], addr_5406_7);

wire[31:0] addr_5407_7;

Selector_2 s5407_7(wires_1351_6[3], addr_1351_6, addr_positional[21631:21628], addr_5407_7);

wire[31:0] addr_5408_7;

Selector_2 s5408_7(wires_1352_6[0], addr_1352_6, addr_positional[21635:21632], addr_5408_7);

wire[31:0] addr_5409_7;

Selector_2 s5409_7(wires_1352_6[1], addr_1352_6, addr_positional[21639:21636], addr_5409_7);

wire[31:0] addr_5410_7;

Selector_2 s5410_7(wires_1352_6[2], addr_1352_6, addr_positional[21643:21640], addr_5410_7);

wire[31:0] addr_5411_7;

Selector_2 s5411_7(wires_1352_6[3], addr_1352_6, addr_positional[21647:21644], addr_5411_7);

wire[31:0] addr_5412_7;

Selector_2 s5412_7(wires_1353_6[0], addr_1353_6, addr_positional[21651:21648], addr_5412_7);

wire[31:0] addr_5413_7;

Selector_2 s5413_7(wires_1353_6[1], addr_1353_6, addr_positional[21655:21652], addr_5413_7);

wire[31:0] addr_5414_7;

Selector_2 s5414_7(wires_1353_6[2], addr_1353_6, addr_positional[21659:21656], addr_5414_7);

wire[31:0] addr_5415_7;

Selector_2 s5415_7(wires_1353_6[3], addr_1353_6, addr_positional[21663:21660], addr_5415_7);

wire[31:0] addr_5416_7;

Selector_2 s5416_7(wires_1354_6[0], addr_1354_6, addr_positional[21667:21664], addr_5416_7);

wire[31:0] addr_5417_7;

Selector_2 s5417_7(wires_1354_6[1], addr_1354_6, addr_positional[21671:21668], addr_5417_7);

wire[31:0] addr_5418_7;

Selector_2 s5418_7(wires_1354_6[2], addr_1354_6, addr_positional[21675:21672], addr_5418_7);

wire[31:0] addr_5419_7;

Selector_2 s5419_7(wires_1354_6[3], addr_1354_6, addr_positional[21679:21676], addr_5419_7);

wire[31:0] addr_5420_7;

Selector_2 s5420_7(wires_1355_6[0], addr_1355_6, addr_positional[21683:21680], addr_5420_7);

wire[31:0] addr_5421_7;

Selector_2 s5421_7(wires_1355_6[1], addr_1355_6, addr_positional[21687:21684], addr_5421_7);

wire[31:0] addr_5422_7;

Selector_2 s5422_7(wires_1355_6[2], addr_1355_6, addr_positional[21691:21688], addr_5422_7);

wire[31:0] addr_5423_7;

Selector_2 s5423_7(wires_1355_6[3], addr_1355_6, addr_positional[21695:21692], addr_5423_7);

wire[31:0] addr_5424_7;

Selector_2 s5424_7(wires_1356_6[0], addr_1356_6, addr_positional[21699:21696], addr_5424_7);

wire[31:0] addr_5425_7;

Selector_2 s5425_7(wires_1356_6[1], addr_1356_6, addr_positional[21703:21700], addr_5425_7);

wire[31:0] addr_5426_7;

Selector_2 s5426_7(wires_1356_6[2], addr_1356_6, addr_positional[21707:21704], addr_5426_7);

wire[31:0] addr_5427_7;

Selector_2 s5427_7(wires_1356_6[3], addr_1356_6, addr_positional[21711:21708], addr_5427_7);

wire[31:0] addr_5428_7;

Selector_2 s5428_7(wires_1357_6[0], addr_1357_6, addr_positional[21715:21712], addr_5428_7);

wire[31:0] addr_5429_7;

Selector_2 s5429_7(wires_1357_6[1], addr_1357_6, addr_positional[21719:21716], addr_5429_7);

wire[31:0] addr_5430_7;

Selector_2 s5430_7(wires_1357_6[2], addr_1357_6, addr_positional[21723:21720], addr_5430_7);

wire[31:0] addr_5431_7;

Selector_2 s5431_7(wires_1357_6[3], addr_1357_6, addr_positional[21727:21724], addr_5431_7);

wire[31:0] addr_5432_7;

Selector_2 s5432_7(wires_1358_6[0], addr_1358_6, addr_positional[21731:21728], addr_5432_7);

wire[31:0] addr_5433_7;

Selector_2 s5433_7(wires_1358_6[1], addr_1358_6, addr_positional[21735:21732], addr_5433_7);

wire[31:0] addr_5434_7;

Selector_2 s5434_7(wires_1358_6[2], addr_1358_6, addr_positional[21739:21736], addr_5434_7);

wire[31:0] addr_5435_7;

Selector_2 s5435_7(wires_1358_6[3], addr_1358_6, addr_positional[21743:21740], addr_5435_7);

wire[31:0] addr_5436_7;

Selector_2 s5436_7(wires_1359_6[0], addr_1359_6, addr_positional[21747:21744], addr_5436_7);

wire[31:0] addr_5437_7;

Selector_2 s5437_7(wires_1359_6[1], addr_1359_6, addr_positional[21751:21748], addr_5437_7);

wire[31:0] addr_5438_7;

Selector_2 s5438_7(wires_1359_6[2], addr_1359_6, addr_positional[21755:21752], addr_5438_7);

wire[31:0] addr_5439_7;

Selector_2 s5439_7(wires_1359_6[3], addr_1359_6, addr_positional[21759:21756], addr_5439_7);

wire[31:0] addr_5440_7;

Selector_2 s5440_7(wires_1360_6[0], addr_1360_6, addr_positional[21763:21760], addr_5440_7);

wire[31:0] addr_5441_7;

Selector_2 s5441_7(wires_1360_6[1], addr_1360_6, addr_positional[21767:21764], addr_5441_7);

wire[31:0] addr_5442_7;

Selector_2 s5442_7(wires_1360_6[2], addr_1360_6, addr_positional[21771:21768], addr_5442_7);

wire[31:0] addr_5443_7;

Selector_2 s5443_7(wires_1360_6[3], addr_1360_6, addr_positional[21775:21772], addr_5443_7);

wire[31:0] addr_5444_7;

Selector_2 s5444_7(wires_1361_6[0], addr_1361_6, addr_positional[21779:21776], addr_5444_7);

wire[31:0] addr_5445_7;

Selector_2 s5445_7(wires_1361_6[1], addr_1361_6, addr_positional[21783:21780], addr_5445_7);

wire[31:0] addr_5446_7;

Selector_2 s5446_7(wires_1361_6[2], addr_1361_6, addr_positional[21787:21784], addr_5446_7);

wire[31:0] addr_5447_7;

Selector_2 s5447_7(wires_1361_6[3], addr_1361_6, addr_positional[21791:21788], addr_5447_7);

wire[31:0] addr_5448_7;

Selector_2 s5448_7(wires_1362_6[0], addr_1362_6, addr_positional[21795:21792], addr_5448_7);

wire[31:0] addr_5449_7;

Selector_2 s5449_7(wires_1362_6[1], addr_1362_6, addr_positional[21799:21796], addr_5449_7);

wire[31:0] addr_5450_7;

Selector_2 s5450_7(wires_1362_6[2], addr_1362_6, addr_positional[21803:21800], addr_5450_7);

wire[31:0] addr_5451_7;

Selector_2 s5451_7(wires_1362_6[3], addr_1362_6, addr_positional[21807:21804], addr_5451_7);

wire[31:0] addr_5452_7;

Selector_2 s5452_7(wires_1363_6[0], addr_1363_6, addr_positional[21811:21808], addr_5452_7);

wire[31:0] addr_5453_7;

Selector_2 s5453_7(wires_1363_6[1], addr_1363_6, addr_positional[21815:21812], addr_5453_7);

wire[31:0] addr_5454_7;

Selector_2 s5454_7(wires_1363_6[2], addr_1363_6, addr_positional[21819:21816], addr_5454_7);

wire[31:0] addr_5455_7;

Selector_2 s5455_7(wires_1363_6[3], addr_1363_6, addr_positional[21823:21820], addr_5455_7);

wire[31:0] addr_5456_7;

Selector_2 s5456_7(wires_1364_6[0], addr_1364_6, addr_positional[21827:21824], addr_5456_7);

wire[31:0] addr_5457_7;

Selector_2 s5457_7(wires_1364_6[1], addr_1364_6, addr_positional[21831:21828], addr_5457_7);

wire[31:0] addr_5458_7;

Selector_2 s5458_7(wires_1364_6[2], addr_1364_6, addr_positional[21835:21832], addr_5458_7);

wire[31:0] addr_5459_7;

Selector_2 s5459_7(wires_1364_6[3], addr_1364_6, addr_positional[21839:21836], addr_5459_7);

wire[31:0] addr_5460_7;

Selector_2 s5460_7(wires_1365_6[0], addr_1365_6, addr_positional[21843:21840], addr_5460_7);

wire[31:0] addr_5461_7;

Selector_2 s5461_7(wires_1365_6[1], addr_1365_6, addr_positional[21847:21844], addr_5461_7);

wire[31:0] addr_5462_7;

Selector_2 s5462_7(wires_1365_6[2], addr_1365_6, addr_positional[21851:21848], addr_5462_7);

wire[31:0] addr_5463_7;

Selector_2 s5463_7(wires_1365_6[3], addr_1365_6, addr_positional[21855:21852], addr_5463_7);

wire[31:0] addr_5464_7;

Selector_2 s5464_7(wires_1366_6[0], addr_1366_6, addr_positional[21859:21856], addr_5464_7);

wire[31:0] addr_5465_7;

Selector_2 s5465_7(wires_1366_6[1], addr_1366_6, addr_positional[21863:21860], addr_5465_7);

wire[31:0] addr_5466_7;

Selector_2 s5466_7(wires_1366_6[2], addr_1366_6, addr_positional[21867:21864], addr_5466_7);

wire[31:0] addr_5467_7;

Selector_2 s5467_7(wires_1366_6[3], addr_1366_6, addr_positional[21871:21868], addr_5467_7);

wire[31:0] addr_5468_7;

Selector_2 s5468_7(wires_1367_6[0], addr_1367_6, addr_positional[21875:21872], addr_5468_7);

wire[31:0] addr_5469_7;

Selector_2 s5469_7(wires_1367_6[1], addr_1367_6, addr_positional[21879:21876], addr_5469_7);

wire[31:0] addr_5470_7;

Selector_2 s5470_7(wires_1367_6[2], addr_1367_6, addr_positional[21883:21880], addr_5470_7);

wire[31:0] addr_5471_7;

Selector_2 s5471_7(wires_1367_6[3], addr_1367_6, addr_positional[21887:21884], addr_5471_7);

wire[31:0] addr_5472_7;

Selector_2 s5472_7(wires_1368_6[0], addr_1368_6, addr_positional[21891:21888], addr_5472_7);

wire[31:0] addr_5473_7;

Selector_2 s5473_7(wires_1368_6[1], addr_1368_6, addr_positional[21895:21892], addr_5473_7);

wire[31:0] addr_5474_7;

Selector_2 s5474_7(wires_1368_6[2], addr_1368_6, addr_positional[21899:21896], addr_5474_7);

wire[31:0] addr_5475_7;

Selector_2 s5475_7(wires_1368_6[3], addr_1368_6, addr_positional[21903:21900], addr_5475_7);

wire[31:0] addr_5476_7;

Selector_2 s5476_7(wires_1369_6[0], addr_1369_6, addr_positional[21907:21904], addr_5476_7);

wire[31:0] addr_5477_7;

Selector_2 s5477_7(wires_1369_6[1], addr_1369_6, addr_positional[21911:21908], addr_5477_7);

wire[31:0] addr_5478_7;

Selector_2 s5478_7(wires_1369_6[2], addr_1369_6, addr_positional[21915:21912], addr_5478_7);

wire[31:0] addr_5479_7;

Selector_2 s5479_7(wires_1369_6[3], addr_1369_6, addr_positional[21919:21916], addr_5479_7);

wire[31:0] addr_5480_7;

Selector_2 s5480_7(wires_1370_6[0], addr_1370_6, addr_positional[21923:21920], addr_5480_7);

wire[31:0] addr_5481_7;

Selector_2 s5481_7(wires_1370_6[1], addr_1370_6, addr_positional[21927:21924], addr_5481_7);

wire[31:0] addr_5482_7;

Selector_2 s5482_7(wires_1370_6[2], addr_1370_6, addr_positional[21931:21928], addr_5482_7);

wire[31:0] addr_5483_7;

Selector_2 s5483_7(wires_1370_6[3], addr_1370_6, addr_positional[21935:21932], addr_5483_7);

wire[31:0] addr_5484_7;

Selector_2 s5484_7(wires_1371_6[0], addr_1371_6, addr_positional[21939:21936], addr_5484_7);

wire[31:0] addr_5485_7;

Selector_2 s5485_7(wires_1371_6[1], addr_1371_6, addr_positional[21943:21940], addr_5485_7);

wire[31:0] addr_5486_7;

Selector_2 s5486_7(wires_1371_6[2], addr_1371_6, addr_positional[21947:21944], addr_5486_7);

wire[31:0] addr_5487_7;

Selector_2 s5487_7(wires_1371_6[3], addr_1371_6, addr_positional[21951:21948], addr_5487_7);

wire[31:0] addr_5488_7;

Selector_2 s5488_7(wires_1372_6[0], addr_1372_6, addr_positional[21955:21952], addr_5488_7);

wire[31:0] addr_5489_7;

Selector_2 s5489_7(wires_1372_6[1], addr_1372_6, addr_positional[21959:21956], addr_5489_7);

wire[31:0] addr_5490_7;

Selector_2 s5490_7(wires_1372_6[2], addr_1372_6, addr_positional[21963:21960], addr_5490_7);

wire[31:0] addr_5491_7;

Selector_2 s5491_7(wires_1372_6[3], addr_1372_6, addr_positional[21967:21964], addr_5491_7);

wire[31:0] addr_5492_7;

Selector_2 s5492_7(wires_1373_6[0], addr_1373_6, addr_positional[21971:21968], addr_5492_7);

wire[31:0] addr_5493_7;

Selector_2 s5493_7(wires_1373_6[1], addr_1373_6, addr_positional[21975:21972], addr_5493_7);

wire[31:0] addr_5494_7;

Selector_2 s5494_7(wires_1373_6[2], addr_1373_6, addr_positional[21979:21976], addr_5494_7);

wire[31:0] addr_5495_7;

Selector_2 s5495_7(wires_1373_6[3], addr_1373_6, addr_positional[21983:21980], addr_5495_7);

wire[31:0] addr_5496_7;

Selector_2 s5496_7(wires_1374_6[0], addr_1374_6, addr_positional[21987:21984], addr_5496_7);

wire[31:0] addr_5497_7;

Selector_2 s5497_7(wires_1374_6[1], addr_1374_6, addr_positional[21991:21988], addr_5497_7);

wire[31:0] addr_5498_7;

Selector_2 s5498_7(wires_1374_6[2], addr_1374_6, addr_positional[21995:21992], addr_5498_7);

wire[31:0] addr_5499_7;

Selector_2 s5499_7(wires_1374_6[3], addr_1374_6, addr_positional[21999:21996], addr_5499_7);

wire[31:0] addr_5500_7;

Selector_2 s5500_7(wires_1375_6[0], addr_1375_6, addr_positional[22003:22000], addr_5500_7);

wire[31:0] addr_5501_7;

Selector_2 s5501_7(wires_1375_6[1], addr_1375_6, addr_positional[22007:22004], addr_5501_7);

wire[31:0] addr_5502_7;

Selector_2 s5502_7(wires_1375_6[2], addr_1375_6, addr_positional[22011:22008], addr_5502_7);

wire[31:0] addr_5503_7;

Selector_2 s5503_7(wires_1375_6[3], addr_1375_6, addr_positional[22015:22012], addr_5503_7);

wire[31:0] addr_5504_7;

Selector_2 s5504_7(wires_1376_6[0], addr_1376_6, addr_positional[22019:22016], addr_5504_7);

wire[31:0] addr_5505_7;

Selector_2 s5505_7(wires_1376_6[1], addr_1376_6, addr_positional[22023:22020], addr_5505_7);

wire[31:0] addr_5506_7;

Selector_2 s5506_7(wires_1376_6[2], addr_1376_6, addr_positional[22027:22024], addr_5506_7);

wire[31:0] addr_5507_7;

Selector_2 s5507_7(wires_1376_6[3], addr_1376_6, addr_positional[22031:22028], addr_5507_7);

wire[31:0] addr_5508_7;

Selector_2 s5508_7(wires_1377_6[0], addr_1377_6, addr_positional[22035:22032], addr_5508_7);

wire[31:0] addr_5509_7;

Selector_2 s5509_7(wires_1377_6[1], addr_1377_6, addr_positional[22039:22036], addr_5509_7);

wire[31:0] addr_5510_7;

Selector_2 s5510_7(wires_1377_6[2], addr_1377_6, addr_positional[22043:22040], addr_5510_7);

wire[31:0] addr_5511_7;

Selector_2 s5511_7(wires_1377_6[3], addr_1377_6, addr_positional[22047:22044], addr_5511_7);

wire[31:0] addr_5512_7;

Selector_2 s5512_7(wires_1378_6[0], addr_1378_6, addr_positional[22051:22048], addr_5512_7);

wire[31:0] addr_5513_7;

Selector_2 s5513_7(wires_1378_6[1], addr_1378_6, addr_positional[22055:22052], addr_5513_7);

wire[31:0] addr_5514_7;

Selector_2 s5514_7(wires_1378_6[2], addr_1378_6, addr_positional[22059:22056], addr_5514_7);

wire[31:0] addr_5515_7;

Selector_2 s5515_7(wires_1378_6[3], addr_1378_6, addr_positional[22063:22060], addr_5515_7);

wire[31:0] addr_5516_7;

Selector_2 s5516_7(wires_1379_6[0], addr_1379_6, addr_positional[22067:22064], addr_5516_7);

wire[31:0] addr_5517_7;

Selector_2 s5517_7(wires_1379_6[1], addr_1379_6, addr_positional[22071:22068], addr_5517_7);

wire[31:0] addr_5518_7;

Selector_2 s5518_7(wires_1379_6[2], addr_1379_6, addr_positional[22075:22072], addr_5518_7);

wire[31:0] addr_5519_7;

Selector_2 s5519_7(wires_1379_6[3], addr_1379_6, addr_positional[22079:22076], addr_5519_7);

wire[31:0] addr_5520_7;

Selector_2 s5520_7(wires_1380_6[0], addr_1380_6, addr_positional[22083:22080], addr_5520_7);

wire[31:0] addr_5521_7;

Selector_2 s5521_7(wires_1380_6[1], addr_1380_6, addr_positional[22087:22084], addr_5521_7);

wire[31:0] addr_5522_7;

Selector_2 s5522_7(wires_1380_6[2], addr_1380_6, addr_positional[22091:22088], addr_5522_7);

wire[31:0] addr_5523_7;

Selector_2 s5523_7(wires_1380_6[3], addr_1380_6, addr_positional[22095:22092], addr_5523_7);

wire[31:0] addr_5524_7;

Selector_2 s5524_7(wires_1381_6[0], addr_1381_6, addr_positional[22099:22096], addr_5524_7);

wire[31:0] addr_5525_7;

Selector_2 s5525_7(wires_1381_6[1], addr_1381_6, addr_positional[22103:22100], addr_5525_7);

wire[31:0] addr_5526_7;

Selector_2 s5526_7(wires_1381_6[2], addr_1381_6, addr_positional[22107:22104], addr_5526_7);

wire[31:0] addr_5527_7;

Selector_2 s5527_7(wires_1381_6[3], addr_1381_6, addr_positional[22111:22108], addr_5527_7);

wire[31:0] addr_5528_7;

Selector_2 s5528_7(wires_1382_6[0], addr_1382_6, addr_positional[22115:22112], addr_5528_7);

wire[31:0] addr_5529_7;

Selector_2 s5529_7(wires_1382_6[1], addr_1382_6, addr_positional[22119:22116], addr_5529_7);

wire[31:0] addr_5530_7;

Selector_2 s5530_7(wires_1382_6[2], addr_1382_6, addr_positional[22123:22120], addr_5530_7);

wire[31:0] addr_5531_7;

Selector_2 s5531_7(wires_1382_6[3], addr_1382_6, addr_positional[22127:22124], addr_5531_7);

wire[31:0] addr_5532_7;

Selector_2 s5532_7(wires_1383_6[0], addr_1383_6, addr_positional[22131:22128], addr_5532_7);

wire[31:0] addr_5533_7;

Selector_2 s5533_7(wires_1383_6[1], addr_1383_6, addr_positional[22135:22132], addr_5533_7);

wire[31:0] addr_5534_7;

Selector_2 s5534_7(wires_1383_6[2], addr_1383_6, addr_positional[22139:22136], addr_5534_7);

wire[31:0] addr_5535_7;

Selector_2 s5535_7(wires_1383_6[3], addr_1383_6, addr_positional[22143:22140], addr_5535_7);

wire[31:0] addr_5536_7;

Selector_2 s5536_7(wires_1384_6[0], addr_1384_6, addr_positional[22147:22144], addr_5536_7);

wire[31:0] addr_5537_7;

Selector_2 s5537_7(wires_1384_6[1], addr_1384_6, addr_positional[22151:22148], addr_5537_7);

wire[31:0] addr_5538_7;

Selector_2 s5538_7(wires_1384_6[2], addr_1384_6, addr_positional[22155:22152], addr_5538_7);

wire[31:0] addr_5539_7;

Selector_2 s5539_7(wires_1384_6[3], addr_1384_6, addr_positional[22159:22156], addr_5539_7);

wire[31:0] addr_5540_7;

Selector_2 s5540_7(wires_1385_6[0], addr_1385_6, addr_positional[22163:22160], addr_5540_7);

wire[31:0] addr_5541_7;

Selector_2 s5541_7(wires_1385_6[1], addr_1385_6, addr_positional[22167:22164], addr_5541_7);

wire[31:0] addr_5542_7;

Selector_2 s5542_7(wires_1385_6[2], addr_1385_6, addr_positional[22171:22168], addr_5542_7);

wire[31:0] addr_5543_7;

Selector_2 s5543_7(wires_1385_6[3], addr_1385_6, addr_positional[22175:22172], addr_5543_7);

wire[31:0] addr_5544_7;

Selector_2 s5544_7(wires_1386_6[0], addr_1386_6, addr_positional[22179:22176], addr_5544_7);

wire[31:0] addr_5545_7;

Selector_2 s5545_7(wires_1386_6[1], addr_1386_6, addr_positional[22183:22180], addr_5545_7);

wire[31:0] addr_5546_7;

Selector_2 s5546_7(wires_1386_6[2], addr_1386_6, addr_positional[22187:22184], addr_5546_7);

wire[31:0] addr_5547_7;

Selector_2 s5547_7(wires_1386_6[3], addr_1386_6, addr_positional[22191:22188], addr_5547_7);

wire[31:0] addr_5548_7;

Selector_2 s5548_7(wires_1387_6[0], addr_1387_6, addr_positional[22195:22192], addr_5548_7);

wire[31:0] addr_5549_7;

Selector_2 s5549_7(wires_1387_6[1], addr_1387_6, addr_positional[22199:22196], addr_5549_7);

wire[31:0] addr_5550_7;

Selector_2 s5550_7(wires_1387_6[2], addr_1387_6, addr_positional[22203:22200], addr_5550_7);

wire[31:0] addr_5551_7;

Selector_2 s5551_7(wires_1387_6[3], addr_1387_6, addr_positional[22207:22204], addr_5551_7);

wire[31:0] addr_5552_7;

Selector_2 s5552_7(wires_1388_6[0], addr_1388_6, addr_positional[22211:22208], addr_5552_7);

wire[31:0] addr_5553_7;

Selector_2 s5553_7(wires_1388_6[1], addr_1388_6, addr_positional[22215:22212], addr_5553_7);

wire[31:0] addr_5554_7;

Selector_2 s5554_7(wires_1388_6[2], addr_1388_6, addr_positional[22219:22216], addr_5554_7);

wire[31:0] addr_5555_7;

Selector_2 s5555_7(wires_1388_6[3], addr_1388_6, addr_positional[22223:22220], addr_5555_7);

wire[31:0] addr_5556_7;

Selector_2 s5556_7(wires_1389_6[0], addr_1389_6, addr_positional[22227:22224], addr_5556_7);

wire[31:0] addr_5557_7;

Selector_2 s5557_7(wires_1389_6[1], addr_1389_6, addr_positional[22231:22228], addr_5557_7);

wire[31:0] addr_5558_7;

Selector_2 s5558_7(wires_1389_6[2], addr_1389_6, addr_positional[22235:22232], addr_5558_7);

wire[31:0] addr_5559_7;

Selector_2 s5559_7(wires_1389_6[3], addr_1389_6, addr_positional[22239:22236], addr_5559_7);

wire[31:0] addr_5560_7;

Selector_2 s5560_7(wires_1390_6[0], addr_1390_6, addr_positional[22243:22240], addr_5560_7);

wire[31:0] addr_5561_7;

Selector_2 s5561_7(wires_1390_6[1], addr_1390_6, addr_positional[22247:22244], addr_5561_7);

wire[31:0] addr_5562_7;

Selector_2 s5562_7(wires_1390_6[2], addr_1390_6, addr_positional[22251:22248], addr_5562_7);

wire[31:0] addr_5563_7;

Selector_2 s5563_7(wires_1390_6[3], addr_1390_6, addr_positional[22255:22252], addr_5563_7);

wire[31:0] addr_5564_7;

Selector_2 s5564_7(wires_1391_6[0], addr_1391_6, addr_positional[22259:22256], addr_5564_7);

wire[31:0] addr_5565_7;

Selector_2 s5565_7(wires_1391_6[1], addr_1391_6, addr_positional[22263:22260], addr_5565_7);

wire[31:0] addr_5566_7;

Selector_2 s5566_7(wires_1391_6[2], addr_1391_6, addr_positional[22267:22264], addr_5566_7);

wire[31:0] addr_5567_7;

Selector_2 s5567_7(wires_1391_6[3], addr_1391_6, addr_positional[22271:22268], addr_5567_7);

wire[31:0] addr_5568_7;

Selector_2 s5568_7(wires_1392_6[0], addr_1392_6, addr_positional[22275:22272], addr_5568_7);

wire[31:0] addr_5569_7;

Selector_2 s5569_7(wires_1392_6[1], addr_1392_6, addr_positional[22279:22276], addr_5569_7);

wire[31:0] addr_5570_7;

Selector_2 s5570_7(wires_1392_6[2], addr_1392_6, addr_positional[22283:22280], addr_5570_7);

wire[31:0] addr_5571_7;

Selector_2 s5571_7(wires_1392_6[3], addr_1392_6, addr_positional[22287:22284], addr_5571_7);

wire[31:0] addr_5572_7;

Selector_2 s5572_7(wires_1393_6[0], addr_1393_6, addr_positional[22291:22288], addr_5572_7);

wire[31:0] addr_5573_7;

Selector_2 s5573_7(wires_1393_6[1], addr_1393_6, addr_positional[22295:22292], addr_5573_7);

wire[31:0] addr_5574_7;

Selector_2 s5574_7(wires_1393_6[2], addr_1393_6, addr_positional[22299:22296], addr_5574_7);

wire[31:0] addr_5575_7;

Selector_2 s5575_7(wires_1393_6[3], addr_1393_6, addr_positional[22303:22300], addr_5575_7);

wire[31:0] addr_5576_7;

Selector_2 s5576_7(wires_1394_6[0], addr_1394_6, addr_positional[22307:22304], addr_5576_7);

wire[31:0] addr_5577_7;

Selector_2 s5577_7(wires_1394_6[1], addr_1394_6, addr_positional[22311:22308], addr_5577_7);

wire[31:0] addr_5578_7;

Selector_2 s5578_7(wires_1394_6[2], addr_1394_6, addr_positional[22315:22312], addr_5578_7);

wire[31:0] addr_5579_7;

Selector_2 s5579_7(wires_1394_6[3], addr_1394_6, addr_positional[22319:22316], addr_5579_7);

wire[31:0] addr_5580_7;

Selector_2 s5580_7(wires_1395_6[0], addr_1395_6, addr_positional[22323:22320], addr_5580_7);

wire[31:0] addr_5581_7;

Selector_2 s5581_7(wires_1395_6[1], addr_1395_6, addr_positional[22327:22324], addr_5581_7);

wire[31:0] addr_5582_7;

Selector_2 s5582_7(wires_1395_6[2], addr_1395_6, addr_positional[22331:22328], addr_5582_7);

wire[31:0] addr_5583_7;

Selector_2 s5583_7(wires_1395_6[3], addr_1395_6, addr_positional[22335:22332], addr_5583_7);

wire[31:0] addr_5584_7;

Selector_2 s5584_7(wires_1396_6[0], addr_1396_6, addr_positional[22339:22336], addr_5584_7);

wire[31:0] addr_5585_7;

Selector_2 s5585_7(wires_1396_6[1], addr_1396_6, addr_positional[22343:22340], addr_5585_7);

wire[31:0] addr_5586_7;

Selector_2 s5586_7(wires_1396_6[2], addr_1396_6, addr_positional[22347:22344], addr_5586_7);

wire[31:0] addr_5587_7;

Selector_2 s5587_7(wires_1396_6[3], addr_1396_6, addr_positional[22351:22348], addr_5587_7);

wire[31:0] addr_5588_7;

Selector_2 s5588_7(wires_1397_6[0], addr_1397_6, addr_positional[22355:22352], addr_5588_7);

wire[31:0] addr_5589_7;

Selector_2 s5589_7(wires_1397_6[1], addr_1397_6, addr_positional[22359:22356], addr_5589_7);

wire[31:0] addr_5590_7;

Selector_2 s5590_7(wires_1397_6[2], addr_1397_6, addr_positional[22363:22360], addr_5590_7);

wire[31:0] addr_5591_7;

Selector_2 s5591_7(wires_1397_6[3], addr_1397_6, addr_positional[22367:22364], addr_5591_7);

wire[31:0] addr_5592_7;

Selector_2 s5592_7(wires_1398_6[0], addr_1398_6, addr_positional[22371:22368], addr_5592_7);

wire[31:0] addr_5593_7;

Selector_2 s5593_7(wires_1398_6[1], addr_1398_6, addr_positional[22375:22372], addr_5593_7);

wire[31:0] addr_5594_7;

Selector_2 s5594_7(wires_1398_6[2], addr_1398_6, addr_positional[22379:22376], addr_5594_7);

wire[31:0] addr_5595_7;

Selector_2 s5595_7(wires_1398_6[3], addr_1398_6, addr_positional[22383:22380], addr_5595_7);

wire[31:0] addr_5596_7;

Selector_2 s5596_7(wires_1399_6[0], addr_1399_6, addr_positional[22387:22384], addr_5596_7);

wire[31:0] addr_5597_7;

Selector_2 s5597_7(wires_1399_6[1], addr_1399_6, addr_positional[22391:22388], addr_5597_7);

wire[31:0] addr_5598_7;

Selector_2 s5598_7(wires_1399_6[2], addr_1399_6, addr_positional[22395:22392], addr_5598_7);

wire[31:0] addr_5599_7;

Selector_2 s5599_7(wires_1399_6[3], addr_1399_6, addr_positional[22399:22396], addr_5599_7);

wire[31:0] addr_5600_7;

Selector_2 s5600_7(wires_1400_6[0], addr_1400_6, addr_positional[22403:22400], addr_5600_7);

wire[31:0] addr_5601_7;

Selector_2 s5601_7(wires_1400_6[1], addr_1400_6, addr_positional[22407:22404], addr_5601_7);

wire[31:0] addr_5602_7;

Selector_2 s5602_7(wires_1400_6[2], addr_1400_6, addr_positional[22411:22408], addr_5602_7);

wire[31:0] addr_5603_7;

Selector_2 s5603_7(wires_1400_6[3], addr_1400_6, addr_positional[22415:22412], addr_5603_7);

wire[31:0] addr_5604_7;

Selector_2 s5604_7(wires_1401_6[0], addr_1401_6, addr_positional[22419:22416], addr_5604_7);

wire[31:0] addr_5605_7;

Selector_2 s5605_7(wires_1401_6[1], addr_1401_6, addr_positional[22423:22420], addr_5605_7);

wire[31:0] addr_5606_7;

Selector_2 s5606_7(wires_1401_6[2], addr_1401_6, addr_positional[22427:22424], addr_5606_7);

wire[31:0] addr_5607_7;

Selector_2 s5607_7(wires_1401_6[3], addr_1401_6, addr_positional[22431:22428], addr_5607_7);

wire[31:0] addr_5608_7;

Selector_2 s5608_7(wires_1402_6[0], addr_1402_6, addr_positional[22435:22432], addr_5608_7);

wire[31:0] addr_5609_7;

Selector_2 s5609_7(wires_1402_6[1], addr_1402_6, addr_positional[22439:22436], addr_5609_7);

wire[31:0] addr_5610_7;

Selector_2 s5610_7(wires_1402_6[2], addr_1402_6, addr_positional[22443:22440], addr_5610_7);

wire[31:0] addr_5611_7;

Selector_2 s5611_7(wires_1402_6[3], addr_1402_6, addr_positional[22447:22444], addr_5611_7);

wire[31:0] addr_5612_7;

Selector_2 s5612_7(wires_1403_6[0], addr_1403_6, addr_positional[22451:22448], addr_5612_7);

wire[31:0] addr_5613_7;

Selector_2 s5613_7(wires_1403_6[1], addr_1403_6, addr_positional[22455:22452], addr_5613_7);

wire[31:0] addr_5614_7;

Selector_2 s5614_7(wires_1403_6[2], addr_1403_6, addr_positional[22459:22456], addr_5614_7);

wire[31:0] addr_5615_7;

Selector_2 s5615_7(wires_1403_6[3], addr_1403_6, addr_positional[22463:22460], addr_5615_7);

wire[31:0] addr_5616_7;

Selector_2 s5616_7(wires_1404_6[0], addr_1404_6, addr_positional[22467:22464], addr_5616_7);

wire[31:0] addr_5617_7;

Selector_2 s5617_7(wires_1404_6[1], addr_1404_6, addr_positional[22471:22468], addr_5617_7);

wire[31:0] addr_5618_7;

Selector_2 s5618_7(wires_1404_6[2], addr_1404_6, addr_positional[22475:22472], addr_5618_7);

wire[31:0] addr_5619_7;

Selector_2 s5619_7(wires_1404_6[3], addr_1404_6, addr_positional[22479:22476], addr_5619_7);

wire[31:0] addr_5620_7;

Selector_2 s5620_7(wires_1405_6[0], addr_1405_6, addr_positional[22483:22480], addr_5620_7);

wire[31:0] addr_5621_7;

Selector_2 s5621_7(wires_1405_6[1], addr_1405_6, addr_positional[22487:22484], addr_5621_7);

wire[31:0] addr_5622_7;

Selector_2 s5622_7(wires_1405_6[2], addr_1405_6, addr_positional[22491:22488], addr_5622_7);

wire[31:0] addr_5623_7;

Selector_2 s5623_7(wires_1405_6[3], addr_1405_6, addr_positional[22495:22492], addr_5623_7);

wire[31:0] addr_5624_7;

Selector_2 s5624_7(wires_1406_6[0], addr_1406_6, addr_positional[22499:22496], addr_5624_7);

wire[31:0] addr_5625_7;

Selector_2 s5625_7(wires_1406_6[1], addr_1406_6, addr_positional[22503:22500], addr_5625_7);

wire[31:0] addr_5626_7;

Selector_2 s5626_7(wires_1406_6[2], addr_1406_6, addr_positional[22507:22504], addr_5626_7);

wire[31:0] addr_5627_7;

Selector_2 s5627_7(wires_1406_6[3], addr_1406_6, addr_positional[22511:22508], addr_5627_7);

wire[31:0] addr_5628_7;

Selector_2 s5628_7(wires_1407_6[0], addr_1407_6, addr_positional[22515:22512], addr_5628_7);

wire[31:0] addr_5629_7;

Selector_2 s5629_7(wires_1407_6[1], addr_1407_6, addr_positional[22519:22516], addr_5629_7);

wire[31:0] addr_5630_7;

Selector_2 s5630_7(wires_1407_6[2], addr_1407_6, addr_positional[22523:22520], addr_5630_7);

wire[31:0] addr_5631_7;

Selector_2 s5631_7(wires_1407_6[3], addr_1407_6, addr_positional[22527:22524], addr_5631_7);

wire[31:0] addr_5632_7;

Selector_2 s5632_7(wires_1408_6[0], addr_1408_6, addr_positional[22531:22528], addr_5632_7);

wire[31:0] addr_5633_7;

Selector_2 s5633_7(wires_1408_6[1], addr_1408_6, addr_positional[22535:22532], addr_5633_7);

wire[31:0] addr_5634_7;

Selector_2 s5634_7(wires_1408_6[2], addr_1408_6, addr_positional[22539:22536], addr_5634_7);

wire[31:0] addr_5635_7;

Selector_2 s5635_7(wires_1408_6[3], addr_1408_6, addr_positional[22543:22540], addr_5635_7);

wire[31:0] addr_5636_7;

Selector_2 s5636_7(wires_1409_6[0], addr_1409_6, addr_positional[22547:22544], addr_5636_7);

wire[31:0] addr_5637_7;

Selector_2 s5637_7(wires_1409_6[1], addr_1409_6, addr_positional[22551:22548], addr_5637_7);

wire[31:0] addr_5638_7;

Selector_2 s5638_7(wires_1409_6[2], addr_1409_6, addr_positional[22555:22552], addr_5638_7);

wire[31:0] addr_5639_7;

Selector_2 s5639_7(wires_1409_6[3], addr_1409_6, addr_positional[22559:22556], addr_5639_7);

wire[31:0] addr_5640_7;

Selector_2 s5640_7(wires_1410_6[0], addr_1410_6, addr_positional[22563:22560], addr_5640_7);

wire[31:0] addr_5641_7;

Selector_2 s5641_7(wires_1410_6[1], addr_1410_6, addr_positional[22567:22564], addr_5641_7);

wire[31:0] addr_5642_7;

Selector_2 s5642_7(wires_1410_6[2], addr_1410_6, addr_positional[22571:22568], addr_5642_7);

wire[31:0] addr_5643_7;

Selector_2 s5643_7(wires_1410_6[3], addr_1410_6, addr_positional[22575:22572], addr_5643_7);

wire[31:0] addr_5644_7;

Selector_2 s5644_7(wires_1411_6[0], addr_1411_6, addr_positional[22579:22576], addr_5644_7);

wire[31:0] addr_5645_7;

Selector_2 s5645_7(wires_1411_6[1], addr_1411_6, addr_positional[22583:22580], addr_5645_7);

wire[31:0] addr_5646_7;

Selector_2 s5646_7(wires_1411_6[2], addr_1411_6, addr_positional[22587:22584], addr_5646_7);

wire[31:0] addr_5647_7;

Selector_2 s5647_7(wires_1411_6[3], addr_1411_6, addr_positional[22591:22588], addr_5647_7);

wire[31:0] addr_5648_7;

Selector_2 s5648_7(wires_1412_6[0], addr_1412_6, addr_positional[22595:22592], addr_5648_7);

wire[31:0] addr_5649_7;

Selector_2 s5649_7(wires_1412_6[1], addr_1412_6, addr_positional[22599:22596], addr_5649_7);

wire[31:0] addr_5650_7;

Selector_2 s5650_7(wires_1412_6[2], addr_1412_6, addr_positional[22603:22600], addr_5650_7);

wire[31:0] addr_5651_7;

Selector_2 s5651_7(wires_1412_6[3], addr_1412_6, addr_positional[22607:22604], addr_5651_7);

wire[31:0] addr_5652_7;

Selector_2 s5652_7(wires_1413_6[0], addr_1413_6, addr_positional[22611:22608], addr_5652_7);

wire[31:0] addr_5653_7;

Selector_2 s5653_7(wires_1413_6[1], addr_1413_6, addr_positional[22615:22612], addr_5653_7);

wire[31:0] addr_5654_7;

Selector_2 s5654_7(wires_1413_6[2], addr_1413_6, addr_positional[22619:22616], addr_5654_7);

wire[31:0] addr_5655_7;

Selector_2 s5655_7(wires_1413_6[3], addr_1413_6, addr_positional[22623:22620], addr_5655_7);

wire[31:0] addr_5656_7;

Selector_2 s5656_7(wires_1414_6[0], addr_1414_6, addr_positional[22627:22624], addr_5656_7);

wire[31:0] addr_5657_7;

Selector_2 s5657_7(wires_1414_6[1], addr_1414_6, addr_positional[22631:22628], addr_5657_7);

wire[31:0] addr_5658_7;

Selector_2 s5658_7(wires_1414_6[2], addr_1414_6, addr_positional[22635:22632], addr_5658_7);

wire[31:0] addr_5659_7;

Selector_2 s5659_7(wires_1414_6[3], addr_1414_6, addr_positional[22639:22636], addr_5659_7);

wire[31:0] addr_5660_7;

Selector_2 s5660_7(wires_1415_6[0], addr_1415_6, addr_positional[22643:22640], addr_5660_7);

wire[31:0] addr_5661_7;

Selector_2 s5661_7(wires_1415_6[1], addr_1415_6, addr_positional[22647:22644], addr_5661_7);

wire[31:0] addr_5662_7;

Selector_2 s5662_7(wires_1415_6[2], addr_1415_6, addr_positional[22651:22648], addr_5662_7);

wire[31:0] addr_5663_7;

Selector_2 s5663_7(wires_1415_6[3], addr_1415_6, addr_positional[22655:22652], addr_5663_7);

wire[31:0] addr_5664_7;

Selector_2 s5664_7(wires_1416_6[0], addr_1416_6, addr_positional[22659:22656], addr_5664_7);

wire[31:0] addr_5665_7;

Selector_2 s5665_7(wires_1416_6[1], addr_1416_6, addr_positional[22663:22660], addr_5665_7);

wire[31:0] addr_5666_7;

Selector_2 s5666_7(wires_1416_6[2], addr_1416_6, addr_positional[22667:22664], addr_5666_7);

wire[31:0] addr_5667_7;

Selector_2 s5667_7(wires_1416_6[3], addr_1416_6, addr_positional[22671:22668], addr_5667_7);

wire[31:0] addr_5668_7;

Selector_2 s5668_7(wires_1417_6[0], addr_1417_6, addr_positional[22675:22672], addr_5668_7);

wire[31:0] addr_5669_7;

Selector_2 s5669_7(wires_1417_6[1], addr_1417_6, addr_positional[22679:22676], addr_5669_7);

wire[31:0] addr_5670_7;

Selector_2 s5670_7(wires_1417_6[2], addr_1417_6, addr_positional[22683:22680], addr_5670_7);

wire[31:0] addr_5671_7;

Selector_2 s5671_7(wires_1417_6[3], addr_1417_6, addr_positional[22687:22684], addr_5671_7);

wire[31:0] addr_5672_7;

Selector_2 s5672_7(wires_1418_6[0], addr_1418_6, addr_positional[22691:22688], addr_5672_7);

wire[31:0] addr_5673_7;

Selector_2 s5673_7(wires_1418_6[1], addr_1418_6, addr_positional[22695:22692], addr_5673_7);

wire[31:0] addr_5674_7;

Selector_2 s5674_7(wires_1418_6[2], addr_1418_6, addr_positional[22699:22696], addr_5674_7);

wire[31:0] addr_5675_7;

Selector_2 s5675_7(wires_1418_6[3], addr_1418_6, addr_positional[22703:22700], addr_5675_7);

wire[31:0] addr_5676_7;

Selector_2 s5676_7(wires_1419_6[0], addr_1419_6, addr_positional[22707:22704], addr_5676_7);

wire[31:0] addr_5677_7;

Selector_2 s5677_7(wires_1419_6[1], addr_1419_6, addr_positional[22711:22708], addr_5677_7);

wire[31:0] addr_5678_7;

Selector_2 s5678_7(wires_1419_6[2], addr_1419_6, addr_positional[22715:22712], addr_5678_7);

wire[31:0] addr_5679_7;

Selector_2 s5679_7(wires_1419_6[3], addr_1419_6, addr_positional[22719:22716], addr_5679_7);

wire[31:0] addr_5680_7;

Selector_2 s5680_7(wires_1420_6[0], addr_1420_6, addr_positional[22723:22720], addr_5680_7);

wire[31:0] addr_5681_7;

Selector_2 s5681_7(wires_1420_6[1], addr_1420_6, addr_positional[22727:22724], addr_5681_7);

wire[31:0] addr_5682_7;

Selector_2 s5682_7(wires_1420_6[2], addr_1420_6, addr_positional[22731:22728], addr_5682_7);

wire[31:0] addr_5683_7;

Selector_2 s5683_7(wires_1420_6[3], addr_1420_6, addr_positional[22735:22732], addr_5683_7);

wire[31:0] addr_5684_7;

Selector_2 s5684_7(wires_1421_6[0], addr_1421_6, addr_positional[22739:22736], addr_5684_7);

wire[31:0] addr_5685_7;

Selector_2 s5685_7(wires_1421_6[1], addr_1421_6, addr_positional[22743:22740], addr_5685_7);

wire[31:0] addr_5686_7;

Selector_2 s5686_7(wires_1421_6[2], addr_1421_6, addr_positional[22747:22744], addr_5686_7);

wire[31:0] addr_5687_7;

Selector_2 s5687_7(wires_1421_6[3], addr_1421_6, addr_positional[22751:22748], addr_5687_7);

wire[31:0] addr_5688_7;

Selector_2 s5688_7(wires_1422_6[0], addr_1422_6, addr_positional[22755:22752], addr_5688_7);

wire[31:0] addr_5689_7;

Selector_2 s5689_7(wires_1422_6[1], addr_1422_6, addr_positional[22759:22756], addr_5689_7);

wire[31:0] addr_5690_7;

Selector_2 s5690_7(wires_1422_6[2], addr_1422_6, addr_positional[22763:22760], addr_5690_7);

wire[31:0] addr_5691_7;

Selector_2 s5691_7(wires_1422_6[3], addr_1422_6, addr_positional[22767:22764], addr_5691_7);

wire[31:0] addr_5692_7;

Selector_2 s5692_7(wires_1423_6[0], addr_1423_6, addr_positional[22771:22768], addr_5692_7);

wire[31:0] addr_5693_7;

Selector_2 s5693_7(wires_1423_6[1], addr_1423_6, addr_positional[22775:22772], addr_5693_7);

wire[31:0] addr_5694_7;

Selector_2 s5694_7(wires_1423_6[2], addr_1423_6, addr_positional[22779:22776], addr_5694_7);

wire[31:0] addr_5695_7;

Selector_2 s5695_7(wires_1423_6[3], addr_1423_6, addr_positional[22783:22780], addr_5695_7);

wire[31:0] addr_5696_7;

Selector_2 s5696_7(wires_1424_6[0], addr_1424_6, addr_positional[22787:22784], addr_5696_7);

wire[31:0] addr_5697_7;

Selector_2 s5697_7(wires_1424_6[1], addr_1424_6, addr_positional[22791:22788], addr_5697_7);

wire[31:0] addr_5698_7;

Selector_2 s5698_7(wires_1424_6[2], addr_1424_6, addr_positional[22795:22792], addr_5698_7);

wire[31:0] addr_5699_7;

Selector_2 s5699_7(wires_1424_6[3], addr_1424_6, addr_positional[22799:22796], addr_5699_7);

wire[31:0] addr_5700_7;

Selector_2 s5700_7(wires_1425_6[0], addr_1425_6, addr_positional[22803:22800], addr_5700_7);

wire[31:0] addr_5701_7;

Selector_2 s5701_7(wires_1425_6[1], addr_1425_6, addr_positional[22807:22804], addr_5701_7);

wire[31:0] addr_5702_7;

Selector_2 s5702_7(wires_1425_6[2], addr_1425_6, addr_positional[22811:22808], addr_5702_7);

wire[31:0] addr_5703_7;

Selector_2 s5703_7(wires_1425_6[3], addr_1425_6, addr_positional[22815:22812], addr_5703_7);

wire[31:0] addr_5704_7;

Selector_2 s5704_7(wires_1426_6[0], addr_1426_6, addr_positional[22819:22816], addr_5704_7);

wire[31:0] addr_5705_7;

Selector_2 s5705_7(wires_1426_6[1], addr_1426_6, addr_positional[22823:22820], addr_5705_7);

wire[31:0] addr_5706_7;

Selector_2 s5706_7(wires_1426_6[2], addr_1426_6, addr_positional[22827:22824], addr_5706_7);

wire[31:0] addr_5707_7;

Selector_2 s5707_7(wires_1426_6[3], addr_1426_6, addr_positional[22831:22828], addr_5707_7);

wire[31:0] addr_5708_7;

Selector_2 s5708_7(wires_1427_6[0], addr_1427_6, addr_positional[22835:22832], addr_5708_7);

wire[31:0] addr_5709_7;

Selector_2 s5709_7(wires_1427_6[1], addr_1427_6, addr_positional[22839:22836], addr_5709_7);

wire[31:0] addr_5710_7;

Selector_2 s5710_7(wires_1427_6[2], addr_1427_6, addr_positional[22843:22840], addr_5710_7);

wire[31:0] addr_5711_7;

Selector_2 s5711_7(wires_1427_6[3], addr_1427_6, addr_positional[22847:22844], addr_5711_7);

wire[31:0] addr_5712_7;

Selector_2 s5712_7(wires_1428_6[0], addr_1428_6, addr_positional[22851:22848], addr_5712_7);

wire[31:0] addr_5713_7;

Selector_2 s5713_7(wires_1428_6[1], addr_1428_6, addr_positional[22855:22852], addr_5713_7);

wire[31:0] addr_5714_7;

Selector_2 s5714_7(wires_1428_6[2], addr_1428_6, addr_positional[22859:22856], addr_5714_7);

wire[31:0] addr_5715_7;

Selector_2 s5715_7(wires_1428_6[3], addr_1428_6, addr_positional[22863:22860], addr_5715_7);

wire[31:0] addr_5716_7;

Selector_2 s5716_7(wires_1429_6[0], addr_1429_6, addr_positional[22867:22864], addr_5716_7);

wire[31:0] addr_5717_7;

Selector_2 s5717_7(wires_1429_6[1], addr_1429_6, addr_positional[22871:22868], addr_5717_7);

wire[31:0] addr_5718_7;

Selector_2 s5718_7(wires_1429_6[2], addr_1429_6, addr_positional[22875:22872], addr_5718_7);

wire[31:0] addr_5719_7;

Selector_2 s5719_7(wires_1429_6[3], addr_1429_6, addr_positional[22879:22876], addr_5719_7);

wire[31:0] addr_5720_7;

Selector_2 s5720_7(wires_1430_6[0], addr_1430_6, addr_positional[22883:22880], addr_5720_7);

wire[31:0] addr_5721_7;

Selector_2 s5721_7(wires_1430_6[1], addr_1430_6, addr_positional[22887:22884], addr_5721_7);

wire[31:0] addr_5722_7;

Selector_2 s5722_7(wires_1430_6[2], addr_1430_6, addr_positional[22891:22888], addr_5722_7);

wire[31:0] addr_5723_7;

Selector_2 s5723_7(wires_1430_6[3], addr_1430_6, addr_positional[22895:22892], addr_5723_7);

wire[31:0] addr_5724_7;

Selector_2 s5724_7(wires_1431_6[0], addr_1431_6, addr_positional[22899:22896], addr_5724_7);

wire[31:0] addr_5725_7;

Selector_2 s5725_7(wires_1431_6[1], addr_1431_6, addr_positional[22903:22900], addr_5725_7);

wire[31:0] addr_5726_7;

Selector_2 s5726_7(wires_1431_6[2], addr_1431_6, addr_positional[22907:22904], addr_5726_7);

wire[31:0] addr_5727_7;

Selector_2 s5727_7(wires_1431_6[3], addr_1431_6, addr_positional[22911:22908], addr_5727_7);

wire[31:0] addr_5728_7;

Selector_2 s5728_7(wires_1432_6[0], addr_1432_6, addr_positional[22915:22912], addr_5728_7);

wire[31:0] addr_5729_7;

Selector_2 s5729_7(wires_1432_6[1], addr_1432_6, addr_positional[22919:22916], addr_5729_7);

wire[31:0] addr_5730_7;

Selector_2 s5730_7(wires_1432_6[2], addr_1432_6, addr_positional[22923:22920], addr_5730_7);

wire[31:0] addr_5731_7;

Selector_2 s5731_7(wires_1432_6[3], addr_1432_6, addr_positional[22927:22924], addr_5731_7);

wire[31:0] addr_5732_7;

Selector_2 s5732_7(wires_1433_6[0], addr_1433_6, addr_positional[22931:22928], addr_5732_7);

wire[31:0] addr_5733_7;

Selector_2 s5733_7(wires_1433_6[1], addr_1433_6, addr_positional[22935:22932], addr_5733_7);

wire[31:0] addr_5734_7;

Selector_2 s5734_7(wires_1433_6[2], addr_1433_6, addr_positional[22939:22936], addr_5734_7);

wire[31:0] addr_5735_7;

Selector_2 s5735_7(wires_1433_6[3], addr_1433_6, addr_positional[22943:22940], addr_5735_7);

wire[31:0] addr_5736_7;

Selector_2 s5736_7(wires_1434_6[0], addr_1434_6, addr_positional[22947:22944], addr_5736_7);

wire[31:0] addr_5737_7;

Selector_2 s5737_7(wires_1434_6[1], addr_1434_6, addr_positional[22951:22948], addr_5737_7);

wire[31:0] addr_5738_7;

Selector_2 s5738_7(wires_1434_6[2], addr_1434_6, addr_positional[22955:22952], addr_5738_7);

wire[31:0] addr_5739_7;

Selector_2 s5739_7(wires_1434_6[3], addr_1434_6, addr_positional[22959:22956], addr_5739_7);

wire[31:0] addr_5740_7;

Selector_2 s5740_7(wires_1435_6[0], addr_1435_6, addr_positional[22963:22960], addr_5740_7);

wire[31:0] addr_5741_7;

Selector_2 s5741_7(wires_1435_6[1], addr_1435_6, addr_positional[22967:22964], addr_5741_7);

wire[31:0] addr_5742_7;

Selector_2 s5742_7(wires_1435_6[2], addr_1435_6, addr_positional[22971:22968], addr_5742_7);

wire[31:0] addr_5743_7;

Selector_2 s5743_7(wires_1435_6[3], addr_1435_6, addr_positional[22975:22972], addr_5743_7);

wire[31:0] addr_5744_7;

Selector_2 s5744_7(wires_1436_6[0], addr_1436_6, addr_positional[22979:22976], addr_5744_7);

wire[31:0] addr_5745_7;

Selector_2 s5745_7(wires_1436_6[1], addr_1436_6, addr_positional[22983:22980], addr_5745_7);

wire[31:0] addr_5746_7;

Selector_2 s5746_7(wires_1436_6[2], addr_1436_6, addr_positional[22987:22984], addr_5746_7);

wire[31:0] addr_5747_7;

Selector_2 s5747_7(wires_1436_6[3], addr_1436_6, addr_positional[22991:22988], addr_5747_7);

wire[31:0] addr_5748_7;

Selector_2 s5748_7(wires_1437_6[0], addr_1437_6, addr_positional[22995:22992], addr_5748_7);

wire[31:0] addr_5749_7;

Selector_2 s5749_7(wires_1437_6[1], addr_1437_6, addr_positional[22999:22996], addr_5749_7);

wire[31:0] addr_5750_7;

Selector_2 s5750_7(wires_1437_6[2], addr_1437_6, addr_positional[23003:23000], addr_5750_7);

wire[31:0] addr_5751_7;

Selector_2 s5751_7(wires_1437_6[3], addr_1437_6, addr_positional[23007:23004], addr_5751_7);

wire[31:0] addr_5752_7;

Selector_2 s5752_7(wires_1438_6[0], addr_1438_6, addr_positional[23011:23008], addr_5752_7);

wire[31:0] addr_5753_7;

Selector_2 s5753_7(wires_1438_6[1], addr_1438_6, addr_positional[23015:23012], addr_5753_7);

wire[31:0] addr_5754_7;

Selector_2 s5754_7(wires_1438_6[2], addr_1438_6, addr_positional[23019:23016], addr_5754_7);

wire[31:0] addr_5755_7;

Selector_2 s5755_7(wires_1438_6[3], addr_1438_6, addr_positional[23023:23020], addr_5755_7);

wire[31:0] addr_5756_7;

Selector_2 s5756_7(wires_1439_6[0], addr_1439_6, addr_positional[23027:23024], addr_5756_7);

wire[31:0] addr_5757_7;

Selector_2 s5757_7(wires_1439_6[1], addr_1439_6, addr_positional[23031:23028], addr_5757_7);

wire[31:0] addr_5758_7;

Selector_2 s5758_7(wires_1439_6[2], addr_1439_6, addr_positional[23035:23032], addr_5758_7);

wire[31:0] addr_5759_7;

Selector_2 s5759_7(wires_1439_6[3], addr_1439_6, addr_positional[23039:23036], addr_5759_7);

wire[31:0] addr_5760_7;

Selector_2 s5760_7(wires_1440_6[0], addr_1440_6, addr_positional[23043:23040], addr_5760_7);

wire[31:0] addr_5761_7;

Selector_2 s5761_7(wires_1440_6[1], addr_1440_6, addr_positional[23047:23044], addr_5761_7);

wire[31:0] addr_5762_7;

Selector_2 s5762_7(wires_1440_6[2], addr_1440_6, addr_positional[23051:23048], addr_5762_7);

wire[31:0] addr_5763_7;

Selector_2 s5763_7(wires_1440_6[3], addr_1440_6, addr_positional[23055:23052], addr_5763_7);

wire[31:0] addr_5764_7;

Selector_2 s5764_7(wires_1441_6[0], addr_1441_6, addr_positional[23059:23056], addr_5764_7);

wire[31:0] addr_5765_7;

Selector_2 s5765_7(wires_1441_6[1], addr_1441_6, addr_positional[23063:23060], addr_5765_7);

wire[31:0] addr_5766_7;

Selector_2 s5766_7(wires_1441_6[2], addr_1441_6, addr_positional[23067:23064], addr_5766_7);

wire[31:0] addr_5767_7;

Selector_2 s5767_7(wires_1441_6[3], addr_1441_6, addr_positional[23071:23068], addr_5767_7);

wire[31:0] addr_5768_7;

Selector_2 s5768_7(wires_1442_6[0], addr_1442_6, addr_positional[23075:23072], addr_5768_7);

wire[31:0] addr_5769_7;

Selector_2 s5769_7(wires_1442_6[1], addr_1442_6, addr_positional[23079:23076], addr_5769_7);

wire[31:0] addr_5770_7;

Selector_2 s5770_7(wires_1442_6[2], addr_1442_6, addr_positional[23083:23080], addr_5770_7);

wire[31:0] addr_5771_7;

Selector_2 s5771_7(wires_1442_6[3], addr_1442_6, addr_positional[23087:23084], addr_5771_7);

wire[31:0] addr_5772_7;

Selector_2 s5772_7(wires_1443_6[0], addr_1443_6, addr_positional[23091:23088], addr_5772_7);

wire[31:0] addr_5773_7;

Selector_2 s5773_7(wires_1443_6[1], addr_1443_6, addr_positional[23095:23092], addr_5773_7);

wire[31:0] addr_5774_7;

Selector_2 s5774_7(wires_1443_6[2], addr_1443_6, addr_positional[23099:23096], addr_5774_7);

wire[31:0] addr_5775_7;

Selector_2 s5775_7(wires_1443_6[3], addr_1443_6, addr_positional[23103:23100], addr_5775_7);

wire[31:0] addr_5776_7;

Selector_2 s5776_7(wires_1444_6[0], addr_1444_6, addr_positional[23107:23104], addr_5776_7);

wire[31:0] addr_5777_7;

Selector_2 s5777_7(wires_1444_6[1], addr_1444_6, addr_positional[23111:23108], addr_5777_7);

wire[31:0] addr_5778_7;

Selector_2 s5778_7(wires_1444_6[2], addr_1444_6, addr_positional[23115:23112], addr_5778_7);

wire[31:0] addr_5779_7;

Selector_2 s5779_7(wires_1444_6[3], addr_1444_6, addr_positional[23119:23116], addr_5779_7);

wire[31:0] addr_5780_7;

Selector_2 s5780_7(wires_1445_6[0], addr_1445_6, addr_positional[23123:23120], addr_5780_7);

wire[31:0] addr_5781_7;

Selector_2 s5781_7(wires_1445_6[1], addr_1445_6, addr_positional[23127:23124], addr_5781_7);

wire[31:0] addr_5782_7;

Selector_2 s5782_7(wires_1445_6[2], addr_1445_6, addr_positional[23131:23128], addr_5782_7);

wire[31:0] addr_5783_7;

Selector_2 s5783_7(wires_1445_6[3], addr_1445_6, addr_positional[23135:23132], addr_5783_7);

wire[31:0] addr_5784_7;

Selector_2 s5784_7(wires_1446_6[0], addr_1446_6, addr_positional[23139:23136], addr_5784_7);

wire[31:0] addr_5785_7;

Selector_2 s5785_7(wires_1446_6[1], addr_1446_6, addr_positional[23143:23140], addr_5785_7);

wire[31:0] addr_5786_7;

Selector_2 s5786_7(wires_1446_6[2], addr_1446_6, addr_positional[23147:23144], addr_5786_7);

wire[31:0] addr_5787_7;

Selector_2 s5787_7(wires_1446_6[3], addr_1446_6, addr_positional[23151:23148], addr_5787_7);

wire[31:0] addr_5788_7;

Selector_2 s5788_7(wires_1447_6[0], addr_1447_6, addr_positional[23155:23152], addr_5788_7);

wire[31:0] addr_5789_7;

Selector_2 s5789_7(wires_1447_6[1], addr_1447_6, addr_positional[23159:23156], addr_5789_7);

wire[31:0] addr_5790_7;

Selector_2 s5790_7(wires_1447_6[2], addr_1447_6, addr_positional[23163:23160], addr_5790_7);

wire[31:0] addr_5791_7;

Selector_2 s5791_7(wires_1447_6[3], addr_1447_6, addr_positional[23167:23164], addr_5791_7);

wire[31:0] addr_5792_7;

Selector_2 s5792_7(wires_1448_6[0], addr_1448_6, addr_positional[23171:23168], addr_5792_7);

wire[31:0] addr_5793_7;

Selector_2 s5793_7(wires_1448_6[1], addr_1448_6, addr_positional[23175:23172], addr_5793_7);

wire[31:0] addr_5794_7;

Selector_2 s5794_7(wires_1448_6[2], addr_1448_6, addr_positional[23179:23176], addr_5794_7);

wire[31:0] addr_5795_7;

Selector_2 s5795_7(wires_1448_6[3], addr_1448_6, addr_positional[23183:23180], addr_5795_7);

wire[31:0] addr_5796_7;

Selector_2 s5796_7(wires_1449_6[0], addr_1449_6, addr_positional[23187:23184], addr_5796_7);

wire[31:0] addr_5797_7;

Selector_2 s5797_7(wires_1449_6[1], addr_1449_6, addr_positional[23191:23188], addr_5797_7);

wire[31:0] addr_5798_7;

Selector_2 s5798_7(wires_1449_6[2], addr_1449_6, addr_positional[23195:23192], addr_5798_7);

wire[31:0] addr_5799_7;

Selector_2 s5799_7(wires_1449_6[3], addr_1449_6, addr_positional[23199:23196], addr_5799_7);

wire[31:0] addr_5800_7;

Selector_2 s5800_7(wires_1450_6[0], addr_1450_6, addr_positional[23203:23200], addr_5800_7);

wire[31:0] addr_5801_7;

Selector_2 s5801_7(wires_1450_6[1], addr_1450_6, addr_positional[23207:23204], addr_5801_7);

wire[31:0] addr_5802_7;

Selector_2 s5802_7(wires_1450_6[2], addr_1450_6, addr_positional[23211:23208], addr_5802_7);

wire[31:0] addr_5803_7;

Selector_2 s5803_7(wires_1450_6[3], addr_1450_6, addr_positional[23215:23212], addr_5803_7);

wire[31:0] addr_5804_7;

Selector_2 s5804_7(wires_1451_6[0], addr_1451_6, addr_positional[23219:23216], addr_5804_7);

wire[31:0] addr_5805_7;

Selector_2 s5805_7(wires_1451_6[1], addr_1451_6, addr_positional[23223:23220], addr_5805_7);

wire[31:0] addr_5806_7;

Selector_2 s5806_7(wires_1451_6[2], addr_1451_6, addr_positional[23227:23224], addr_5806_7);

wire[31:0] addr_5807_7;

Selector_2 s5807_7(wires_1451_6[3], addr_1451_6, addr_positional[23231:23228], addr_5807_7);

wire[31:0] addr_5808_7;

Selector_2 s5808_7(wires_1452_6[0], addr_1452_6, addr_positional[23235:23232], addr_5808_7);

wire[31:0] addr_5809_7;

Selector_2 s5809_7(wires_1452_6[1], addr_1452_6, addr_positional[23239:23236], addr_5809_7);

wire[31:0] addr_5810_7;

Selector_2 s5810_7(wires_1452_6[2], addr_1452_6, addr_positional[23243:23240], addr_5810_7);

wire[31:0] addr_5811_7;

Selector_2 s5811_7(wires_1452_6[3], addr_1452_6, addr_positional[23247:23244], addr_5811_7);

wire[31:0] addr_5812_7;

Selector_2 s5812_7(wires_1453_6[0], addr_1453_6, addr_positional[23251:23248], addr_5812_7);

wire[31:0] addr_5813_7;

Selector_2 s5813_7(wires_1453_6[1], addr_1453_6, addr_positional[23255:23252], addr_5813_7);

wire[31:0] addr_5814_7;

Selector_2 s5814_7(wires_1453_6[2], addr_1453_6, addr_positional[23259:23256], addr_5814_7);

wire[31:0] addr_5815_7;

Selector_2 s5815_7(wires_1453_6[3], addr_1453_6, addr_positional[23263:23260], addr_5815_7);

wire[31:0] addr_5816_7;

Selector_2 s5816_7(wires_1454_6[0], addr_1454_6, addr_positional[23267:23264], addr_5816_7);

wire[31:0] addr_5817_7;

Selector_2 s5817_7(wires_1454_6[1], addr_1454_6, addr_positional[23271:23268], addr_5817_7);

wire[31:0] addr_5818_7;

Selector_2 s5818_7(wires_1454_6[2], addr_1454_6, addr_positional[23275:23272], addr_5818_7);

wire[31:0] addr_5819_7;

Selector_2 s5819_7(wires_1454_6[3], addr_1454_6, addr_positional[23279:23276], addr_5819_7);

wire[31:0] addr_5820_7;

Selector_2 s5820_7(wires_1455_6[0], addr_1455_6, addr_positional[23283:23280], addr_5820_7);

wire[31:0] addr_5821_7;

Selector_2 s5821_7(wires_1455_6[1], addr_1455_6, addr_positional[23287:23284], addr_5821_7);

wire[31:0] addr_5822_7;

Selector_2 s5822_7(wires_1455_6[2], addr_1455_6, addr_positional[23291:23288], addr_5822_7);

wire[31:0] addr_5823_7;

Selector_2 s5823_7(wires_1455_6[3], addr_1455_6, addr_positional[23295:23292], addr_5823_7);

wire[31:0] addr_5824_7;

Selector_2 s5824_7(wires_1456_6[0], addr_1456_6, addr_positional[23299:23296], addr_5824_7);

wire[31:0] addr_5825_7;

Selector_2 s5825_7(wires_1456_6[1], addr_1456_6, addr_positional[23303:23300], addr_5825_7);

wire[31:0] addr_5826_7;

Selector_2 s5826_7(wires_1456_6[2], addr_1456_6, addr_positional[23307:23304], addr_5826_7);

wire[31:0] addr_5827_7;

Selector_2 s5827_7(wires_1456_6[3], addr_1456_6, addr_positional[23311:23308], addr_5827_7);

wire[31:0] addr_5828_7;

Selector_2 s5828_7(wires_1457_6[0], addr_1457_6, addr_positional[23315:23312], addr_5828_7);

wire[31:0] addr_5829_7;

Selector_2 s5829_7(wires_1457_6[1], addr_1457_6, addr_positional[23319:23316], addr_5829_7);

wire[31:0] addr_5830_7;

Selector_2 s5830_7(wires_1457_6[2], addr_1457_6, addr_positional[23323:23320], addr_5830_7);

wire[31:0] addr_5831_7;

Selector_2 s5831_7(wires_1457_6[3], addr_1457_6, addr_positional[23327:23324], addr_5831_7);

wire[31:0] addr_5832_7;

Selector_2 s5832_7(wires_1458_6[0], addr_1458_6, addr_positional[23331:23328], addr_5832_7);

wire[31:0] addr_5833_7;

Selector_2 s5833_7(wires_1458_6[1], addr_1458_6, addr_positional[23335:23332], addr_5833_7);

wire[31:0] addr_5834_7;

Selector_2 s5834_7(wires_1458_6[2], addr_1458_6, addr_positional[23339:23336], addr_5834_7);

wire[31:0] addr_5835_7;

Selector_2 s5835_7(wires_1458_6[3], addr_1458_6, addr_positional[23343:23340], addr_5835_7);

wire[31:0] addr_5836_7;

Selector_2 s5836_7(wires_1459_6[0], addr_1459_6, addr_positional[23347:23344], addr_5836_7);

wire[31:0] addr_5837_7;

Selector_2 s5837_7(wires_1459_6[1], addr_1459_6, addr_positional[23351:23348], addr_5837_7);

wire[31:0] addr_5838_7;

Selector_2 s5838_7(wires_1459_6[2], addr_1459_6, addr_positional[23355:23352], addr_5838_7);

wire[31:0] addr_5839_7;

Selector_2 s5839_7(wires_1459_6[3], addr_1459_6, addr_positional[23359:23356], addr_5839_7);

wire[31:0] addr_5840_7;

Selector_2 s5840_7(wires_1460_6[0], addr_1460_6, addr_positional[23363:23360], addr_5840_7);

wire[31:0] addr_5841_7;

Selector_2 s5841_7(wires_1460_6[1], addr_1460_6, addr_positional[23367:23364], addr_5841_7);

wire[31:0] addr_5842_7;

Selector_2 s5842_7(wires_1460_6[2], addr_1460_6, addr_positional[23371:23368], addr_5842_7);

wire[31:0] addr_5843_7;

Selector_2 s5843_7(wires_1460_6[3], addr_1460_6, addr_positional[23375:23372], addr_5843_7);

wire[31:0] addr_5844_7;

Selector_2 s5844_7(wires_1461_6[0], addr_1461_6, addr_positional[23379:23376], addr_5844_7);

wire[31:0] addr_5845_7;

Selector_2 s5845_7(wires_1461_6[1], addr_1461_6, addr_positional[23383:23380], addr_5845_7);

wire[31:0] addr_5846_7;

Selector_2 s5846_7(wires_1461_6[2], addr_1461_6, addr_positional[23387:23384], addr_5846_7);

wire[31:0] addr_5847_7;

Selector_2 s5847_7(wires_1461_6[3], addr_1461_6, addr_positional[23391:23388], addr_5847_7);

wire[31:0] addr_5848_7;

Selector_2 s5848_7(wires_1462_6[0], addr_1462_6, addr_positional[23395:23392], addr_5848_7);

wire[31:0] addr_5849_7;

Selector_2 s5849_7(wires_1462_6[1], addr_1462_6, addr_positional[23399:23396], addr_5849_7);

wire[31:0] addr_5850_7;

Selector_2 s5850_7(wires_1462_6[2], addr_1462_6, addr_positional[23403:23400], addr_5850_7);

wire[31:0] addr_5851_7;

Selector_2 s5851_7(wires_1462_6[3], addr_1462_6, addr_positional[23407:23404], addr_5851_7);

wire[31:0] addr_5852_7;

Selector_2 s5852_7(wires_1463_6[0], addr_1463_6, addr_positional[23411:23408], addr_5852_7);

wire[31:0] addr_5853_7;

Selector_2 s5853_7(wires_1463_6[1], addr_1463_6, addr_positional[23415:23412], addr_5853_7);

wire[31:0] addr_5854_7;

Selector_2 s5854_7(wires_1463_6[2], addr_1463_6, addr_positional[23419:23416], addr_5854_7);

wire[31:0] addr_5855_7;

Selector_2 s5855_7(wires_1463_6[3], addr_1463_6, addr_positional[23423:23420], addr_5855_7);

wire[31:0] addr_5856_7;

Selector_2 s5856_7(wires_1464_6[0], addr_1464_6, addr_positional[23427:23424], addr_5856_7);

wire[31:0] addr_5857_7;

Selector_2 s5857_7(wires_1464_6[1], addr_1464_6, addr_positional[23431:23428], addr_5857_7);

wire[31:0] addr_5858_7;

Selector_2 s5858_7(wires_1464_6[2], addr_1464_6, addr_positional[23435:23432], addr_5858_7);

wire[31:0] addr_5859_7;

Selector_2 s5859_7(wires_1464_6[3], addr_1464_6, addr_positional[23439:23436], addr_5859_7);

wire[31:0] addr_5860_7;

Selector_2 s5860_7(wires_1465_6[0], addr_1465_6, addr_positional[23443:23440], addr_5860_7);

wire[31:0] addr_5861_7;

Selector_2 s5861_7(wires_1465_6[1], addr_1465_6, addr_positional[23447:23444], addr_5861_7);

wire[31:0] addr_5862_7;

Selector_2 s5862_7(wires_1465_6[2], addr_1465_6, addr_positional[23451:23448], addr_5862_7);

wire[31:0] addr_5863_7;

Selector_2 s5863_7(wires_1465_6[3], addr_1465_6, addr_positional[23455:23452], addr_5863_7);

wire[31:0] addr_5864_7;

Selector_2 s5864_7(wires_1466_6[0], addr_1466_6, addr_positional[23459:23456], addr_5864_7);

wire[31:0] addr_5865_7;

Selector_2 s5865_7(wires_1466_6[1], addr_1466_6, addr_positional[23463:23460], addr_5865_7);

wire[31:0] addr_5866_7;

Selector_2 s5866_7(wires_1466_6[2], addr_1466_6, addr_positional[23467:23464], addr_5866_7);

wire[31:0] addr_5867_7;

Selector_2 s5867_7(wires_1466_6[3], addr_1466_6, addr_positional[23471:23468], addr_5867_7);

wire[31:0] addr_5868_7;

Selector_2 s5868_7(wires_1467_6[0], addr_1467_6, addr_positional[23475:23472], addr_5868_7);

wire[31:0] addr_5869_7;

Selector_2 s5869_7(wires_1467_6[1], addr_1467_6, addr_positional[23479:23476], addr_5869_7);

wire[31:0] addr_5870_7;

Selector_2 s5870_7(wires_1467_6[2], addr_1467_6, addr_positional[23483:23480], addr_5870_7);

wire[31:0] addr_5871_7;

Selector_2 s5871_7(wires_1467_6[3], addr_1467_6, addr_positional[23487:23484], addr_5871_7);

wire[31:0] addr_5872_7;

Selector_2 s5872_7(wires_1468_6[0], addr_1468_6, addr_positional[23491:23488], addr_5872_7);

wire[31:0] addr_5873_7;

Selector_2 s5873_7(wires_1468_6[1], addr_1468_6, addr_positional[23495:23492], addr_5873_7);

wire[31:0] addr_5874_7;

Selector_2 s5874_7(wires_1468_6[2], addr_1468_6, addr_positional[23499:23496], addr_5874_7);

wire[31:0] addr_5875_7;

Selector_2 s5875_7(wires_1468_6[3], addr_1468_6, addr_positional[23503:23500], addr_5875_7);

wire[31:0] addr_5876_7;

Selector_2 s5876_7(wires_1469_6[0], addr_1469_6, addr_positional[23507:23504], addr_5876_7);

wire[31:0] addr_5877_7;

Selector_2 s5877_7(wires_1469_6[1], addr_1469_6, addr_positional[23511:23508], addr_5877_7);

wire[31:0] addr_5878_7;

Selector_2 s5878_7(wires_1469_6[2], addr_1469_6, addr_positional[23515:23512], addr_5878_7);

wire[31:0] addr_5879_7;

Selector_2 s5879_7(wires_1469_6[3], addr_1469_6, addr_positional[23519:23516], addr_5879_7);

wire[31:0] addr_5880_7;

Selector_2 s5880_7(wires_1470_6[0], addr_1470_6, addr_positional[23523:23520], addr_5880_7);

wire[31:0] addr_5881_7;

Selector_2 s5881_7(wires_1470_6[1], addr_1470_6, addr_positional[23527:23524], addr_5881_7);

wire[31:0] addr_5882_7;

Selector_2 s5882_7(wires_1470_6[2], addr_1470_6, addr_positional[23531:23528], addr_5882_7);

wire[31:0] addr_5883_7;

Selector_2 s5883_7(wires_1470_6[3], addr_1470_6, addr_positional[23535:23532], addr_5883_7);

wire[31:0] addr_5884_7;

Selector_2 s5884_7(wires_1471_6[0], addr_1471_6, addr_positional[23539:23536], addr_5884_7);

wire[31:0] addr_5885_7;

Selector_2 s5885_7(wires_1471_6[1], addr_1471_6, addr_positional[23543:23540], addr_5885_7);

wire[31:0] addr_5886_7;

Selector_2 s5886_7(wires_1471_6[2], addr_1471_6, addr_positional[23547:23544], addr_5886_7);

wire[31:0] addr_5887_7;

Selector_2 s5887_7(wires_1471_6[3], addr_1471_6, addr_positional[23551:23548], addr_5887_7);

wire[31:0] addr_5888_7;

Selector_2 s5888_7(wires_1472_6[0], addr_1472_6, addr_positional[23555:23552], addr_5888_7);

wire[31:0] addr_5889_7;

Selector_2 s5889_7(wires_1472_6[1], addr_1472_6, addr_positional[23559:23556], addr_5889_7);

wire[31:0] addr_5890_7;

Selector_2 s5890_7(wires_1472_6[2], addr_1472_6, addr_positional[23563:23560], addr_5890_7);

wire[31:0] addr_5891_7;

Selector_2 s5891_7(wires_1472_6[3], addr_1472_6, addr_positional[23567:23564], addr_5891_7);

wire[31:0] addr_5892_7;

Selector_2 s5892_7(wires_1473_6[0], addr_1473_6, addr_positional[23571:23568], addr_5892_7);

wire[31:0] addr_5893_7;

Selector_2 s5893_7(wires_1473_6[1], addr_1473_6, addr_positional[23575:23572], addr_5893_7);

wire[31:0] addr_5894_7;

Selector_2 s5894_7(wires_1473_6[2], addr_1473_6, addr_positional[23579:23576], addr_5894_7);

wire[31:0] addr_5895_7;

Selector_2 s5895_7(wires_1473_6[3], addr_1473_6, addr_positional[23583:23580], addr_5895_7);

wire[31:0] addr_5896_7;

Selector_2 s5896_7(wires_1474_6[0], addr_1474_6, addr_positional[23587:23584], addr_5896_7);

wire[31:0] addr_5897_7;

Selector_2 s5897_7(wires_1474_6[1], addr_1474_6, addr_positional[23591:23588], addr_5897_7);

wire[31:0] addr_5898_7;

Selector_2 s5898_7(wires_1474_6[2], addr_1474_6, addr_positional[23595:23592], addr_5898_7);

wire[31:0] addr_5899_7;

Selector_2 s5899_7(wires_1474_6[3], addr_1474_6, addr_positional[23599:23596], addr_5899_7);

wire[31:0] addr_5900_7;

Selector_2 s5900_7(wires_1475_6[0], addr_1475_6, addr_positional[23603:23600], addr_5900_7);

wire[31:0] addr_5901_7;

Selector_2 s5901_7(wires_1475_6[1], addr_1475_6, addr_positional[23607:23604], addr_5901_7);

wire[31:0] addr_5902_7;

Selector_2 s5902_7(wires_1475_6[2], addr_1475_6, addr_positional[23611:23608], addr_5902_7);

wire[31:0] addr_5903_7;

Selector_2 s5903_7(wires_1475_6[3], addr_1475_6, addr_positional[23615:23612], addr_5903_7);

wire[31:0] addr_5904_7;

Selector_2 s5904_7(wires_1476_6[0], addr_1476_6, addr_positional[23619:23616], addr_5904_7);

wire[31:0] addr_5905_7;

Selector_2 s5905_7(wires_1476_6[1], addr_1476_6, addr_positional[23623:23620], addr_5905_7);

wire[31:0] addr_5906_7;

Selector_2 s5906_7(wires_1476_6[2], addr_1476_6, addr_positional[23627:23624], addr_5906_7);

wire[31:0] addr_5907_7;

Selector_2 s5907_7(wires_1476_6[3], addr_1476_6, addr_positional[23631:23628], addr_5907_7);

wire[31:0] addr_5908_7;

Selector_2 s5908_7(wires_1477_6[0], addr_1477_6, addr_positional[23635:23632], addr_5908_7);

wire[31:0] addr_5909_7;

Selector_2 s5909_7(wires_1477_6[1], addr_1477_6, addr_positional[23639:23636], addr_5909_7);

wire[31:0] addr_5910_7;

Selector_2 s5910_7(wires_1477_6[2], addr_1477_6, addr_positional[23643:23640], addr_5910_7);

wire[31:0] addr_5911_7;

Selector_2 s5911_7(wires_1477_6[3], addr_1477_6, addr_positional[23647:23644], addr_5911_7);

wire[31:0] addr_5912_7;

Selector_2 s5912_7(wires_1478_6[0], addr_1478_6, addr_positional[23651:23648], addr_5912_7);

wire[31:0] addr_5913_7;

Selector_2 s5913_7(wires_1478_6[1], addr_1478_6, addr_positional[23655:23652], addr_5913_7);

wire[31:0] addr_5914_7;

Selector_2 s5914_7(wires_1478_6[2], addr_1478_6, addr_positional[23659:23656], addr_5914_7);

wire[31:0] addr_5915_7;

Selector_2 s5915_7(wires_1478_6[3], addr_1478_6, addr_positional[23663:23660], addr_5915_7);

wire[31:0] addr_5916_7;

Selector_2 s5916_7(wires_1479_6[0], addr_1479_6, addr_positional[23667:23664], addr_5916_7);

wire[31:0] addr_5917_7;

Selector_2 s5917_7(wires_1479_6[1], addr_1479_6, addr_positional[23671:23668], addr_5917_7);

wire[31:0] addr_5918_7;

Selector_2 s5918_7(wires_1479_6[2], addr_1479_6, addr_positional[23675:23672], addr_5918_7);

wire[31:0] addr_5919_7;

Selector_2 s5919_7(wires_1479_6[3], addr_1479_6, addr_positional[23679:23676], addr_5919_7);

wire[31:0] addr_5920_7;

Selector_2 s5920_7(wires_1480_6[0], addr_1480_6, addr_positional[23683:23680], addr_5920_7);

wire[31:0] addr_5921_7;

Selector_2 s5921_7(wires_1480_6[1], addr_1480_6, addr_positional[23687:23684], addr_5921_7);

wire[31:0] addr_5922_7;

Selector_2 s5922_7(wires_1480_6[2], addr_1480_6, addr_positional[23691:23688], addr_5922_7);

wire[31:0] addr_5923_7;

Selector_2 s5923_7(wires_1480_6[3], addr_1480_6, addr_positional[23695:23692], addr_5923_7);

wire[31:0] addr_5924_7;

Selector_2 s5924_7(wires_1481_6[0], addr_1481_6, addr_positional[23699:23696], addr_5924_7);

wire[31:0] addr_5925_7;

Selector_2 s5925_7(wires_1481_6[1], addr_1481_6, addr_positional[23703:23700], addr_5925_7);

wire[31:0] addr_5926_7;

Selector_2 s5926_7(wires_1481_6[2], addr_1481_6, addr_positional[23707:23704], addr_5926_7);

wire[31:0] addr_5927_7;

Selector_2 s5927_7(wires_1481_6[3], addr_1481_6, addr_positional[23711:23708], addr_5927_7);

wire[31:0] addr_5928_7;

Selector_2 s5928_7(wires_1482_6[0], addr_1482_6, addr_positional[23715:23712], addr_5928_7);

wire[31:0] addr_5929_7;

Selector_2 s5929_7(wires_1482_6[1], addr_1482_6, addr_positional[23719:23716], addr_5929_7);

wire[31:0] addr_5930_7;

Selector_2 s5930_7(wires_1482_6[2], addr_1482_6, addr_positional[23723:23720], addr_5930_7);

wire[31:0] addr_5931_7;

Selector_2 s5931_7(wires_1482_6[3], addr_1482_6, addr_positional[23727:23724], addr_5931_7);

wire[31:0] addr_5932_7;

Selector_2 s5932_7(wires_1483_6[0], addr_1483_6, addr_positional[23731:23728], addr_5932_7);

wire[31:0] addr_5933_7;

Selector_2 s5933_7(wires_1483_6[1], addr_1483_6, addr_positional[23735:23732], addr_5933_7);

wire[31:0] addr_5934_7;

Selector_2 s5934_7(wires_1483_6[2], addr_1483_6, addr_positional[23739:23736], addr_5934_7);

wire[31:0] addr_5935_7;

Selector_2 s5935_7(wires_1483_6[3], addr_1483_6, addr_positional[23743:23740], addr_5935_7);

wire[31:0] addr_5936_7;

Selector_2 s5936_7(wires_1484_6[0], addr_1484_6, addr_positional[23747:23744], addr_5936_7);

wire[31:0] addr_5937_7;

Selector_2 s5937_7(wires_1484_6[1], addr_1484_6, addr_positional[23751:23748], addr_5937_7);

wire[31:0] addr_5938_7;

Selector_2 s5938_7(wires_1484_6[2], addr_1484_6, addr_positional[23755:23752], addr_5938_7);

wire[31:0] addr_5939_7;

Selector_2 s5939_7(wires_1484_6[3], addr_1484_6, addr_positional[23759:23756], addr_5939_7);

wire[31:0] addr_5940_7;

Selector_2 s5940_7(wires_1485_6[0], addr_1485_6, addr_positional[23763:23760], addr_5940_7);

wire[31:0] addr_5941_7;

Selector_2 s5941_7(wires_1485_6[1], addr_1485_6, addr_positional[23767:23764], addr_5941_7);

wire[31:0] addr_5942_7;

Selector_2 s5942_7(wires_1485_6[2], addr_1485_6, addr_positional[23771:23768], addr_5942_7);

wire[31:0] addr_5943_7;

Selector_2 s5943_7(wires_1485_6[3], addr_1485_6, addr_positional[23775:23772], addr_5943_7);

wire[31:0] addr_5944_7;

Selector_2 s5944_7(wires_1486_6[0], addr_1486_6, addr_positional[23779:23776], addr_5944_7);

wire[31:0] addr_5945_7;

Selector_2 s5945_7(wires_1486_6[1], addr_1486_6, addr_positional[23783:23780], addr_5945_7);

wire[31:0] addr_5946_7;

Selector_2 s5946_7(wires_1486_6[2], addr_1486_6, addr_positional[23787:23784], addr_5946_7);

wire[31:0] addr_5947_7;

Selector_2 s5947_7(wires_1486_6[3], addr_1486_6, addr_positional[23791:23788], addr_5947_7);

wire[31:0] addr_5948_7;

Selector_2 s5948_7(wires_1487_6[0], addr_1487_6, addr_positional[23795:23792], addr_5948_7);

wire[31:0] addr_5949_7;

Selector_2 s5949_7(wires_1487_6[1], addr_1487_6, addr_positional[23799:23796], addr_5949_7);

wire[31:0] addr_5950_7;

Selector_2 s5950_7(wires_1487_6[2], addr_1487_6, addr_positional[23803:23800], addr_5950_7);

wire[31:0] addr_5951_7;

Selector_2 s5951_7(wires_1487_6[3], addr_1487_6, addr_positional[23807:23804], addr_5951_7);

wire[31:0] addr_5952_7;

Selector_2 s5952_7(wires_1488_6[0], addr_1488_6, addr_positional[23811:23808], addr_5952_7);

wire[31:0] addr_5953_7;

Selector_2 s5953_7(wires_1488_6[1], addr_1488_6, addr_positional[23815:23812], addr_5953_7);

wire[31:0] addr_5954_7;

Selector_2 s5954_7(wires_1488_6[2], addr_1488_6, addr_positional[23819:23816], addr_5954_7);

wire[31:0] addr_5955_7;

Selector_2 s5955_7(wires_1488_6[3], addr_1488_6, addr_positional[23823:23820], addr_5955_7);

wire[31:0] addr_5956_7;

Selector_2 s5956_7(wires_1489_6[0], addr_1489_6, addr_positional[23827:23824], addr_5956_7);

wire[31:0] addr_5957_7;

Selector_2 s5957_7(wires_1489_6[1], addr_1489_6, addr_positional[23831:23828], addr_5957_7);

wire[31:0] addr_5958_7;

Selector_2 s5958_7(wires_1489_6[2], addr_1489_6, addr_positional[23835:23832], addr_5958_7);

wire[31:0] addr_5959_7;

Selector_2 s5959_7(wires_1489_6[3], addr_1489_6, addr_positional[23839:23836], addr_5959_7);

wire[31:0] addr_5960_7;

Selector_2 s5960_7(wires_1490_6[0], addr_1490_6, addr_positional[23843:23840], addr_5960_7);

wire[31:0] addr_5961_7;

Selector_2 s5961_7(wires_1490_6[1], addr_1490_6, addr_positional[23847:23844], addr_5961_7);

wire[31:0] addr_5962_7;

Selector_2 s5962_7(wires_1490_6[2], addr_1490_6, addr_positional[23851:23848], addr_5962_7);

wire[31:0] addr_5963_7;

Selector_2 s5963_7(wires_1490_6[3], addr_1490_6, addr_positional[23855:23852], addr_5963_7);

wire[31:0] addr_5964_7;

Selector_2 s5964_7(wires_1491_6[0], addr_1491_6, addr_positional[23859:23856], addr_5964_7);

wire[31:0] addr_5965_7;

Selector_2 s5965_7(wires_1491_6[1], addr_1491_6, addr_positional[23863:23860], addr_5965_7);

wire[31:0] addr_5966_7;

Selector_2 s5966_7(wires_1491_6[2], addr_1491_6, addr_positional[23867:23864], addr_5966_7);

wire[31:0] addr_5967_7;

Selector_2 s5967_7(wires_1491_6[3], addr_1491_6, addr_positional[23871:23868], addr_5967_7);

wire[31:0] addr_5968_7;

Selector_2 s5968_7(wires_1492_6[0], addr_1492_6, addr_positional[23875:23872], addr_5968_7);

wire[31:0] addr_5969_7;

Selector_2 s5969_7(wires_1492_6[1], addr_1492_6, addr_positional[23879:23876], addr_5969_7);

wire[31:0] addr_5970_7;

Selector_2 s5970_7(wires_1492_6[2], addr_1492_6, addr_positional[23883:23880], addr_5970_7);

wire[31:0] addr_5971_7;

Selector_2 s5971_7(wires_1492_6[3], addr_1492_6, addr_positional[23887:23884], addr_5971_7);

wire[31:0] addr_5972_7;

Selector_2 s5972_7(wires_1493_6[0], addr_1493_6, addr_positional[23891:23888], addr_5972_7);

wire[31:0] addr_5973_7;

Selector_2 s5973_7(wires_1493_6[1], addr_1493_6, addr_positional[23895:23892], addr_5973_7);

wire[31:0] addr_5974_7;

Selector_2 s5974_7(wires_1493_6[2], addr_1493_6, addr_positional[23899:23896], addr_5974_7);

wire[31:0] addr_5975_7;

Selector_2 s5975_7(wires_1493_6[3], addr_1493_6, addr_positional[23903:23900], addr_5975_7);

wire[31:0] addr_5976_7;

Selector_2 s5976_7(wires_1494_6[0], addr_1494_6, addr_positional[23907:23904], addr_5976_7);

wire[31:0] addr_5977_7;

Selector_2 s5977_7(wires_1494_6[1], addr_1494_6, addr_positional[23911:23908], addr_5977_7);

wire[31:0] addr_5978_7;

Selector_2 s5978_7(wires_1494_6[2], addr_1494_6, addr_positional[23915:23912], addr_5978_7);

wire[31:0] addr_5979_7;

Selector_2 s5979_7(wires_1494_6[3], addr_1494_6, addr_positional[23919:23916], addr_5979_7);

wire[31:0] addr_5980_7;

Selector_2 s5980_7(wires_1495_6[0], addr_1495_6, addr_positional[23923:23920], addr_5980_7);

wire[31:0] addr_5981_7;

Selector_2 s5981_7(wires_1495_6[1], addr_1495_6, addr_positional[23927:23924], addr_5981_7);

wire[31:0] addr_5982_7;

Selector_2 s5982_7(wires_1495_6[2], addr_1495_6, addr_positional[23931:23928], addr_5982_7);

wire[31:0] addr_5983_7;

Selector_2 s5983_7(wires_1495_6[3], addr_1495_6, addr_positional[23935:23932], addr_5983_7);

wire[31:0] addr_5984_7;

Selector_2 s5984_7(wires_1496_6[0], addr_1496_6, addr_positional[23939:23936], addr_5984_7);

wire[31:0] addr_5985_7;

Selector_2 s5985_7(wires_1496_6[1], addr_1496_6, addr_positional[23943:23940], addr_5985_7);

wire[31:0] addr_5986_7;

Selector_2 s5986_7(wires_1496_6[2], addr_1496_6, addr_positional[23947:23944], addr_5986_7);

wire[31:0] addr_5987_7;

Selector_2 s5987_7(wires_1496_6[3], addr_1496_6, addr_positional[23951:23948], addr_5987_7);

wire[31:0] addr_5988_7;

Selector_2 s5988_7(wires_1497_6[0], addr_1497_6, addr_positional[23955:23952], addr_5988_7);

wire[31:0] addr_5989_7;

Selector_2 s5989_7(wires_1497_6[1], addr_1497_6, addr_positional[23959:23956], addr_5989_7);

wire[31:0] addr_5990_7;

Selector_2 s5990_7(wires_1497_6[2], addr_1497_6, addr_positional[23963:23960], addr_5990_7);

wire[31:0] addr_5991_7;

Selector_2 s5991_7(wires_1497_6[3], addr_1497_6, addr_positional[23967:23964], addr_5991_7);

wire[31:0] addr_5992_7;

Selector_2 s5992_7(wires_1498_6[0], addr_1498_6, addr_positional[23971:23968], addr_5992_7);

wire[31:0] addr_5993_7;

Selector_2 s5993_7(wires_1498_6[1], addr_1498_6, addr_positional[23975:23972], addr_5993_7);

wire[31:0] addr_5994_7;

Selector_2 s5994_7(wires_1498_6[2], addr_1498_6, addr_positional[23979:23976], addr_5994_7);

wire[31:0] addr_5995_7;

Selector_2 s5995_7(wires_1498_6[3], addr_1498_6, addr_positional[23983:23980], addr_5995_7);

wire[31:0] addr_5996_7;

Selector_2 s5996_7(wires_1499_6[0], addr_1499_6, addr_positional[23987:23984], addr_5996_7);

wire[31:0] addr_5997_7;

Selector_2 s5997_7(wires_1499_6[1], addr_1499_6, addr_positional[23991:23988], addr_5997_7);

wire[31:0] addr_5998_7;

Selector_2 s5998_7(wires_1499_6[2], addr_1499_6, addr_positional[23995:23992], addr_5998_7);

wire[31:0] addr_5999_7;

Selector_2 s5999_7(wires_1499_6[3], addr_1499_6, addr_positional[23999:23996], addr_5999_7);

wire[31:0] addr_6000_7;

Selector_2 s6000_7(wires_1500_6[0], addr_1500_6, addr_positional[24003:24000], addr_6000_7);

wire[31:0] addr_6001_7;

Selector_2 s6001_7(wires_1500_6[1], addr_1500_6, addr_positional[24007:24004], addr_6001_7);

wire[31:0] addr_6002_7;

Selector_2 s6002_7(wires_1500_6[2], addr_1500_6, addr_positional[24011:24008], addr_6002_7);

wire[31:0] addr_6003_7;

Selector_2 s6003_7(wires_1500_6[3], addr_1500_6, addr_positional[24015:24012], addr_6003_7);

wire[31:0] addr_6004_7;

Selector_2 s6004_7(wires_1501_6[0], addr_1501_6, addr_positional[24019:24016], addr_6004_7);

wire[31:0] addr_6005_7;

Selector_2 s6005_7(wires_1501_6[1], addr_1501_6, addr_positional[24023:24020], addr_6005_7);

wire[31:0] addr_6006_7;

Selector_2 s6006_7(wires_1501_6[2], addr_1501_6, addr_positional[24027:24024], addr_6006_7);

wire[31:0] addr_6007_7;

Selector_2 s6007_7(wires_1501_6[3], addr_1501_6, addr_positional[24031:24028], addr_6007_7);

wire[31:0] addr_6008_7;

Selector_2 s6008_7(wires_1502_6[0], addr_1502_6, addr_positional[24035:24032], addr_6008_7);

wire[31:0] addr_6009_7;

Selector_2 s6009_7(wires_1502_6[1], addr_1502_6, addr_positional[24039:24036], addr_6009_7);

wire[31:0] addr_6010_7;

Selector_2 s6010_7(wires_1502_6[2], addr_1502_6, addr_positional[24043:24040], addr_6010_7);

wire[31:0] addr_6011_7;

Selector_2 s6011_7(wires_1502_6[3], addr_1502_6, addr_positional[24047:24044], addr_6011_7);

wire[31:0] addr_6012_7;

Selector_2 s6012_7(wires_1503_6[0], addr_1503_6, addr_positional[24051:24048], addr_6012_7);

wire[31:0] addr_6013_7;

Selector_2 s6013_7(wires_1503_6[1], addr_1503_6, addr_positional[24055:24052], addr_6013_7);

wire[31:0] addr_6014_7;

Selector_2 s6014_7(wires_1503_6[2], addr_1503_6, addr_positional[24059:24056], addr_6014_7);

wire[31:0] addr_6015_7;

Selector_2 s6015_7(wires_1503_6[3], addr_1503_6, addr_positional[24063:24060], addr_6015_7);

wire[31:0] addr_6016_7;

Selector_2 s6016_7(wires_1504_6[0], addr_1504_6, addr_positional[24067:24064], addr_6016_7);

wire[31:0] addr_6017_7;

Selector_2 s6017_7(wires_1504_6[1], addr_1504_6, addr_positional[24071:24068], addr_6017_7);

wire[31:0] addr_6018_7;

Selector_2 s6018_7(wires_1504_6[2], addr_1504_6, addr_positional[24075:24072], addr_6018_7);

wire[31:0] addr_6019_7;

Selector_2 s6019_7(wires_1504_6[3], addr_1504_6, addr_positional[24079:24076], addr_6019_7);

wire[31:0] addr_6020_7;

Selector_2 s6020_7(wires_1505_6[0], addr_1505_6, addr_positional[24083:24080], addr_6020_7);

wire[31:0] addr_6021_7;

Selector_2 s6021_7(wires_1505_6[1], addr_1505_6, addr_positional[24087:24084], addr_6021_7);

wire[31:0] addr_6022_7;

Selector_2 s6022_7(wires_1505_6[2], addr_1505_6, addr_positional[24091:24088], addr_6022_7);

wire[31:0] addr_6023_7;

Selector_2 s6023_7(wires_1505_6[3], addr_1505_6, addr_positional[24095:24092], addr_6023_7);

wire[31:0] addr_6024_7;

Selector_2 s6024_7(wires_1506_6[0], addr_1506_6, addr_positional[24099:24096], addr_6024_7);

wire[31:0] addr_6025_7;

Selector_2 s6025_7(wires_1506_6[1], addr_1506_6, addr_positional[24103:24100], addr_6025_7);

wire[31:0] addr_6026_7;

Selector_2 s6026_7(wires_1506_6[2], addr_1506_6, addr_positional[24107:24104], addr_6026_7);

wire[31:0] addr_6027_7;

Selector_2 s6027_7(wires_1506_6[3], addr_1506_6, addr_positional[24111:24108], addr_6027_7);

wire[31:0] addr_6028_7;

Selector_2 s6028_7(wires_1507_6[0], addr_1507_6, addr_positional[24115:24112], addr_6028_7);

wire[31:0] addr_6029_7;

Selector_2 s6029_7(wires_1507_6[1], addr_1507_6, addr_positional[24119:24116], addr_6029_7);

wire[31:0] addr_6030_7;

Selector_2 s6030_7(wires_1507_6[2], addr_1507_6, addr_positional[24123:24120], addr_6030_7);

wire[31:0] addr_6031_7;

Selector_2 s6031_7(wires_1507_6[3], addr_1507_6, addr_positional[24127:24124], addr_6031_7);

wire[31:0] addr_6032_7;

Selector_2 s6032_7(wires_1508_6[0], addr_1508_6, addr_positional[24131:24128], addr_6032_7);

wire[31:0] addr_6033_7;

Selector_2 s6033_7(wires_1508_6[1], addr_1508_6, addr_positional[24135:24132], addr_6033_7);

wire[31:0] addr_6034_7;

Selector_2 s6034_7(wires_1508_6[2], addr_1508_6, addr_positional[24139:24136], addr_6034_7);

wire[31:0] addr_6035_7;

Selector_2 s6035_7(wires_1508_6[3], addr_1508_6, addr_positional[24143:24140], addr_6035_7);

wire[31:0] addr_6036_7;

Selector_2 s6036_7(wires_1509_6[0], addr_1509_6, addr_positional[24147:24144], addr_6036_7);

wire[31:0] addr_6037_7;

Selector_2 s6037_7(wires_1509_6[1], addr_1509_6, addr_positional[24151:24148], addr_6037_7);

wire[31:0] addr_6038_7;

Selector_2 s6038_7(wires_1509_6[2], addr_1509_6, addr_positional[24155:24152], addr_6038_7);

wire[31:0] addr_6039_7;

Selector_2 s6039_7(wires_1509_6[3], addr_1509_6, addr_positional[24159:24156], addr_6039_7);

wire[31:0] addr_6040_7;

Selector_2 s6040_7(wires_1510_6[0], addr_1510_6, addr_positional[24163:24160], addr_6040_7);

wire[31:0] addr_6041_7;

Selector_2 s6041_7(wires_1510_6[1], addr_1510_6, addr_positional[24167:24164], addr_6041_7);

wire[31:0] addr_6042_7;

Selector_2 s6042_7(wires_1510_6[2], addr_1510_6, addr_positional[24171:24168], addr_6042_7);

wire[31:0] addr_6043_7;

Selector_2 s6043_7(wires_1510_6[3], addr_1510_6, addr_positional[24175:24172], addr_6043_7);

wire[31:0] addr_6044_7;

Selector_2 s6044_7(wires_1511_6[0], addr_1511_6, addr_positional[24179:24176], addr_6044_7);

wire[31:0] addr_6045_7;

Selector_2 s6045_7(wires_1511_6[1], addr_1511_6, addr_positional[24183:24180], addr_6045_7);

wire[31:0] addr_6046_7;

Selector_2 s6046_7(wires_1511_6[2], addr_1511_6, addr_positional[24187:24184], addr_6046_7);

wire[31:0] addr_6047_7;

Selector_2 s6047_7(wires_1511_6[3], addr_1511_6, addr_positional[24191:24188], addr_6047_7);

wire[31:0] addr_6048_7;

Selector_2 s6048_7(wires_1512_6[0], addr_1512_6, addr_positional[24195:24192], addr_6048_7);

wire[31:0] addr_6049_7;

Selector_2 s6049_7(wires_1512_6[1], addr_1512_6, addr_positional[24199:24196], addr_6049_7);

wire[31:0] addr_6050_7;

Selector_2 s6050_7(wires_1512_6[2], addr_1512_6, addr_positional[24203:24200], addr_6050_7);

wire[31:0] addr_6051_7;

Selector_2 s6051_7(wires_1512_6[3], addr_1512_6, addr_positional[24207:24204], addr_6051_7);

wire[31:0] addr_6052_7;

Selector_2 s6052_7(wires_1513_6[0], addr_1513_6, addr_positional[24211:24208], addr_6052_7);

wire[31:0] addr_6053_7;

Selector_2 s6053_7(wires_1513_6[1], addr_1513_6, addr_positional[24215:24212], addr_6053_7);

wire[31:0] addr_6054_7;

Selector_2 s6054_7(wires_1513_6[2], addr_1513_6, addr_positional[24219:24216], addr_6054_7);

wire[31:0] addr_6055_7;

Selector_2 s6055_7(wires_1513_6[3], addr_1513_6, addr_positional[24223:24220], addr_6055_7);

wire[31:0] addr_6056_7;

Selector_2 s6056_7(wires_1514_6[0], addr_1514_6, addr_positional[24227:24224], addr_6056_7);

wire[31:0] addr_6057_7;

Selector_2 s6057_7(wires_1514_6[1], addr_1514_6, addr_positional[24231:24228], addr_6057_7);

wire[31:0] addr_6058_7;

Selector_2 s6058_7(wires_1514_6[2], addr_1514_6, addr_positional[24235:24232], addr_6058_7);

wire[31:0] addr_6059_7;

Selector_2 s6059_7(wires_1514_6[3], addr_1514_6, addr_positional[24239:24236], addr_6059_7);

wire[31:0] addr_6060_7;

Selector_2 s6060_7(wires_1515_6[0], addr_1515_6, addr_positional[24243:24240], addr_6060_7);

wire[31:0] addr_6061_7;

Selector_2 s6061_7(wires_1515_6[1], addr_1515_6, addr_positional[24247:24244], addr_6061_7);

wire[31:0] addr_6062_7;

Selector_2 s6062_7(wires_1515_6[2], addr_1515_6, addr_positional[24251:24248], addr_6062_7);

wire[31:0] addr_6063_7;

Selector_2 s6063_7(wires_1515_6[3], addr_1515_6, addr_positional[24255:24252], addr_6063_7);

wire[31:0] addr_6064_7;

Selector_2 s6064_7(wires_1516_6[0], addr_1516_6, addr_positional[24259:24256], addr_6064_7);

wire[31:0] addr_6065_7;

Selector_2 s6065_7(wires_1516_6[1], addr_1516_6, addr_positional[24263:24260], addr_6065_7);

wire[31:0] addr_6066_7;

Selector_2 s6066_7(wires_1516_6[2], addr_1516_6, addr_positional[24267:24264], addr_6066_7);

wire[31:0] addr_6067_7;

Selector_2 s6067_7(wires_1516_6[3], addr_1516_6, addr_positional[24271:24268], addr_6067_7);

wire[31:0] addr_6068_7;

Selector_2 s6068_7(wires_1517_6[0], addr_1517_6, addr_positional[24275:24272], addr_6068_7);

wire[31:0] addr_6069_7;

Selector_2 s6069_7(wires_1517_6[1], addr_1517_6, addr_positional[24279:24276], addr_6069_7);

wire[31:0] addr_6070_7;

Selector_2 s6070_7(wires_1517_6[2], addr_1517_6, addr_positional[24283:24280], addr_6070_7);

wire[31:0] addr_6071_7;

Selector_2 s6071_7(wires_1517_6[3], addr_1517_6, addr_positional[24287:24284], addr_6071_7);

wire[31:0] addr_6072_7;

Selector_2 s6072_7(wires_1518_6[0], addr_1518_6, addr_positional[24291:24288], addr_6072_7);

wire[31:0] addr_6073_7;

Selector_2 s6073_7(wires_1518_6[1], addr_1518_6, addr_positional[24295:24292], addr_6073_7);

wire[31:0] addr_6074_7;

Selector_2 s6074_7(wires_1518_6[2], addr_1518_6, addr_positional[24299:24296], addr_6074_7);

wire[31:0] addr_6075_7;

Selector_2 s6075_7(wires_1518_6[3], addr_1518_6, addr_positional[24303:24300], addr_6075_7);

wire[31:0] addr_6076_7;

Selector_2 s6076_7(wires_1519_6[0], addr_1519_6, addr_positional[24307:24304], addr_6076_7);

wire[31:0] addr_6077_7;

Selector_2 s6077_7(wires_1519_6[1], addr_1519_6, addr_positional[24311:24308], addr_6077_7);

wire[31:0] addr_6078_7;

Selector_2 s6078_7(wires_1519_6[2], addr_1519_6, addr_positional[24315:24312], addr_6078_7);

wire[31:0] addr_6079_7;

Selector_2 s6079_7(wires_1519_6[3], addr_1519_6, addr_positional[24319:24316], addr_6079_7);

wire[31:0] addr_6080_7;

Selector_2 s6080_7(wires_1520_6[0], addr_1520_6, addr_positional[24323:24320], addr_6080_7);

wire[31:0] addr_6081_7;

Selector_2 s6081_7(wires_1520_6[1], addr_1520_6, addr_positional[24327:24324], addr_6081_7);

wire[31:0] addr_6082_7;

Selector_2 s6082_7(wires_1520_6[2], addr_1520_6, addr_positional[24331:24328], addr_6082_7);

wire[31:0] addr_6083_7;

Selector_2 s6083_7(wires_1520_6[3], addr_1520_6, addr_positional[24335:24332], addr_6083_7);

wire[31:0] addr_6084_7;

Selector_2 s6084_7(wires_1521_6[0], addr_1521_6, addr_positional[24339:24336], addr_6084_7);

wire[31:0] addr_6085_7;

Selector_2 s6085_7(wires_1521_6[1], addr_1521_6, addr_positional[24343:24340], addr_6085_7);

wire[31:0] addr_6086_7;

Selector_2 s6086_7(wires_1521_6[2], addr_1521_6, addr_positional[24347:24344], addr_6086_7);

wire[31:0] addr_6087_7;

Selector_2 s6087_7(wires_1521_6[3], addr_1521_6, addr_positional[24351:24348], addr_6087_7);

wire[31:0] addr_6088_7;

Selector_2 s6088_7(wires_1522_6[0], addr_1522_6, addr_positional[24355:24352], addr_6088_7);

wire[31:0] addr_6089_7;

Selector_2 s6089_7(wires_1522_6[1], addr_1522_6, addr_positional[24359:24356], addr_6089_7);

wire[31:0] addr_6090_7;

Selector_2 s6090_7(wires_1522_6[2], addr_1522_6, addr_positional[24363:24360], addr_6090_7);

wire[31:0] addr_6091_7;

Selector_2 s6091_7(wires_1522_6[3], addr_1522_6, addr_positional[24367:24364], addr_6091_7);

wire[31:0] addr_6092_7;

Selector_2 s6092_7(wires_1523_6[0], addr_1523_6, addr_positional[24371:24368], addr_6092_7);

wire[31:0] addr_6093_7;

Selector_2 s6093_7(wires_1523_6[1], addr_1523_6, addr_positional[24375:24372], addr_6093_7);

wire[31:0] addr_6094_7;

Selector_2 s6094_7(wires_1523_6[2], addr_1523_6, addr_positional[24379:24376], addr_6094_7);

wire[31:0] addr_6095_7;

Selector_2 s6095_7(wires_1523_6[3], addr_1523_6, addr_positional[24383:24380], addr_6095_7);

wire[31:0] addr_6096_7;

Selector_2 s6096_7(wires_1524_6[0], addr_1524_6, addr_positional[24387:24384], addr_6096_7);

wire[31:0] addr_6097_7;

Selector_2 s6097_7(wires_1524_6[1], addr_1524_6, addr_positional[24391:24388], addr_6097_7);

wire[31:0] addr_6098_7;

Selector_2 s6098_7(wires_1524_6[2], addr_1524_6, addr_positional[24395:24392], addr_6098_7);

wire[31:0] addr_6099_7;

Selector_2 s6099_7(wires_1524_6[3], addr_1524_6, addr_positional[24399:24396], addr_6099_7);

wire[31:0] addr_6100_7;

Selector_2 s6100_7(wires_1525_6[0], addr_1525_6, addr_positional[24403:24400], addr_6100_7);

wire[31:0] addr_6101_7;

Selector_2 s6101_7(wires_1525_6[1], addr_1525_6, addr_positional[24407:24404], addr_6101_7);

wire[31:0] addr_6102_7;

Selector_2 s6102_7(wires_1525_6[2], addr_1525_6, addr_positional[24411:24408], addr_6102_7);

wire[31:0] addr_6103_7;

Selector_2 s6103_7(wires_1525_6[3], addr_1525_6, addr_positional[24415:24412], addr_6103_7);

wire[31:0] addr_6104_7;

Selector_2 s6104_7(wires_1526_6[0], addr_1526_6, addr_positional[24419:24416], addr_6104_7);

wire[31:0] addr_6105_7;

Selector_2 s6105_7(wires_1526_6[1], addr_1526_6, addr_positional[24423:24420], addr_6105_7);

wire[31:0] addr_6106_7;

Selector_2 s6106_7(wires_1526_6[2], addr_1526_6, addr_positional[24427:24424], addr_6106_7);

wire[31:0] addr_6107_7;

Selector_2 s6107_7(wires_1526_6[3], addr_1526_6, addr_positional[24431:24428], addr_6107_7);

wire[31:0] addr_6108_7;

Selector_2 s6108_7(wires_1527_6[0], addr_1527_6, addr_positional[24435:24432], addr_6108_7);

wire[31:0] addr_6109_7;

Selector_2 s6109_7(wires_1527_6[1], addr_1527_6, addr_positional[24439:24436], addr_6109_7);

wire[31:0] addr_6110_7;

Selector_2 s6110_7(wires_1527_6[2], addr_1527_6, addr_positional[24443:24440], addr_6110_7);

wire[31:0] addr_6111_7;

Selector_2 s6111_7(wires_1527_6[3], addr_1527_6, addr_positional[24447:24444], addr_6111_7);

wire[31:0] addr_6112_7;

Selector_2 s6112_7(wires_1528_6[0], addr_1528_6, addr_positional[24451:24448], addr_6112_7);

wire[31:0] addr_6113_7;

Selector_2 s6113_7(wires_1528_6[1], addr_1528_6, addr_positional[24455:24452], addr_6113_7);

wire[31:0] addr_6114_7;

Selector_2 s6114_7(wires_1528_6[2], addr_1528_6, addr_positional[24459:24456], addr_6114_7);

wire[31:0] addr_6115_7;

Selector_2 s6115_7(wires_1528_6[3], addr_1528_6, addr_positional[24463:24460], addr_6115_7);

wire[31:0] addr_6116_7;

Selector_2 s6116_7(wires_1529_6[0], addr_1529_6, addr_positional[24467:24464], addr_6116_7);

wire[31:0] addr_6117_7;

Selector_2 s6117_7(wires_1529_6[1], addr_1529_6, addr_positional[24471:24468], addr_6117_7);

wire[31:0] addr_6118_7;

Selector_2 s6118_7(wires_1529_6[2], addr_1529_6, addr_positional[24475:24472], addr_6118_7);

wire[31:0] addr_6119_7;

Selector_2 s6119_7(wires_1529_6[3], addr_1529_6, addr_positional[24479:24476], addr_6119_7);

wire[31:0] addr_6120_7;

Selector_2 s6120_7(wires_1530_6[0], addr_1530_6, addr_positional[24483:24480], addr_6120_7);

wire[31:0] addr_6121_7;

Selector_2 s6121_7(wires_1530_6[1], addr_1530_6, addr_positional[24487:24484], addr_6121_7);

wire[31:0] addr_6122_7;

Selector_2 s6122_7(wires_1530_6[2], addr_1530_6, addr_positional[24491:24488], addr_6122_7);

wire[31:0] addr_6123_7;

Selector_2 s6123_7(wires_1530_6[3], addr_1530_6, addr_positional[24495:24492], addr_6123_7);

wire[31:0] addr_6124_7;

Selector_2 s6124_7(wires_1531_6[0], addr_1531_6, addr_positional[24499:24496], addr_6124_7);

wire[31:0] addr_6125_7;

Selector_2 s6125_7(wires_1531_6[1], addr_1531_6, addr_positional[24503:24500], addr_6125_7);

wire[31:0] addr_6126_7;

Selector_2 s6126_7(wires_1531_6[2], addr_1531_6, addr_positional[24507:24504], addr_6126_7);

wire[31:0] addr_6127_7;

Selector_2 s6127_7(wires_1531_6[3], addr_1531_6, addr_positional[24511:24508], addr_6127_7);

wire[31:0] addr_6128_7;

Selector_2 s6128_7(wires_1532_6[0], addr_1532_6, addr_positional[24515:24512], addr_6128_7);

wire[31:0] addr_6129_7;

Selector_2 s6129_7(wires_1532_6[1], addr_1532_6, addr_positional[24519:24516], addr_6129_7);

wire[31:0] addr_6130_7;

Selector_2 s6130_7(wires_1532_6[2], addr_1532_6, addr_positional[24523:24520], addr_6130_7);

wire[31:0] addr_6131_7;

Selector_2 s6131_7(wires_1532_6[3], addr_1532_6, addr_positional[24527:24524], addr_6131_7);

wire[31:0] addr_6132_7;

Selector_2 s6132_7(wires_1533_6[0], addr_1533_6, addr_positional[24531:24528], addr_6132_7);

wire[31:0] addr_6133_7;

Selector_2 s6133_7(wires_1533_6[1], addr_1533_6, addr_positional[24535:24532], addr_6133_7);

wire[31:0] addr_6134_7;

Selector_2 s6134_7(wires_1533_6[2], addr_1533_6, addr_positional[24539:24536], addr_6134_7);

wire[31:0] addr_6135_7;

Selector_2 s6135_7(wires_1533_6[3], addr_1533_6, addr_positional[24543:24540], addr_6135_7);

wire[31:0] addr_6136_7;

Selector_2 s6136_7(wires_1534_6[0], addr_1534_6, addr_positional[24547:24544], addr_6136_7);

wire[31:0] addr_6137_7;

Selector_2 s6137_7(wires_1534_6[1], addr_1534_6, addr_positional[24551:24548], addr_6137_7);

wire[31:0] addr_6138_7;

Selector_2 s6138_7(wires_1534_6[2], addr_1534_6, addr_positional[24555:24552], addr_6138_7);

wire[31:0] addr_6139_7;

Selector_2 s6139_7(wires_1534_6[3], addr_1534_6, addr_positional[24559:24556], addr_6139_7);

wire[31:0] addr_6140_7;

Selector_2 s6140_7(wires_1535_6[0], addr_1535_6, addr_positional[24563:24560], addr_6140_7);

wire[31:0] addr_6141_7;

Selector_2 s6141_7(wires_1535_6[1], addr_1535_6, addr_positional[24567:24564], addr_6141_7);

wire[31:0] addr_6142_7;

Selector_2 s6142_7(wires_1535_6[2], addr_1535_6, addr_positional[24571:24568], addr_6142_7);

wire[31:0] addr_6143_7;

Selector_2 s6143_7(wires_1535_6[3], addr_1535_6, addr_positional[24575:24572], addr_6143_7);

wire[31:0] addr_6144_7;

Selector_2 s6144_7(wires_1536_6[0], addr_1536_6, addr_positional[24579:24576], addr_6144_7);

wire[31:0] addr_6145_7;

Selector_2 s6145_7(wires_1536_6[1], addr_1536_6, addr_positional[24583:24580], addr_6145_7);

wire[31:0] addr_6146_7;

Selector_2 s6146_7(wires_1536_6[2], addr_1536_6, addr_positional[24587:24584], addr_6146_7);

wire[31:0] addr_6147_7;

Selector_2 s6147_7(wires_1536_6[3], addr_1536_6, addr_positional[24591:24588], addr_6147_7);

wire[31:0] addr_6148_7;

Selector_2 s6148_7(wires_1537_6[0], addr_1537_6, addr_positional[24595:24592], addr_6148_7);

wire[31:0] addr_6149_7;

Selector_2 s6149_7(wires_1537_6[1], addr_1537_6, addr_positional[24599:24596], addr_6149_7);

wire[31:0] addr_6150_7;

Selector_2 s6150_7(wires_1537_6[2], addr_1537_6, addr_positional[24603:24600], addr_6150_7);

wire[31:0] addr_6151_7;

Selector_2 s6151_7(wires_1537_6[3], addr_1537_6, addr_positional[24607:24604], addr_6151_7);

wire[31:0] addr_6152_7;

Selector_2 s6152_7(wires_1538_6[0], addr_1538_6, addr_positional[24611:24608], addr_6152_7);

wire[31:0] addr_6153_7;

Selector_2 s6153_7(wires_1538_6[1], addr_1538_6, addr_positional[24615:24612], addr_6153_7);

wire[31:0] addr_6154_7;

Selector_2 s6154_7(wires_1538_6[2], addr_1538_6, addr_positional[24619:24616], addr_6154_7);

wire[31:0] addr_6155_7;

Selector_2 s6155_7(wires_1538_6[3], addr_1538_6, addr_positional[24623:24620], addr_6155_7);

wire[31:0] addr_6156_7;

Selector_2 s6156_7(wires_1539_6[0], addr_1539_6, addr_positional[24627:24624], addr_6156_7);

wire[31:0] addr_6157_7;

Selector_2 s6157_7(wires_1539_6[1], addr_1539_6, addr_positional[24631:24628], addr_6157_7);

wire[31:0] addr_6158_7;

Selector_2 s6158_7(wires_1539_6[2], addr_1539_6, addr_positional[24635:24632], addr_6158_7);

wire[31:0] addr_6159_7;

Selector_2 s6159_7(wires_1539_6[3], addr_1539_6, addr_positional[24639:24636], addr_6159_7);

wire[31:0] addr_6160_7;

Selector_2 s6160_7(wires_1540_6[0], addr_1540_6, addr_positional[24643:24640], addr_6160_7);

wire[31:0] addr_6161_7;

Selector_2 s6161_7(wires_1540_6[1], addr_1540_6, addr_positional[24647:24644], addr_6161_7);

wire[31:0] addr_6162_7;

Selector_2 s6162_7(wires_1540_6[2], addr_1540_6, addr_positional[24651:24648], addr_6162_7);

wire[31:0] addr_6163_7;

Selector_2 s6163_7(wires_1540_6[3], addr_1540_6, addr_positional[24655:24652], addr_6163_7);

wire[31:0] addr_6164_7;

Selector_2 s6164_7(wires_1541_6[0], addr_1541_6, addr_positional[24659:24656], addr_6164_7);

wire[31:0] addr_6165_7;

Selector_2 s6165_7(wires_1541_6[1], addr_1541_6, addr_positional[24663:24660], addr_6165_7);

wire[31:0] addr_6166_7;

Selector_2 s6166_7(wires_1541_6[2], addr_1541_6, addr_positional[24667:24664], addr_6166_7);

wire[31:0] addr_6167_7;

Selector_2 s6167_7(wires_1541_6[3], addr_1541_6, addr_positional[24671:24668], addr_6167_7);

wire[31:0] addr_6168_7;

Selector_2 s6168_7(wires_1542_6[0], addr_1542_6, addr_positional[24675:24672], addr_6168_7);

wire[31:0] addr_6169_7;

Selector_2 s6169_7(wires_1542_6[1], addr_1542_6, addr_positional[24679:24676], addr_6169_7);

wire[31:0] addr_6170_7;

Selector_2 s6170_7(wires_1542_6[2], addr_1542_6, addr_positional[24683:24680], addr_6170_7);

wire[31:0] addr_6171_7;

Selector_2 s6171_7(wires_1542_6[3], addr_1542_6, addr_positional[24687:24684], addr_6171_7);

wire[31:0] addr_6172_7;

Selector_2 s6172_7(wires_1543_6[0], addr_1543_6, addr_positional[24691:24688], addr_6172_7);

wire[31:0] addr_6173_7;

Selector_2 s6173_7(wires_1543_6[1], addr_1543_6, addr_positional[24695:24692], addr_6173_7);

wire[31:0] addr_6174_7;

Selector_2 s6174_7(wires_1543_6[2], addr_1543_6, addr_positional[24699:24696], addr_6174_7);

wire[31:0] addr_6175_7;

Selector_2 s6175_7(wires_1543_6[3], addr_1543_6, addr_positional[24703:24700], addr_6175_7);

wire[31:0] addr_6176_7;

Selector_2 s6176_7(wires_1544_6[0], addr_1544_6, addr_positional[24707:24704], addr_6176_7);

wire[31:0] addr_6177_7;

Selector_2 s6177_7(wires_1544_6[1], addr_1544_6, addr_positional[24711:24708], addr_6177_7);

wire[31:0] addr_6178_7;

Selector_2 s6178_7(wires_1544_6[2], addr_1544_6, addr_positional[24715:24712], addr_6178_7);

wire[31:0] addr_6179_7;

Selector_2 s6179_7(wires_1544_6[3], addr_1544_6, addr_positional[24719:24716], addr_6179_7);

wire[31:0] addr_6180_7;

Selector_2 s6180_7(wires_1545_6[0], addr_1545_6, addr_positional[24723:24720], addr_6180_7);

wire[31:0] addr_6181_7;

Selector_2 s6181_7(wires_1545_6[1], addr_1545_6, addr_positional[24727:24724], addr_6181_7);

wire[31:0] addr_6182_7;

Selector_2 s6182_7(wires_1545_6[2], addr_1545_6, addr_positional[24731:24728], addr_6182_7);

wire[31:0] addr_6183_7;

Selector_2 s6183_7(wires_1545_6[3], addr_1545_6, addr_positional[24735:24732], addr_6183_7);

wire[31:0] addr_6184_7;

Selector_2 s6184_7(wires_1546_6[0], addr_1546_6, addr_positional[24739:24736], addr_6184_7);

wire[31:0] addr_6185_7;

Selector_2 s6185_7(wires_1546_6[1], addr_1546_6, addr_positional[24743:24740], addr_6185_7);

wire[31:0] addr_6186_7;

Selector_2 s6186_7(wires_1546_6[2], addr_1546_6, addr_positional[24747:24744], addr_6186_7);

wire[31:0] addr_6187_7;

Selector_2 s6187_7(wires_1546_6[3], addr_1546_6, addr_positional[24751:24748], addr_6187_7);

wire[31:0] addr_6188_7;

Selector_2 s6188_7(wires_1547_6[0], addr_1547_6, addr_positional[24755:24752], addr_6188_7);

wire[31:0] addr_6189_7;

Selector_2 s6189_7(wires_1547_6[1], addr_1547_6, addr_positional[24759:24756], addr_6189_7);

wire[31:0] addr_6190_7;

Selector_2 s6190_7(wires_1547_6[2], addr_1547_6, addr_positional[24763:24760], addr_6190_7);

wire[31:0] addr_6191_7;

Selector_2 s6191_7(wires_1547_6[3], addr_1547_6, addr_positional[24767:24764], addr_6191_7);

wire[31:0] addr_6192_7;

Selector_2 s6192_7(wires_1548_6[0], addr_1548_6, addr_positional[24771:24768], addr_6192_7);

wire[31:0] addr_6193_7;

Selector_2 s6193_7(wires_1548_6[1], addr_1548_6, addr_positional[24775:24772], addr_6193_7);

wire[31:0] addr_6194_7;

Selector_2 s6194_7(wires_1548_6[2], addr_1548_6, addr_positional[24779:24776], addr_6194_7);

wire[31:0] addr_6195_7;

Selector_2 s6195_7(wires_1548_6[3], addr_1548_6, addr_positional[24783:24780], addr_6195_7);

wire[31:0] addr_6196_7;

Selector_2 s6196_7(wires_1549_6[0], addr_1549_6, addr_positional[24787:24784], addr_6196_7);

wire[31:0] addr_6197_7;

Selector_2 s6197_7(wires_1549_6[1], addr_1549_6, addr_positional[24791:24788], addr_6197_7);

wire[31:0] addr_6198_7;

Selector_2 s6198_7(wires_1549_6[2], addr_1549_6, addr_positional[24795:24792], addr_6198_7);

wire[31:0] addr_6199_7;

Selector_2 s6199_7(wires_1549_6[3], addr_1549_6, addr_positional[24799:24796], addr_6199_7);

wire[31:0] addr_6200_7;

Selector_2 s6200_7(wires_1550_6[0], addr_1550_6, addr_positional[24803:24800], addr_6200_7);

wire[31:0] addr_6201_7;

Selector_2 s6201_7(wires_1550_6[1], addr_1550_6, addr_positional[24807:24804], addr_6201_7);

wire[31:0] addr_6202_7;

Selector_2 s6202_7(wires_1550_6[2], addr_1550_6, addr_positional[24811:24808], addr_6202_7);

wire[31:0] addr_6203_7;

Selector_2 s6203_7(wires_1550_6[3], addr_1550_6, addr_positional[24815:24812], addr_6203_7);

wire[31:0] addr_6204_7;

Selector_2 s6204_7(wires_1551_6[0], addr_1551_6, addr_positional[24819:24816], addr_6204_7);

wire[31:0] addr_6205_7;

Selector_2 s6205_7(wires_1551_6[1], addr_1551_6, addr_positional[24823:24820], addr_6205_7);

wire[31:0] addr_6206_7;

Selector_2 s6206_7(wires_1551_6[2], addr_1551_6, addr_positional[24827:24824], addr_6206_7);

wire[31:0] addr_6207_7;

Selector_2 s6207_7(wires_1551_6[3], addr_1551_6, addr_positional[24831:24828], addr_6207_7);

wire[31:0] addr_6208_7;

Selector_2 s6208_7(wires_1552_6[0], addr_1552_6, addr_positional[24835:24832], addr_6208_7);

wire[31:0] addr_6209_7;

Selector_2 s6209_7(wires_1552_6[1], addr_1552_6, addr_positional[24839:24836], addr_6209_7);

wire[31:0] addr_6210_7;

Selector_2 s6210_7(wires_1552_6[2], addr_1552_6, addr_positional[24843:24840], addr_6210_7);

wire[31:0] addr_6211_7;

Selector_2 s6211_7(wires_1552_6[3], addr_1552_6, addr_positional[24847:24844], addr_6211_7);

wire[31:0] addr_6212_7;

Selector_2 s6212_7(wires_1553_6[0], addr_1553_6, addr_positional[24851:24848], addr_6212_7);

wire[31:0] addr_6213_7;

Selector_2 s6213_7(wires_1553_6[1], addr_1553_6, addr_positional[24855:24852], addr_6213_7);

wire[31:0] addr_6214_7;

Selector_2 s6214_7(wires_1553_6[2], addr_1553_6, addr_positional[24859:24856], addr_6214_7);

wire[31:0] addr_6215_7;

Selector_2 s6215_7(wires_1553_6[3], addr_1553_6, addr_positional[24863:24860], addr_6215_7);

wire[31:0] addr_6216_7;

Selector_2 s6216_7(wires_1554_6[0], addr_1554_6, addr_positional[24867:24864], addr_6216_7);

wire[31:0] addr_6217_7;

Selector_2 s6217_7(wires_1554_6[1], addr_1554_6, addr_positional[24871:24868], addr_6217_7);

wire[31:0] addr_6218_7;

Selector_2 s6218_7(wires_1554_6[2], addr_1554_6, addr_positional[24875:24872], addr_6218_7);

wire[31:0] addr_6219_7;

Selector_2 s6219_7(wires_1554_6[3], addr_1554_6, addr_positional[24879:24876], addr_6219_7);

wire[31:0] addr_6220_7;

Selector_2 s6220_7(wires_1555_6[0], addr_1555_6, addr_positional[24883:24880], addr_6220_7);

wire[31:0] addr_6221_7;

Selector_2 s6221_7(wires_1555_6[1], addr_1555_6, addr_positional[24887:24884], addr_6221_7);

wire[31:0] addr_6222_7;

Selector_2 s6222_7(wires_1555_6[2], addr_1555_6, addr_positional[24891:24888], addr_6222_7);

wire[31:0] addr_6223_7;

Selector_2 s6223_7(wires_1555_6[3], addr_1555_6, addr_positional[24895:24892], addr_6223_7);

wire[31:0] addr_6224_7;

Selector_2 s6224_7(wires_1556_6[0], addr_1556_6, addr_positional[24899:24896], addr_6224_7);

wire[31:0] addr_6225_7;

Selector_2 s6225_7(wires_1556_6[1], addr_1556_6, addr_positional[24903:24900], addr_6225_7);

wire[31:0] addr_6226_7;

Selector_2 s6226_7(wires_1556_6[2], addr_1556_6, addr_positional[24907:24904], addr_6226_7);

wire[31:0] addr_6227_7;

Selector_2 s6227_7(wires_1556_6[3], addr_1556_6, addr_positional[24911:24908], addr_6227_7);

wire[31:0] addr_6228_7;

Selector_2 s6228_7(wires_1557_6[0], addr_1557_6, addr_positional[24915:24912], addr_6228_7);

wire[31:0] addr_6229_7;

Selector_2 s6229_7(wires_1557_6[1], addr_1557_6, addr_positional[24919:24916], addr_6229_7);

wire[31:0] addr_6230_7;

Selector_2 s6230_7(wires_1557_6[2], addr_1557_6, addr_positional[24923:24920], addr_6230_7);

wire[31:0] addr_6231_7;

Selector_2 s6231_7(wires_1557_6[3], addr_1557_6, addr_positional[24927:24924], addr_6231_7);

wire[31:0] addr_6232_7;

Selector_2 s6232_7(wires_1558_6[0], addr_1558_6, addr_positional[24931:24928], addr_6232_7);

wire[31:0] addr_6233_7;

Selector_2 s6233_7(wires_1558_6[1], addr_1558_6, addr_positional[24935:24932], addr_6233_7);

wire[31:0] addr_6234_7;

Selector_2 s6234_7(wires_1558_6[2], addr_1558_6, addr_positional[24939:24936], addr_6234_7);

wire[31:0] addr_6235_7;

Selector_2 s6235_7(wires_1558_6[3], addr_1558_6, addr_positional[24943:24940], addr_6235_7);

wire[31:0] addr_6236_7;

Selector_2 s6236_7(wires_1559_6[0], addr_1559_6, addr_positional[24947:24944], addr_6236_7);

wire[31:0] addr_6237_7;

Selector_2 s6237_7(wires_1559_6[1], addr_1559_6, addr_positional[24951:24948], addr_6237_7);

wire[31:0] addr_6238_7;

Selector_2 s6238_7(wires_1559_6[2], addr_1559_6, addr_positional[24955:24952], addr_6238_7);

wire[31:0] addr_6239_7;

Selector_2 s6239_7(wires_1559_6[3], addr_1559_6, addr_positional[24959:24956], addr_6239_7);

wire[31:0] addr_6240_7;

Selector_2 s6240_7(wires_1560_6[0], addr_1560_6, addr_positional[24963:24960], addr_6240_7);

wire[31:0] addr_6241_7;

Selector_2 s6241_7(wires_1560_6[1], addr_1560_6, addr_positional[24967:24964], addr_6241_7);

wire[31:0] addr_6242_7;

Selector_2 s6242_7(wires_1560_6[2], addr_1560_6, addr_positional[24971:24968], addr_6242_7);

wire[31:0] addr_6243_7;

Selector_2 s6243_7(wires_1560_6[3], addr_1560_6, addr_positional[24975:24972], addr_6243_7);

wire[31:0] addr_6244_7;

Selector_2 s6244_7(wires_1561_6[0], addr_1561_6, addr_positional[24979:24976], addr_6244_7);

wire[31:0] addr_6245_7;

Selector_2 s6245_7(wires_1561_6[1], addr_1561_6, addr_positional[24983:24980], addr_6245_7);

wire[31:0] addr_6246_7;

Selector_2 s6246_7(wires_1561_6[2], addr_1561_6, addr_positional[24987:24984], addr_6246_7);

wire[31:0] addr_6247_7;

Selector_2 s6247_7(wires_1561_6[3], addr_1561_6, addr_positional[24991:24988], addr_6247_7);

wire[31:0] addr_6248_7;

Selector_2 s6248_7(wires_1562_6[0], addr_1562_6, addr_positional[24995:24992], addr_6248_7);

wire[31:0] addr_6249_7;

Selector_2 s6249_7(wires_1562_6[1], addr_1562_6, addr_positional[24999:24996], addr_6249_7);

wire[31:0] addr_6250_7;

Selector_2 s6250_7(wires_1562_6[2], addr_1562_6, addr_positional[25003:25000], addr_6250_7);

wire[31:0] addr_6251_7;

Selector_2 s6251_7(wires_1562_6[3], addr_1562_6, addr_positional[25007:25004], addr_6251_7);

wire[31:0] addr_6252_7;

Selector_2 s6252_7(wires_1563_6[0], addr_1563_6, addr_positional[25011:25008], addr_6252_7);

wire[31:0] addr_6253_7;

Selector_2 s6253_7(wires_1563_6[1], addr_1563_6, addr_positional[25015:25012], addr_6253_7);

wire[31:0] addr_6254_7;

Selector_2 s6254_7(wires_1563_6[2], addr_1563_6, addr_positional[25019:25016], addr_6254_7);

wire[31:0] addr_6255_7;

Selector_2 s6255_7(wires_1563_6[3], addr_1563_6, addr_positional[25023:25020], addr_6255_7);

wire[31:0] addr_6256_7;

Selector_2 s6256_7(wires_1564_6[0], addr_1564_6, addr_positional[25027:25024], addr_6256_7);

wire[31:0] addr_6257_7;

Selector_2 s6257_7(wires_1564_6[1], addr_1564_6, addr_positional[25031:25028], addr_6257_7);

wire[31:0] addr_6258_7;

Selector_2 s6258_7(wires_1564_6[2], addr_1564_6, addr_positional[25035:25032], addr_6258_7);

wire[31:0] addr_6259_7;

Selector_2 s6259_7(wires_1564_6[3], addr_1564_6, addr_positional[25039:25036], addr_6259_7);

wire[31:0] addr_6260_7;

Selector_2 s6260_7(wires_1565_6[0], addr_1565_6, addr_positional[25043:25040], addr_6260_7);

wire[31:0] addr_6261_7;

Selector_2 s6261_7(wires_1565_6[1], addr_1565_6, addr_positional[25047:25044], addr_6261_7);

wire[31:0] addr_6262_7;

Selector_2 s6262_7(wires_1565_6[2], addr_1565_6, addr_positional[25051:25048], addr_6262_7);

wire[31:0] addr_6263_7;

Selector_2 s6263_7(wires_1565_6[3], addr_1565_6, addr_positional[25055:25052], addr_6263_7);

wire[31:0] addr_6264_7;

Selector_2 s6264_7(wires_1566_6[0], addr_1566_6, addr_positional[25059:25056], addr_6264_7);

wire[31:0] addr_6265_7;

Selector_2 s6265_7(wires_1566_6[1], addr_1566_6, addr_positional[25063:25060], addr_6265_7);

wire[31:0] addr_6266_7;

Selector_2 s6266_7(wires_1566_6[2], addr_1566_6, addr_positional[25067:25064], addr_6266_7);

wire[31:0] addr_6267_7;

Selector_2 s6267_7(wires_1566_6[3], addr_1566_6, addr_positional[25071:25068], addr_6267_7);

wire[31:0] addr_6268_7;

Selector_2 s6268_7(wires_1567_6[0], addr_1567_6, addr_positional[25075:25072], addr_6268_7);

wire[31:0] addr_6269_7;

Selector_2 s6269_7(wires_1567_6[1], addr_1567_6, addr_positional[25079:25076], addr_6269_7);

wire[31:0] addr_6270_7;

Selector_2 s6270_7(wires_1567_6[2], addr_1567_6, addr_positional[25083:25080], addr_6270_7);

wire[31:0] addr_6271_7;

Selector_2 s6271_7(wires_1567_6[3], addr_1567_6, addr_positional[25087:25084], addr_6271_7);

wire[31:0] addr_6272_7;

Selector_2 s6272_7(wires_1568_6[0], addr_1568_6, addr_positional[25091:25088], addr_6272_7);

wire[31:0] addr_6273_7;

Selector_2 s6273_7(wires_1568_6[1], addr_1568_6, addr_positional[25095:25092], addr_6273_7);

wire[31:0] addr_6274_7;

Selector_2 s6274_7(wires_1568_6[2], addr_1568_6, addr_positional[25099:25096], addr_6274_7);

wire[31:0] addr_6275_7;

Selector_2 s6275_7(wires_1568_6[3], addr_1568_6, addr_positional[25103:25100], addr_6275_7);

wire[31:0] addr_6276_7;

Selector_2 s6276_7(wires_1569_6[0], addr_1569_6, addr_positional[25107:25104], addr_6276_7);

wire[31:0] addr_6277_7;

Selector_2 s6277_7(wires_1569_6[1], addr_1569_6, addr_positional[25111:25108], addr_6277_7);

wire[31:0] addr_6278_7;

Selector_2 s6278_7(wires_1569_6[2], addr_1569_6, addr_positional[25115:25112], addr_6278_7);

wire[31:0] addr_6279_7;

Selector_2 s6279_7(wires_1569_6[3], addr_1569_6, addr_positional[25119:25116], addr_6279_7);

wire[31:0] addr_6280_7;

Selector_2 s6280_7(wires_1570_6[0], addr_1570_6, addr_positional[25123:25120], addr_6280_7);

wire[31:0] addr_6281_7;

Selector_2 s6281_7(wires_1570_6[1], addr_1570_6, addr_positional[25127:25124], addr_6281_7);

wire[31:0] addr_6282_7;

Selector_2 s6282_7(wires_1570_6[2], addr_1570_6, addr_positional[25131:25128], addr_6282_7);

wire[31:0] addr_6283_7;

Selector_2 s6283_7(wires_1570_6[3], addr_1570_6, addr_positional[25135:25132], addr_6283_7);

wire[31:0] addr_6284_7;

Selector_2 s6284_7(wires_1571_6[0], addr_1571_6, addr_positional[25139:25136], addr_6284_7);

wire[31:0] addr_6285_7;

Selector_2 s6285_7(wires_1571_6[1], addr_1571_6, addr_positional[25143:25140], addr_6285_7);

wire[31:0] addr_6286_7;

Selector_2 s6286_7(wires_1571_6[2], addr_1571_6, addr_positional[25147:25144], addr_6286_7);

wire[31:0] addr_6287_7;

Selector_2 s6287_7(wires_1571_6[3], addr_1571_6, addr_positional[25151:25148], addr_6287_7);

wire[31:0] addr_6288_7;

Selector_2 s6288_7(wires_1572_6[0], addr_1572_6, addr_positional[25155:25152], addr_6288_7);

wire[31:0] addr_6289_7;

Selector_2 s6289_7(wires_1572_6[1], addr_1572_6, addr_positional[25159:25156], addr_6289_7);

wire[31:0] addr_6290_7;

Selector_2 s6290_7(wires_1572_6[2], addr_1572_6, addr_positional[25163:25160], addr_6290_7);

wire[31:0] addr_6291_7;

Selector_2 s6291_7(wires_1572_6[3], addr_1572_6, addr_positional[25167:25164], addr_6291_7);

wire[31:0] addr_6292_7;

Selector_2 s6292_7(wires_1573_6[0], addr_1573_6, addr_positional[25171:25168], addr_6292_7);

wire[31:0] addr_6293_7;

Selector_2 s6293_7(wires_1573_6[1], addr_1573_6, addr_positional[25175:25172], addr_6293_7);

wire[31:0] addr_6294_7;

Selector_2 s6294_7(wires_1573_6[2], addr_1573_6, addr_positional[25179:25176], addr_6294_7);

wire[31:0] addr_6295_7;

Selector_2 s6295_7(wires_1573_6[3], addr_1573_6, addr_positional[25183:25180], addr_6295_7);

wire[31:0] addr_6296_7;

Selector_2 s6296_7(wires_1574_6[0], addr_1574_6, addr_positional[25187:25184], addr_6296_7);

wire[31:0] addr_6297_7;

Selector_2 s6297_7(wires_1574_6[1], addr_1574_6, addr_positional[25191:25188], addr_6297_7);

wire[31:0] addr_6298_7;

Selector_2 s6298_7(wires_1574_6[2], addr_1574_6, addr_positional[25195:25192], addr_6298_7);

wire[31:0] addr_6299_7;

Selector_2 s6299_7(wires_1574_6[3], addr_1574_6, addr_positional[25199:25196], addr_6299_7);

wire[31:0] addr_6300_7;

Selector_2 s6300_7(wires_1575_6[0], addr_1575_6, addr_positional[25203:25200], addr_6300_7);

wire[31:0] addr_6301_7;

Selector_2 s6301_7(wires_1575_6[1], addr_1575_6, addr_positional[25207:25204], addr_6301_7);

wire[31:0] addr_6302_7;

Selector_2 s6302_7(wires_1575_6[2], addr_1575_6, addr_positional[25211:25208], addr_6302_7);

wire[31:0] addr_6303_7;

Selector_2 s6303_7(wires_1575_6[3], addr_1575_6, addr_positional[25215:25212], addr_6303_7);

wire[31:0] addr_6304_7;

Selector_2 s6304_7(wires_1576_6[0], addr_1576_6, addr_positional[25219:25216], addr_6304_7);

wire[31:0] addr_6305_7;

Selector_2 s6305_7(wires_1576_6[1], addr_1576_6, addr_positional[25223:25220], addr_6305_7);

wire[31:0] addr_6306_7;

Selector_2 s6306_7(wires_1576_6[2], addr_1576_6, addr_positional[25227:25224], addr_6306_7);

wire[31:0] addr_6307_7;

Selector_2 s6307_7(wires_1576_6[3], addr_1576_6, addr_positional[25231:25228], addr_6307_7);

wire[31:0] addr_6308_7;

Selector_2 s6308_7(wires_1577_6[0], addr_1577_6, addr_positional[25235:25232], addr_6308_7);

wire[31:0] addr_6309_7;

Selector_2 s6309_7(wires_1577_6[1], addr_1577_6, addr_positional[25239:25236], addr_6309_7);

wire[31:0] addr_6310_7;

Selector_2 s6310_7(wires_1577_6[2], addr_1577_6, addr_positional[25243:25240], addr_6310_7);

wire[31:0] addr_6311_7;

Selector_2 s6311_7(wires_1577_6[3], addr_1577_6, addr_positional[25247:25244], addr_6311_7);

wire[31:0] addr_6312_7;

Selector_2 s6312_7(wires_1578_6[0], addr_1578_6, addr_positional[25251:25248], addr_6312_7);

wire[31:0] addr_6313_7;

Selector_2 s6313_7(wires_1578_6[1], addr_1578_6, addr_positional[25255:25252], addr_6313_7);

wire[31:0] addr_6314_7;

Selector_2 s6314_7(wires_1578_6[2], addr_1578_6, addr_positional[25259:25256], addr_6314_7);

wire[31:0] addr_6315_7;

Selector_2 s6315_7(wires_1578_6[3], addr_1578_6, addr_positional[25263:25260], addr_6315_7);

wire[31:0] addr_6316_7;

Selector_2 s6316_7(wires_1579_6[0], addr_1579_6, addr_positional[25267:25264], addr_6316_7);

wire[31:0] addr_6317_7;

Selector_2 s6317_7(wires_1579_6[1], addr_1579_6, addr_positional[25271:25268], addr_6317_7);

wire[31:0] addr_6318_7;

Selector_2 s6318_7(wires_1579_6[2], addr_1579_6, addr_positional[25275:25272], addr_6318_7);

wire[31:0] addr_6319_7;

Selector_2 s6319_7(wires_1579_6[3], addr_1579_6, addr_positional[25279:25276], addr_6319_7);

wire[31:0] addr_6320_7;

Selector_2 s6320_7(wires_1580_6[0], addr_1580_6, addr_positional[25283:25280], addr_6320_7);

wire[31:0] addr_6321_7;

Selector_2 s6321_7(wires_1580_6[1], addr_1580_6, addr_positional[25287:25284], addr_6321_7);

wire[31:0] addr_6322_7;

Selector_2 s6322_7(wires_1580_6[2], addr_1580_6, addr_positional[25291:25288], addr_6322_7);

wire[31:0] addr_6323_7;

Selector_2 s6323_7(wires_1580_6[3], addr_1580_6, addr_positional[25295:25292], addr_6323_7);

wire[31:0] addr_6324_7;

Selector_2 s6324_7(wires_1581_6[0], addr_1581_6, addr_positional[25299:25296], addr_6324_7);

wire[31:0] addr_6325_7;

Selector_2 s6325_7(wires_1581_6[1], addr_1581_6, addr_positional[25303:25300], addr_6325_7);

wire[31:0] addr_6326_7;

Selector_2 s6326_7(wires_1581_6[2], addr_1581_6, addr_positional[25307:25304], addr_6326_7);

wire[31:0] addr_6327_7;

Selector_2 s6327_7(wires_1581_6[3], addr_1581_6, addr_positional[25311:25308], addr_6327_7);

wire[31:0] addr_6328_7;

Selector_2 s6328_7(wires_1582_6[0], addr_1582_6, addr_positional[25315:25312], addr_6328_7);

wire[31:0] addr_6329_7;

Selector_2 s6329_7(wires_1582_6[1], addr_1582_6, addr_positional[25319:25316], addr_6329_7);

wire[31:0] addr_6330_7;

Selector_2 s6330_7(wires_1582_6[2], addr_1582_6, addr_positional[25323:25320], addr_6330_7);

wire[31:0] addr_6331_7;

Selector_2 s6331_7(wires_1582_6[3], addr_1582_6, addr_positional[25327:25324], addr_6331_7);

wire[31:0] addr_6332_7;

Selector_2 s6332_7(wires_1583_6[0], addr_1583_6, addr_positional[25331:25328], addr_6332_7);

wire[31:0] addr_6333_7;

Selector_2 s6333_7(wires_1583_6[1], addr_1583_6, addr_positional[25335:25332], addr_6333_7);

wire[31:0] addr_6334_7;

Selector_2 s6334_7(wires_1583_6[2], addr_1583_6, addr_positional[25339:25336], addr_6334_7);

wire[31:0] addr_6335_7;

Selector_2 s6335_7(wires_1583_6[3], addr_1583_6, addr_positional[25343:25340], addr_6335_7);

wire[31:0] addr_6336_7;

Selector_2 s6336_7(wires_1584_6[0], addr_1584_6, addr_positional[25347:25344], addr_6336_7);

wire[31:0] addr_6337_7;

Selector_2 s6337_7(wires_1584_6[1], addr_1584_6, addr_positional[25351:25348], addr_6337_7);

wire[31:0] addr_6338_7;

Selector_2 s6338_7(wires_1584_6[2], addr_1584_6, addr_positional[25355:25352], addr_6338_7);

wire[31:0] addr_6339_7;

Selector_2 s6339_7(wires_1584_6[3], addr_1584_6, addr_positional[25359:25356], addr_6339_7);

wire[31:0] addr_6340_7;

Selector_2 s6340_7(wires_1585_6[0], addr_1585_6, addr_positional[25363:25360], addr_6340_7);

wire[31:0] addr_6341_7;

Selector_2 s6341_7(wires_1585_6[1], addr_1585_6, addr_positional[25367:25364], addr_6341_7);

wire[31:0] addr_6342_7;

Selector_2 s6342_7(wires_1585_6[2], addr_1585_6, addr_positional[25371:25368], addr_6342_7);

wire[31:0] addr_6343_7;

Selector_2 s6343_7(wires_1585_6[3], addr_1585_6, addr_positional[25375:25372], addr_6343_7);

wire[31:0] addr_6344_7;

Selector_2 s6344_7(wires_1586_6[0], addr_1586_6, addr_positional[25379:25376], addr_6344_7);

wire[31:0] addr_6345_7;

Selector_2 s6345_7(wires_1586_6[1], addr_1586_6, addr_positional[25383:25380], addr_6345_7);

wire[31:0] addr_6346_7;

Selector_2 s6346_7(wires_1586_6[2], addr_1586_6, addr_positional[25387:25384], addr_6346_7);

wire[31:0] addr_6347_7;

Selector_2 s6347_7(wires_1586_6[3], addr_1586_6, addr_positional[25391:25388], addr_6347_7);

wire[31:0] addr_6348_7;

Selector_2 s6348_7(wires_1587_6[0], addr_1587_6, addr_positional[25395:25392], addr_6348_7);

wire[31:0] addr_6349_7;

Selector_2 s6349_7(wires_1587_6[1], addr_1587_6, addr_positional[25399:25396], addr_6349_7);

wire[31:0] addr_6350_7;

Selector_2 s6350_7(wires_1587_6[2], addr_1587_6, addr_positional[25403:25400], addr_6350_7);

wire[31:0] addr_6351_7;

Selector_2 s6351_7(wires_1587_6[3], addr_1587_6, addr_positional[25407:25404], addr_6351_7);

wire[31:0] addr_6352_7;

Selector_2 s6352_7(wires_1588_6[0], addr_1588_6, addr_positional[25411:25408], addr_6352_7);

wire[31:0] addr_6353_7;

Selector_2 s6353_7(wires_1588_6[1], addr_1588_6, addr_positional[25415:25412], addr_6353_7);

wire[31:0] addr_6354_7;

Selector_2 s6354_7(wires_1588_6[2], addr_1588_6, addr_positional[25419:25416], addr_6354_7);

wire[31:0] addr_6355_7;

Selector_2 s6355_7(wires_1588_6[3], addr_1588_6, addr_positional[25423:25420], addr_6355_7);

wire[31:0] addr_6356_7;

Selector_2 s6356_7(wires_1589_6[0], addr_1589_6, addr_positional[25427:25424], addr_6356_7);

wire[31:0] addr_6357_7;

Selector_2 s6357_7(wires_1589_6[1], addr_1589_6, addr_positional[25431:25428], addr_6357_7);

wire[31:0] addr_6358_7;

Selector_2 s6358_7(wires_1589_6[2], addr_1589_6, addr_positional[25435:25432], addr_6358_7);

wire[31:0] addr_6359_7;

Selector_2 s6359_7(wires_1589_6[3], addr_1589_6, addr_positional[25439:25436], addr_6359_7);

wire[31:0] addr_6360_7;

Selector_2 s6360_7(wires_1590_6[0], addr_1590_6, addr_positional[25443:25440], addr_6360_7);

wire[31:0] addr_6361_7;

Selector_2 s6361_7(wires_1590_6[1], addr_1590_6, addr_positional[25447:25444], addr_6361_7);

wire[31:0] addr_6362_7;

Selector_2 s6362_7(wires_1590_6[2], addr_1590_6, addr_positional[25451:25448], addr_6362_7);

wire[31:0] addr_6363_7;

Selector_2 s6363_7(wires_1590_6[3], addr_1590_6, addr_positional[25455:25452], addr_6363_7);

wire[31:0] addr_6364_7;

Selector_2 s6364_7(wires_1591_6[0], addr_1591_6, addr_positional[25459:25456], addr_6364_7);

wire[31:0] addr_6365_7;

Selector_2 s6365_7(wires_1591_6[1], addr_1591_6, addr_positional[25463:25460], addr_6365_7);

wire[31:0] addr_6366_7;

Selector_2 s6366_7(wires_1591_6[2], addr_1591_6, addr_positional[25467:25464], addr_6366_7);

wire[31:0] addr_6367_7;

Selector_2 s6367_7(wires_1591_6[3], addr_1591_6, addr_positional[25471:25468], addr_6367_7);

wire[31:0] addr_6368_7;

Selector_2 s6368_7(wires_1592_6[0], addr_1592_6, addr_positional[25475:25472], addr_6368_7);

wire[31:0] addr_6369_7;

Selector_2 s6369_7(wires_1592_6[1], addr_1592_6, addr_positional[25479:25476], addr_6369_7);

wire[31:0] addr_6370_7;

Selector_2 s6370_7(wires_1592_6[2], addr_1592_6, addr_positional[25483:25480], addr_6370_7);

wire[31:0] addr_6371_7;

Selector_2 s6371_7(wires_1592_6[3], addr_1592_6, addr_positional[25487:25484], addr_6371_7);

wire[31:0] addr_6372_7;

Selector_2 s6372_7(wires_1593_6[0], addr_1593_6, addr_positional[25491:25488], addr_6372_7);

wire[31:0] addr_6373_7;

Selector_2 s6373_7(wires_1593_6[1], addr_1593_6, addr_positional[25495:25492], addr_6373_7);

wire[31:0] addr_6374_7;

Selector_2 s6374_7(wires_1593_6[2], addr_1593_6, addr_positional[25499:25496], addr_6374_7);

wire[31:0] addr_6375_7;

Selector_2 s6375_7(wires_1593_6[3], addr_1593_6, addr_positional[25503:25500], addr_6375_7);

wire[31:0] addr_6376_7;

Selector_2 s6376_7(wires_1594_6[0], addr_1594_6, addr_positional[25507:25504], addr_6376_7);

wire[31:0] addr_6377_7;

Selector_2 s6377_7(wires_1594_6[1], addr_1594_6, addr_positional[25511:25508], addr_6377_7);

wire[31:0] addr_6378_7;

Selector_2 s6378_7(wires_1594_6[2], addr_1594_6, addr_positional[25515:25512], addr_6378_7);

wire[31:0] addr_6379_7;

Selector_2 s6379_7(wires_1594_6[3], addr_1594_6, addr_positional[25519:25516], addr_6379_7);

wire[31:0] addr_6380_7;

Selector_2 s6380_7(wires_1595_6[0], addr_1595_6, addr_positional[25523:25520], addr_6380_7);

wire[31:0] addr_6381_7;

Selector_2 s6381_7(wires_1595_6[1], addr_1595_6, addr_positional[25527:25524], addr_6381_7);

wire[31:0] addr_6382_7;

Selector_2 s6382_7(wires_1595_6[2], addr_1595_6, addr_positional[25531:25528], addr_6382_7);

wire[31:0] addr_6383_7;

Selector_2 s6383_7(wires_1595_6[3], addr_1595_6, addr_positional[25535:25532], addr_6383_7);

wire[31:0] addr_6384_7;

Selector_2 s6384_7(wires_1596_6[0], addr_1596_6, addr_positional[25539:25536], addr_6384_7);

wire[31:0] addr_6385_7;

Selector_2 s6385_7(wires_1596_6[1], addr_1596_6, addr_positional[25543:25540], addr_6385_7);

wire[31:0] addr_6386_7;

Selector_2 s6386_7(wires_1596_6[2], addr_1596_6, addr_positional[25547:25544], addr_6386_7);

wire[31:0] addr_6387_7;

Selector_2 s6387_7(wires_1596_6[3], addr_1596_6, addr_positional[25551:25548], addr_6387_7);

wire[31:0] addr_6388_7;

Selector_2 s6388_7(wires_1597_6[0], addr_1597_6, addr_positional[25555:25552], addr_6388_7);

wire[31:0] addr_6389_7;

Selector_2 s6389_7(wires_1597_6[1], addr_1597_6, addr_positional[25559:25556], addr_6389_7);

wire[31:0] addr_6390_7;

Selector_2 s6390_7(wires_1597_6[2], addr_1597_6, addr_positional[25563:25560], addr_6390_7);

wire[31:0] addr_6391_7;

Selector_2 s6391_7(wires_1597_6[3], addr_1597_6, addr_positional[25567:25564], addr_6391_7);

wire[31:0] addr_6392_7;

Selector_2 s6392_7(wires_1598_6[0], addr_1598_6, addr_positional[25571:25568], addr_6392_7);

wire[31:0] addr_6393_7;

Selector_2 s6393_7(wires_1598_6[1], addr_1598_6, addr_positional[25575:25572], addr_6393_7);

wire[31:0] addr_6394_7;

Selector_2 s6394_7(wires_1598_6[2], addr_1598_6, addr_positional[25579:25576], addr_6394_7);

wire[31:0] addr_6395_7;

Selector_2 s6395_7(wires_1598_6[3], addr_1598_6, addr_positional[25583:25580], addr_6395_7);

wire[31:0] addr_6396_7;

Selector_2 s6396_7(wires_1599_6[0], addr_1599_6, addr_positional[25587:25584], addr_6396_7);

wire[31:0] addr_6397_7;

Selector_2 s6397_7(wires_1599_6[1], addr_1599_6, addr_positional[25591:25588], addr_6397_7);

wire[31:0] addr_6398_7;

Selector_2 s6398_7(wires_1599_6[2], addr_1599_6, addr_positional[25595:25592], addr_6398_7);

wire[31:0] addr_6399_7;

Selector_2 s6399_7(wires_1599_6[3], addr_1599_6, addr_positional[25599:25596], addr_6399_7);

wire[31:0] addr_6400_7;

Selector_2 s6400_7(wires_1600_6[0], addr_1600_6, addr_positional[25603:25600], addr_6400_7);

wire[31:0] addr_6401_7;

Selector_2 s6401_7(wires_1600_6[1], addr_1600_6, addr_positional[25607:25604], addr_6401_7);

wire[31:0] addr_6402_7;

Selector_2 s6402_7(wires_1600_6[2], addr_1600_6, addr_positional[25611:25608], addr_6402_7);

wire[31:0] addr_6403_7;

Selector_2 s6403_7(wires_1600_6[3], addr_1600_6, addr_positional[25615:25612], addr_6403_7);

wire[31:0] addr_6404_7;

Selector_2 s6404_7(wires_1601_6[0], addr_1601_6, addr_positional[25619:25616], addr_6404_7);

wire[31:0] addr_6405_7;

Selector_2 s6405_7(wires_1601_6[1], addr_1601_6, addr_positional[25623:25620], addr_6405_7);

wire[31:0] addr_6406_7;

Selector_2 s6406_7(wires_1601_6[2], addr_1601_6, addr_positional[25627:25624], addr_6406_7);

wire[31:0] addr_6407_7;

Selector_2 s6407_7(wires_1601_6[3], addr_1601_6, addr_positional[25631:25628], addr_6407_7);

wire[31:0] addr_6408_7;

Selector_2 s6408_7(wires_1602_6[0], addr_1602_6, addr_positional[25635:25632], addr_6408_7);

wire[31:0] addr_6409_7;

Selector_2 s6409_7(wires_1602_6[1], addr_1602_6, addr_positional[25639:25636], addr_6409_7);

wire[31:0] addr_6410_7;

Selector_2 s6410_7(wires_1602_6[2], addr_1602_6, addr_positional[25643:25640], addr_6410_7);

wire[31:0] addr_6411_7;

Selector_2 s6411_7(wires_1602_6[3], addr_1602_6, addr_positional[25647:25644], addr_6411_7);

wire[31:0] addr_6412_7;

Selector_2 s6412_7(wires_1603_6[0], addr_1603_6, addr_positional[25651:25648], addr_6412_7);

wire[31:0] addr_6413_7;

Selector_2 s6413_7(wires_1603_6[1], addr_1603_6, addr_positional[25655:25652], addr_6413_7);

wire[31:0] addr_6414_7;

Selector_2 s6414_7(wires_1603_6[2], addr_1603_6, addr_positional[25659:25656], addr_6414_7);

wire[31:0] addr_6415_7;

Selector_2 s6415_7(wires_1603_6[3], addr_1603_6, addr_positional[25663:25660], addr_6415_7);

wire[31:0] addr_6416_7;

Selector_2 s6416_7(wires_1604_6[0], addr_1604_6, addr_positional[25667:25664], addr_6416_7);

wire[31:0] addr_6417_7;

Selector_2 s6417_7(wires_1604_6[1], addr_1604_6, addr_positional[25671:25668], addr_6417_7);

wire[31:0] addr_6418_7;

Selector_2 s6418_7(wires_1604_6[2], addr_1604_6, addr_positional[25675:25672], addr_6418_7);

wire[31:0] addr_6419_7;

Selector_2 s6419_7(wires_1604_6[3], addr_1604_6, addr_positional[25679:25676], addr_6419_7);

wire[31:0] addr_6420_7;

Selector_2 s6420_7(wires_1605_6[0], addr_1605_6, addr_positional[25683:25680], addr_6420_7);

wire[31:0] addr_6421_7;

Selector_2 s6421_7(wires_1605_6[1], addr_1605_6, addr_positional[25687:25684], addr_6421_7);

wire[31:0] addr_6422_7;

Selector_2 s6422_7(wires_1605_6[2], addr_1605_6, addr_positional[25691:25688], addr_6422_7);

wire[31:0] addr_6423_7;

Selector_2 s6423_7(wires_1605_6[3], addr_1605_6, addr_positional[25695:25692], addr_6423_7);

wire[31:0] addr_6424_7;

Selector_2 s6424_7(wires_1606_6[0], addr_1606_6, addr_positional[25699:25696], addr_6424_7);

wire[31:0] addr_6425_7;

Selector_2 s6425_7(wires_1606_6[1], addr_1606_6, addr_positional[25703:25700], addr_6425_7);

wire[31:0] addr_6426_7;

Selector_2 s6426_7(wires_1606_6[2], addr_1606_6, addr_positional[25707:25704], addr_6426_7);

wire[31:0] addr_6427_7;

Selector_2 s6427_7(wires_1606_6[3], addr_1606_6, addr_positional[25711:25708], addr_6427_7);

wire[31:0] addr_6428_7;

Selector_2 s6428_7(wires_1607_6[0], addr_1607_6, addr_positional[25715:25712], addr_6428_7);

wire[31:0] addr_6429_7;

Selector_2 s6429_7(wires_1607_6[1], addr_1607_6, addr_positional[25719:25716], addr_6429_7);

wire[31:0] addr_6430_7;

Selector_2 s6430_7(wires_1607_6[2], addr_1607_6, addr_positional[25723:25720], addr_6430_7);

wire[31:0] addr_6431_7;

Selector_2 s6431_7(wires_1607_6[3], addr_1607_6, addr_positional[25727:25724], addr_6431_7);

wire[31:0] addr_6432_7;

Selector_2 s6432_7(wires_1608_6[0], addr_1608_6, addr_positional[25731:25728], addr_6432_7);

wire[31:0] addr_6433_7;

Selector_2 s6433_7(wires_1608_6[1], addr_1608_6, addr_positional[25735:25732], addr_6433_7);

wire[31:0] addr_6434_7;

Selector_2 s6434_7(wires_1608_6[2], addr_1608_6, addr_positional[25739:25736], addr_6434_7);

wire[31:0] addr_6435_7;

Selector_2 s6435_7(wires_1608_6[3], addr_1608_6, addr_positional[25743:25740], addr_6435_7);

wire[31:0] addr_6436_7;

Selector_2 s6436_7(wires_1609_6[0], addr_1609_6, addr_positional[25747:25744], addr_6436_7);

wire[31:0] addr_6437_7;

Selector_2 s6437_7(wires_1609_6[1], addr_1609_6, addr_positional[25751:25748], addr_6437_7);

wire[31:0] addr_6438_7;

Selector_2 s6438_7(wires_1609_6[2], addr_1609_6, addr_positional[25755:25752], addr_6438_7);

wire[31:0] addr_6439_7;

Selector_2 s6439_7(wires_1609_6[3], addr_1609_6, addr_positional[25759:25756], addr_6439_7);

wire[31:0] addr_6440_7;

Selector_2 s6440_7(wires_1610_6[0], addr_1610_6, addr_positional[25763:25760], addr_6440_7);

wire[31:0] addr_6441_7;

Selector_2 s6441_7(wires_1610_6[1], addr_1610_6, addr_positional[25767:25764], addr_6441_7);

wire[31:0] addr_6442_7;

Selector_2 s6442_7(wires_1610_6[2], addr_1610_6, addr_positional[25771:25768], addr_6442_7);

wire[31:0] addr_6443_7;

Selector_2 s6443_7(wires_1610_6[3], addr_1610_6, addr_positional[25775:25772], addr_6443_7);

wire[31:0] addr_6444_7;

Selector_2 s6444_7(wires_1611_6[0], addr_1611_6, addr_positional[25779:25776], addr_6444_7);

wire[31:0] addr_6445_7;

Selector_2 s6445_7(wires_1611_6[1], addr_1611_6, addr_positional[25783:25780], addr_6445_7);

wire[31:0] addr_6446_7;

Selector_2 s6446_7(wires_1611_6[2], addr_1611_6, addr_positional[25787:25784], addr_6446_7);

wire[31:0] addr_6447_7;

Selector_2 s6447_7(wires_1611_6[3], addr_1611_6, addr_positional[25791:25788], addr_6447_7);

wire[31:0] addr_6448_7;

Selector_2 s6448_7(wires_1612_6[0], addr_1612_6, addr_positional[25795:25792], addr_6448_7);

wire[31:0] addr_6449_7;

Selector_2 s6449_7(wires_1612_6[1], addr_1612_6, addr_positional[25799:25796], addr_6449_7);

wire[31:0] addr_6450_7;

Selector_2 s6450_7(wires_1612_6[2], addr_1612_6, addr_positional[25803:25800], addr_6450_7);

wire[31:0] addr_6451_7;

Selector_2 s6451_7(wires_1612_6[3], addr_1612_6, addr_positional[25807:25804], addr_6451_7);

wire[31:0] addr_6452_7;

Selector_2 s6452_7(wires_1613_6[0], addr_1613_6, addr_positional[25811:25808], addr_6452_7);

wire[31:0] addr_6453_7;

Selector_2 s6453_7(wires_1613_6[1], addr_1613_6, addr_positional[25815:25812], addr_6453_7);

wire[31:0] addr_6454_7;

Selector_2 s6454_7(wires_1613_6[2], addr_1613_6, addr_positional[25819:25816], addr_6454_7);

wire[31:0] addr_6455_7;

Selector_2 s6455_7(wires_1613_6[3], addr_1613_6, addr_positional[25823:25820], addr_6455_7);

wire[31:0] addr_6456_7;

Selector_2 s6456_7(wires_1614_6[0], addr_1614_6, addr_positional[25827:25824], addr_6456_7);

wire[31:0] addr_6457_7;

Selector_2 s6457_7(wires_1614_6[1], addr_1614_6, addr_positional[25831:25828], addr_6457_7);

wire[31:0] addr_6458_7;

Selector_2 s6458_7(wires_1614_6[2], addr_1614_6, addr_positional[25835:25832], addr_6458_7);

wire[31:0] addr_6459_7;

Selector_2 s6459_7(wires_1614_6[3], addr_1614_6, addr_positional[25839:25836], addr_6459_7);

wire[31:0] addr_6460_7;

Selector_2 s6460_7(wires_1615_6[0], addr_1615_6, addr_positional[25843:25840], addr_6460_7);

wire[31:0] addr_6461_7;

Selector_2 s6461_7(wires_1615_6[1], addr_1615_6, addr_positional[25847:25844], addr_6461_7);

wire[31:0] addr_6462_7;

Selector_2 s6462_7(wires_1615_6[2], addr_1615_6, addr_positional[25851:25848], addr_6462_7);

wire[31:0] addr_6463_7;

Selector_2 s6463_7(wires_1615_6[3], addr_1615_6, addr_positional[25855:25852], addr_6463_7);

wire[31:0] addr_6464_7;

Selector_2 s6464_7(wires_1616_6[0], addr_1616_6, addr_positional[25859:25856], addr_6464_7);

wire[31:0] addr_6465_7;

Selector_2 s6465_7(wires_1616_6[1], addr_1616_6, addr_positional[25863:25860], addr_6465_7);

wire[31:0] addr_6466_7;

Selector_2 s6466_7(wires_1616_6[2], addr_1616_6, addr_positional[25867:25864], addr_6466_7);

wire[31:0] addr_6467_7;

Selector_2 s6467_7(wires_1616_6[3], addr_1616_6, addr_positional[25871:25868], addr_6467_7);

wire[31:0] addr_6468_7;

Selector_2 s6468_7(wires_1617_6[0], addr_1617_6, addr_positional[25875:25872], addr_6468_7);

wire[31:0] addr_6469_7;

Selector_2 s6469_7(wires_1617_6[1], addr_1617_6, addr_positional[25879:25876], addr_6469_7);

wire[31:0] addr_6470_7;

Selector_2 s6470_7(wires_1617_6[2], addr_1617_6, addr_positional[25883:25880], addr_6470_7);

wire[31:0] addr_6471_7;

Selector_2 s6471_7(wires_1617_6[3], addr_1617_6, addr_positional[25887:25884], addr_6471_7);

wire[31:0] addr_6472_7;

Selector_2 s6472_7(wires_1618_6[0], addr_1618_6, addr_positional[25891:25888], addr_6472_7);

wire[31:0] addr_6473_7;

Selector_2 s6473_7(wires_1618_6[1], addr_1618_6, addr_positional[25895:25892], addr_6473_7);

wire[31:0] addr_6474_7;

Selector_2 s6474_7(wires_1618_6[2], addr_1618_6, addr_positional[25899:25896], addr_6474_7);

wire[31:0] addr_6475_7;

Selector_2 s6475_7(wires_1618_6[3], addr_1618_6, addr_positional[25903:25900], addr_6475_7);

wire[31:0] addr_6476_7;

Selector_2 s6476_7(wires_1619_6[0], addr_1619_6, addr_positional[25907:25904], addr_6476_7);

wire[31:0] addr_6477_7;

Selector_2 s6477_7(wires_1619_6[1], addr_1619_6, addr_positional[25911:25908], addr_6477_7);

wire[31:0] addr_6478_7;

Selector_2 s6478_7(wires_1619_6[2], addr_1619_6, addr_positional[25915:25912], addr_6478_7);

wire[31:0] addr_6479_7;

Selector_2 s6479_7(wires_1619_6[3], addr_1619_6, addr_positional[25919:25916], addr_6479_7);

wire[31:0] addr_6480_7;

Selector_2 s6480_7(wires_1620_6[0], addr_1620_6, addr_positional[25923:25920], addr_6480_7);

wire[31:0] addr_6481_7;

Selector_2 s6481_7(wires_1620_6[1], addr_1620_6, addr_positional[25927:25924], addr_6481_7);

wire[31:0] addr_6482_7;

Selector_2 s6482_7(wires_1620_6[2], addr_1620_6, addr_positional[25931:25928], addr_6482_7);

wire[31:0] addr_6483_7;

Selector_2 s6483_7(wires_1620_6[3], addr_1620_6, addr_positional[25935:25932], addr_6483_7);

wire[31:0] addr_6484_7;

Selector_2 s6484_7(wires_1621_6[0], addr_1621_6, addr_positional[25939:25936], addr_6484_7);

wire[31:0] addr_6485_7;

Selector_2 s6485_7(wires_1621_6[1], addr_1621_6, addr_positional[25943:25940], addr_6485_7);

wire[31:0] addr_6486_7;

Selector_2 s6486_7(wires_1621_6[2], addr_1621_6, addr_positional[25947:25944], addr_6486_7);

wire[31:0] addr_6487_7;

Selector_2 s6487_7(wires_1621_6[3], addr_1621_6, addr_positional[25951:25948], addr_6487_7);

wire[31:0] addr_6488_7;

Selector_2 s6488_7(wires_1622_6[0], addr_1622_6, addr_positional[25955:25952], addr_6488_7);

wire[31:0] addr_6489_7;

Selector_2 s6489_7(wires_1622_6[1], addr_1622_6, addr_positional[25959:25956], addr_6489_7);

wire[31:0] addr_6490_7;

Selector_2 s6490_7(wires_1622_6[2], addr_1622_6, addr_positional[25963:25960], addr_6490_7);

wire[31:0] addr_6491_7;

Selector_2 s6491_7(wires_1622_6[3], addr_1622_6, addr_positional[25967:25964], addr_6491_7);

wire[31:0] addr_6492_7;

Selector_2 s6492_7(wires_1623_6[0], addr_1623_6, addr_positional[25971:25968], addr_6492_7);

wire[31:0] addr_6493_7;

Selector_2 s6493_7(wires_1623_6[1], addr_1623_6, addr_positional[25975:25972], addr_6493_7);

wire[31:0] addr_6494_7;

Selector_2 s6494_7(wires_1623_6[2], addr_1623_6, addr_positional[25979:25976], addr_6494_7);

wire[31:0] addr_6495_7;

Selector_2 s6495_7(wires_1623_6[3], addr_1623_6, addr_positional[25983:25980], addr_6495_7);

wire[31:0] addr_6496_7;

Selector_2 s6496_7(wires_1624_6[0], addr_1624_6, addr_positional[25987:25984], addr_6496_7);

wire[31:0] addr_6497_7;

Selector_2 s6497_7(wires_1624_6[1], addr_1624_6, addr_positional[25991:25988], addr_6497_7);

wire[31:0] addr_6498_7;

Selector_2 s6498_7(wires_1624_6[2], addr_1624_6, addr_positional[25995:25992], addr_6498_7);

wire[31:0] addr_6499_7;

Selector_2 s6499_7(wires_1624_6[3], addr_1624_6, addr_positional[25999:25996], addr_6499_7);

wire[31:0] addr_6500_7;

Selector_2 s6500_7(wires_1625_6[0], addr_1625_6, addr_positional[26003:26000], addr_6500_7);

wire[31:0] addr_6501_7;

Selector_2 s6501_7(wires_1625_6[1], addr_1625_6, addr_positional[26007:26004], addr_6501_7);

wire[31:0] addr_6502_7;

Selector_2 s6502_7(wires_1625_6[2], addr_1625_6, addr_positional[26011:26008], addr_6502_7);

wire[31:0] addr_6503_7;

Selector_2 s6503_7(wires_1625_6[3], addr_1625_6, addr_positional[26015:26012], addr_6503_7);

wire[31:0] addr_6504_7;

Selector_2 s6504_7(wires_1626_6[0], addr_1626_6, addr_positional[26019:26016], addr_6504_7);

wire[31:0] addr_6505_7;

Selector_2 s6505_7(wires_1626_6[1], addr_1626_6, addr_positional[26023:26020], addr_6505_7);

wire[31:0] addr_6506_7;

Selector_2 s6506_7(wires_1626_6[2], addr_1626_6, addr_positional[26027:26024], addr_6506_7);

wire[31:0] addr_6507_7;

Selector_2 s6507_7(wires_1626_6[3], addr_1626_6, addr_positional[26031:26028], addr_6507_7);

wire[31:0] addr_6508_7;

Selector_2 s6508_7(wires_1627_6[0], addr_1627_6, addr_positional[26035:26032], addr_6508_7);

wire[31:0] addr_6509_7;

Selector_2 s6509_7(wires_1627_6[1], addr_1627_6, addr_positional[26039:26036], addr_6509_7);

wire[31:0] addr_6510_7;

Selector_2 s6510_7(wires_1627_6[2], addr_1627_6, addr_positional[26043:26040], addr_6510_7);

wire[31:0] addr_6511_7;

Selector_2 s6511_7(wires_1627_6[3], addr_1627_6, addr_positional[26047:26044], addr_6511_7);

wire[31:0] addr_6512_7;

Selector_2 s6512_7(wires_1628_6[0], addr_1628_6, addr_positional[26051:26048], addr_6512_7);

wire[31:0] addr_6513_7;

Selector_2 s6513_7(wires_1628_6[1], addr_1628_6, addr_positional[26055:26052], addr_6513_7);

wire[31:0] addr_6514_7;

Selector_2 s6514_7(wires_1628_6[2], addr_1628_6, addr_positional[26059:26056], addr_6514_7);

wire[31:0] addr_6515_7;

Selector_2 s6515_7(wires_1628_6[3], addr_1628_6, addr_positional[26063:26060], addr_6515_7);

wire[31:0] addr_6516_7;

Selector_2 s6516_7(wires_1629_6[0], addr_1629_6, addr_positional[26067:26064], addr_6516_7);

wire[31:0] addr_6517_7;

Selector_2 s6517_7(wires_1629_6[1], addr_1629_6, addr_positional[26071:26068], addr_6517_7);

wire[31:0] addr_6518_7;

Selector_2 s6518_7(wires_1629_6[2], addr_1629_6, addr_positional[26075:26072], addr_6518_7);

wire[31:0] addr_6519_7;

Selector_2 s6519_7(wires_1629_6[3], addr_1629_6, addr_positional[26079:26076], addr_6519_7);

wire[31:0] addr_6520_7;

Selector_2 s6520_7(wires_1630_6[0], addr_1630_6, addr_positional[26083:26080], addr_6520_7);

wire[31:0] addr_6521_7;

Selector_2 s6521_7(wires_1630_6[1], addr_1630_6, addr_positional[26087:26084], addr_6521_7);

wire[31:0] addr_6522_7;

Selector_2 s6522_7(wires_1630_6[2], addr_1630_6, addr_positional[26091:26088], addr_6522_7);

wire[31:0] addr_6523_7;

Selector_2 s6523_7(wires_1630_6[3], addr_1630_6, addr_positional[26095:26092], addr_6523_7);

wire[31:0] addr_6524_7;

Selector_2 s6524_7(wires_1631_6[0], addr_1631_6, addr_positional[26099:26096], addr_6524_7);

wire[31:0] addr_6525_7;

Selector_2 s6525_7(wires_1631_6[1], addr_1631_6, addr_positional[26103:26100], addr_6525_7);

wire[31:0] addr_6526_7;

Selector_2 s6526_7(wires_1631_6[2], addr_1631_6, addr_positional[26107:26104], addr_6526_7);

wire[31:0] addr_6527_7;

Selector_2 s6527_7(wires_1631_6[3], addr_1631_6, addr_positional[26111:26108], addr_6527_7);

wire[31:0] addr_6528_7;

Selector_2 s6528_7(wires_1632_6[0], addr_1632_6, addr_positional[26115:26112], addr_6528_7);

wire[31:0] addr_6529_7;

Selector_2 s6529_7(wires_1632_6[1], addr_1632_6, addr_positional[26119:26116], addr_6529_7);

wire[31:0] addr_6530_7;

Selector_2 s6530_7(wires_1632_6[2], addr_1632_6, addr_positional[26123:26120], addr_6530_7);

wire[31:0] addr_6531_7;

Selector_2 s6531_7(wires_1632_6[3], addr_1632_6, addr_positional[26127:26124], addr_6531_7);

wire[31:0] addr_6532_7;

Selector_2 s6532_7(wires_1633_6[0], addr_1633_6, addr_positional[26131:26128], addr_6532_7);

wire[31:0] addr_6533_7;

Selector_2 s6533_7(wires_1633_6[1], addr_1633_6, addr_positional[26135:26132], addr_6533_7);

wire[31:0] addr_6534_7;

Selector_2 s6534_7(wires_1633_6[2], addr_1633_6, addr_positional[26139:26136], addr_6534_7);

wire[31:0] addr_6535_7;

Selector_2 s6535_7(wires_1633_6[3], addr_1633_6, addr_positional[26143:26140], addr_6535_7);

wire[31:0] addr_6536_7;

Selector_2 s6536_7(wires_1634_6[0], addr_1634_6, addr_positional[26147:26144], addr_6536_7);

wire[31:0] addr_6537_7;

Selector_2 s6537_7(wires_1634_6[1], addr_1634_6, addr_positional[26151:26148], addr_6537_7);

wire[31:0] addr_6538_7;

Selector_2 s6538_7(wires_1634_6[2], addr_1634_6, addr_positional[26155:26152], addr_6538_7);

wire[31:0] addr_6539_7;

Selector_2 s6539_7(wires_1634_6[3], addr_1634_6, addr_positional[26159:26156], addr_6539_7);

wire[31:0] addr_6540_7;

Selector_2 s6540_7(wires_1635_6[0], addr_1635_6, addr_positional[26163:26160], addr_6540_7);

wire[31:0] addr_6541_7;

Selector_2 s6541_7(wires_1635_6[1], addr_1635_6, addr_positional[26167:26164], addr_6541_7);

wire[31:0] addr_6542_7;

Selector_2 s6542_7(wires_1635_6[2], addr_1635_6, addr_positional[26171:26168], addr_6542_7);

wire[31:0] addr_6543_7;

Selector_2 s6543_7(wires_1635_6[3], addr_1635_6, addr_positional[26175:26172], addr_6543_7);

wire[31:0] addr_6544_7;

Selector_2 s6544_7(wires_1636_6[0], addr_1636_6, addr_positional[26179:26176], addr_6544_7);

wire[31:0] addr_6545_7;

Selector_2 s6545_7(wires_1636_6[1], addr_1636_6, addr_positional[26183:26180], addr_6545_7);

wire[31:0] addr_6546_7;

Selector_2 s6546_7(wires_1636_6[2], addr_1636_6, addr_positional[26187:26184], addr_6546_7);

wire[31:0] addr_6547_7;

Selector_2 s6547_7(wires_1636_6[3], addr_1636_6, addr_positional[26191:26188], addr_6547_7);

wire[31:0] addr_6548_7;

Selector_2 s6548_7(wires_1637_6[0], addr_1637_6, addr_positional[26195:26192], addr_6548_7);

wire[31:0] addr_6549_7;

Selector_2 s6549_7(wires_1637_6[1], addr_1637_6, addr_positional[26199:26196], addr_6549_7);

wire[31:0] addr_6550_7;

Selector_2 s6550_7(wires_1637_6[2], addr_1637_6, addr_positional[26203:26200], addr_6550_7);

wire[31:0] addr_6551_7;

Selector_2 s6551_7(wires_1637_6[3], addr_1637_6, addr_positional[26207:26204], addr_6551_7);

wire[31:0] addr_6552_7;

Selector_2 s6552_7(wires_1638_6[0], addr_1638_6, addr_positional[26211:26208], addr_6552_7);

wire[31:0] addr_6553_7;

Selector_2 s6553_7(wires_1638_6[1], addr_1638_6, addr_positional[26215:26212], addr_6553_7);

wire[31:0] addr_6554_7;

Selector_2 s6554_7(wires_1638_6[2], addr_1638_6, addr_positional[26219:26216], addr_6554_7);

wire[31:0] addr_6555_7;

Selector_2 s6555_7(wires_1638_6[3], addr_1638_6, addr_positional[26223:26220], addr_6555_7);

wire[31:0] addr_6556_7;

Selector_2 s6556_7(wires_1639_6[0], addr_1639_6, addr_positional[26227:26224], addr_6556_7);

wire[31:0] addr_6557_7;

Selector_2 s6557_7(wires_1639_6[1], addr_1639_6, addr_positional[26231:26228], addr_6557_7);

wire[31:0] addr_6558_7;

Selector_2 s6558_7(wires_1639_6[2], addr_1639_6, addr_positional[26235:26232], addr_6558_7);

wire[31:0] addr_6559_7;

Selector_2 s6559_7(wires_1639_6[3], addr_1639_6, addr_positional[26239:26236], addr_6559_7);

wire[31:0] addr_6560_7;

Selector_2 s6560_7(wires_1640_6[0], addr_1640_6, addr_positional[26243:26240], addr_6560_7);

wire[31:0] addr_6561_7;

Selector_2 s6561_7(wires_1640_6[1], addr_1640_6, addr_positional[26247:26244], addr_6561_7);

wire[31:0] addr_6562_7;

Selector_2 s6562_7(wires_1640_6[2], addr_1640_6, addr_positional[26251:26248], addr_6562_7);

wire[31:0] addr_6563_7;

Selector_2 s6563_7(wires_1640_6[3], addr_1640_6, addr_positional[26255:26252], addr_6563_7);

wire[31:0] addr_6564_7;

Selector_2 s6564_7(wires_1641_6[0], addr_1641_6, addr_positional[26259:26256], addr_6564_7);

wire[31:0] addr_6565_7;

Selector_2 s6565_7(wires_1641_6[1], addr_1641_6, addr_positional[26263:26260], addr_6565_7);

wire[31:0] addr_6566_7;

Selector_2 s6566_7(wires_1641_6[2], addr_1641_6, addr_positional[26267:26264], addr_6566_7);

wire[31:0] addr_6567_7;

Selector_2 s6567_7(wires_1641_6[3], addr_1641_6, addr_positional[26271:26268], addr_6567_7);

wire[31:0] addr_6568_7;

Selector_2 s6568_7(wires_1642_6[0], addr_1642_6, addr_positional[26275:26272], addr_6568_7);

wire[31:0] addr_6569_7;

Selector_2 s6569_7(wires_1642_6[1], addr_1642_6, addr_positional[26279:26276], addr_6569_7);

wire[31:0] addr_6570_7;

Selector_2 s6570_7(wires_1642_6[2], addr_1642_6, addr_positional[26283:26280], addr_6570_7);

wire[31:0] addr_6571_7;

Selector_2 s6571_7(wires_1642_6[3], addr_1642_6, addr_positional[26287:26284], addr_6571_7);

wire[31:0] addr_6572_7;

Selector_2 s6572_7(wires_1643_6[0], addr_1643_6, addr_positional[26291:26288], addr_6572_7);

wire[31:0] addr_6573_7;

Selector_2 s6573_7(wires_1643_6[1], addr_1643_6, addr_positional[26295:26292], addr_6573_7);

wire[31:0] addr_6574_7;

Selector_2 s6574_7(wires_1643_6[2], addr_1643_6, addr_positional[26299:26296], addr_6574_7);

wire[31:0] addr_6575_7;

Selector_2 s6575_7(wires_1643_6[3], addr_1643_6, addr_positional[26303:26300], addr_6575_7);

wire[31:0] addr_6576_7;

Selector_2 s6576_7(wires_1644_6[0], addr_1644_6, addr_positional[26307:26304], addr_6576_7);

wire[31:0] addr_6577_7;

Selector_2 s6577_7(wires_1644_6[1], addr_1644_6, addr_positional[26311:26308], addr_6577_7);

wire[31:0] addr_6578_7;

Selector_2 s6578_7(wires_1644_6[2], addr_1644_6, addr_positional[26315:26312], addr_6578_7);

wire[31:0] addr_6579_7;

Selector_2 s6579_7(wires_1644_6[3], addr_1644_6, addr_positional[26319:26316], addr_6579_7);

wire[31:0] addr_6580_7;

Selector_2 s6580_7(wires_1645_6[0], addr_1645_6, addr_positional[26323:26320], addr_6580_7);

wire[31:0] addr_6581_7;

Selector_2 s6581_7(wires_1645_6[1], addr_1645_6, addr_positional[26327:26324], addr_6581_7);

wire[31:0] addr_6582_7;

Selector_2 s6582_7(wires_1645_6[2], addr_1645_6, addr_positional[26331:26328], addr_6582_7);

wire[31:0] addr_6583_7;

Selector_2 s6583_7(wires_1645_6[3], addr_1645_6, addr_positional[26335:26332], addr_6583_7);

wire[31:0] addr_6584_7;

Selector_2 s6584_7(wires_1646_6[0], addr_1646_6, addr_positional[26339:26336], addr_6584_7);

wire[31:0] addr_6585_7;

Selector_2 s6585_7(wires_1646_6[1], addr_1646_6, addr_positional[26343:26340], addr_6585_7);

wire[31:0] addr_6586_7;

Selector_2 s6586_7(wires_1646_6[2], addr_1646_6, addr_positional[26347:26344], addr_6586_7);

wire[31:0] addr_6587_7;

Selector_2 s6587_7(wires_1646_6[3], addr_1646_6, addr_positional[26351:26348], addr_6587_7);

wire[31:0] addr_6588_7;

Selector_2 s6588_7(wires_1647_6[0], addr_1647_6, addr_positional[26355:26352], addr_6588_7);

wire[31:0] addr_6589_7;

Selector_2 s6589_7(wires_1647_6[1], addr_1647_6, addr_positional[26359:26356], addr_6589_7);

wire[31:0] addr_6590_7;

Selector_2 s6590_7(wires_1647_6[2], addr_1647_6, addr_positional[26363:26360], addr_6590_7);

wire[31:0] addr_6591_7;

Selector_2 s6591_7(wires_1647_6[3], addr_1647_6, addr_positional[26367:26364], addr_6591_7);

wire[31:0] addr_6592_7;

Selector_2 s6592_7(wires_1648_6[0], addr_1648_6, addr_positional[26371:26368], addr_6592_7);

wire[31:0] addr_6593_7;

Selector_2 s6593_7(wires_1648_6[1], addr_1648_6, addr_positional[26375:26372], addr_6593_7);

wire[31:0] addr_6594_7;

Selector_2 s6594_7(wires_1648_6[2], addr_1648_6, addr_positional[26379:26376], addr_6594_7);

wire[31:0] addr_6595_7;

Selector_2 s6595_7(wires_1648_6[3], addr_1648_6, addr_positional[26383:26380], addr_6595_7);

wire[31:0] addr_6596_7;

Selector_2 s6596_7(wires_1649_6[0], addr_1649_6, addr_positional[26387:26384], addr_6596_7);

wire[31:0] addr_6597_7;

Selector_2 s6597_7(wires_1649_6[1], addr_1649_6, addr_positional[26391:26388], addr_6597_7);

wire[31:0] addr_6598_7;

Selector_2 s6598_7(wires_1649_6[2], addr_1649_6, addr_positional[26395:26392], addr_6598_7);

wire[31:0] addr_6599_7;

Selector_2 s6599_7(wires_1649_6[3], addr_1649_6, addr_positional[26399:26396], addr_6599_7);

wire[31:0] addr_6600_7;

Selector_2 s6600_7(wires_1650_6[0], addr_1650_6, addr_positional[26403:26400], addr_6600_7);

wire[31:0] addr_6601_7;

Selector_2 s6601_7(wires_1650_6[1], addr_1650_6, addr_positional[26407:26404], addr_6601_7);

wire[31:0] addr_6602_7;

Selector_2 s6602_7(wires_1650_6[2], addr_1650_6, addr_positional[26411:26408], addr_6602_7);

wire[31:0] addr_6603_7;

Selector_2 s6603_7(wires_1650_6[3], addr_1650_6, addr_positional[26415:26412], addr_6603_7);

wire[31:0] addr_6604_7;

Selector_2 s6604_7(wires_1651_6[0], addr_1651_6, addr_positional[26419:26416], addr_6604_7);

wire[31:0] addr_6605_7;

Selector_2 s6605_7(wires_1651_6[1], addr_1651_6, addr_positional[26423:26420], addr_6605_7);

wire[31:0] addr_6606_7;

Selector_2 s6606_7(wires_1651_6[2], addr_1651_6, addr_positional[26427:26424], addr_6606_7);

wire[31:0] addr_6607_7;

Selector_2 s6607_7(wires_1651_6[3], addr_1651_6, addr_positional[26431:26428], addr_6607_7);

wire[31:0] addr_6608_7;

Selector_2 s6608_7(wires_1652_6[0], addr_1652_6, addr_positional[26435:26432], addr_6608_7);

wire[31:0] addr_6609_7;

Selector_2 s6609_7(wires_1652_6[1], addr_1652_6, addr_positional[26439:26436], addr_6609_7);

wire[31:0] addr_6610_7;

Selector_2 s6610_7(wires_1652_6[2], addr_1652_6, addr_positional[26443:26440], addr_6610_7);

wire[31:0] addr_6611_7;

Selector_2 s6611_7(wires_1652_6[3], addr_1652_6, addr_positional[26447:26444], addr_6611_7);

wire[31:0] addr_6612_7;

Selector_2 s6612_7(wires_1653_6[0], addr_1653_6, addr_positional[26451:26448], addr_6612_7);

wire[31:0] addr_6613_7;

Selector_2 s6613_7(wires_1653_6[1], addr_1653_6, addr_positional[26455:26452], addr_6613_7);

wire[31:0] addr_6614_7;

Selector_2 s6614_7(wires_1653_6[2], addr_1653_6, addr_positional[26459:26456], addr_6614_7);

wire[31:0] addr_6615_7;

Selector_2 s6615_7(wires_1653_6[3], addr_1653_6, addr_positional[26463:26460], addr_6615_7);

wire[31:0] addr_6616_7;

Selector_2 s6616_7(wires_1654_6[0], addr_1654_6, addr_positional[26467:26464], addr_6616_7);

wire[31:0] addr_6617_7;

Selector_2 s6617_7(wires_1654_6[1], addr_1654_6, addr_positional[26471:26468], addr_6617_7);

wire[31:0] addr_6618_7;

Selector_2 s6618_7(wires_1654_6[2], addr_1654_6, addr_positional[26475:26472], addr_6618_7);

wire[31:0] addr_6619_7;

Selector_2 s6619_7(wires_1654_6[3], addr_1654_6, addr_positional[26479:26476], addr_6619_7);

wire[31:0] addr_6620_7;

Selector_2 s6620_7(wires_1655_6[0], addr_1655_6, addr_positional[26483:26480], addr_6620_7);

wire[31:0] addr_6621_7;

Selector_2 s6621_7(wires_1655_6[1], addr_1655_6, addr_positional[26487:26484], addr_6621_7);

wire[31:0] addr_6622_7;

Selector_2 s6622_7(wires_1655_6[2], addr_1655_6, addr_positional[26491:26488], addr_6622_7);

wire[31:0] addr_6623_7;

Selector_2 s6623_7(wires_1655_6[3], addr_1655_6, addr_positional[26495:26492], addr_6623_7);

wire[31:0] addr_6624_7;

Selector_2 s6624_7(wires_1656_6[0], addr_1656_6, addr_positional[26499:26496], addr_6624_7);

wire[31:0] addr_6625_7;

Selector_2 s6625_7(wires_1656_6[1], addr_1656_6, addr_positional[26503:26500], addr_6625_7);

wire[31:0] addr_6626_7;

Selector_2 s6626_7(wires_1656_6[2], addr_1656_6, addr_positional[26507:26504], addr_6626_7);

wire[31:0] addr_6627_7;

Selector_2 s6627_7(wires_1656_6[3], addr_1656_6, addr_positional[26511:26508], addr_6627_7);

wire[31:0] addr_6628_7;

Selector_2 s6628_7(wires_1657_6[0], addr_1657_6, addr_positional[26515:26512], addr_6628_7);

wire[31:0] addr_6629_7;

Selector_2 s6629_7(wires_1657_6[1], addr_1657_6, addr_positional[26519:26516], addr_6629_7);

wire[31:0] addr_6630_7;

Selector_2 s6630_7(wires_1657_6[2], addr_1657_6, addr_positional[26523:26520], addr_6630_7);

wire[31:0] addr_6631_7;

Selector_2 s6631_7(wires_1657_6[3], addr_1657_6, addr_positional[26527:26524], addr_6631_7);

wire[31:0] addr_6632_7;

Selector_2 s6632_7(wires_1658_6[0], addr_1658_6, addr_positional[26531:26528], addr_6632_7);

wire[31:0] addr_6633_7;

Selector_2 s6633_7(wires_1658_6[1], addr_1658_6, addr_positional[26535:26532], addr_6633_7);

wire[31:0] addr_6634_7;

Selector_2 s6634_7(wires_1658_6[2], addr_1658_6, addr_positional[26539:26536], addr_6634_7);

wire[31:0] addr_6635_7;

Selector_2 s6635_7(wires_1658_6[3], addr_1658_6, addr_positional[26543:26540], addr_6635_7);

wire[31:0] addr_6636_7;

Selector_2 s6636_7(wires_1659_6[0], addr_1659_6, addr_positional[26547:26544], addr_6636_7);

wire[31:0] addr_6637_7;

Selector_2 s6637_7(wires_1659_6[1], addr_1659_6, addr_positional[26551:26548], addr_6637_7);

wire[31:0] addr_6638_7;

Selector_2 s6638_7(wires_1659_6[2], addr_1659_6, addr_positional[26555:26552], addr_6638_7);

wire[31:0] addr_6639_7;

Selector_2 s6639_7(wires_1659_6[3], addr_1659_6, addr_positional[26559:26556], addr_6639_7);

wire[31:0] addr_6640_7;

Selector_2 s6640_7(wires_1660_6[0], addr_1660_6, addr_positional[26563:26560], addr_6640_7);

wire[31:0] addr_6641_7;

Selector_2 s6641_7(wires_1660_6[1], addr_1660_6, addr_positional[26567:26564], addr_6641_7);

wire[31:0] addr_6642_7;

Selector_2 s6642_7(wires_1660_6[2], addr_1660_6, addr_positional[26571:26568], addr_6642_7);

wire[31:0] addr_6643_7;

Selector_2 s6643_7(wires_1660_6[3], addr_1660_6, addr_positional[26575:26572], addr_6643_7);

wire[31:0] addr_6644_7;

Selector_2 s6644_7(wires_1661_6[0], addr_1661_6, addr_positional[26579:26576], addr_6644_7);

wire[31:0] addr_6645_7;

Selector_2 s6645_7(wires_1661_6[1], addr_1661_6, addr_positional[26583:26580], addr_6645_7);

wire[31:0] addr_6646_7;

Selector_2 s6646_7(wires_1661_6[2], addr_1661_6, addr_positional[26587:26584], addr_6646_7);

wire[31:0] addr_6647_7;

Selector_2 s6647_7(wires_1661_6[3], addr_1661_6, addr_positional[26591:26588], addr_6647_7);

wire[31:0] addr_6648_7;

Selector_2 s6648_7(wires_1662_6[0], addr_1662_6, addr_positional[26595:26592], addr_6648_7);

wire[31:0] addr_6649_7;

Selector_2 s6649_7(wires_1662_6[1], addr_1662_6, addr_positional[26599:26596], addr_6649_7);

wire[31:0] addr_6650_7;

Selector_2 s6650_7(wires_1662_6[2], addr_1662_6, addr_positional[26603:26600], addr_6650_7);

wire[31:0] addr_6651_7;

Selector_2 s6651_7(wires_1662_6[3], addr_1662_6, addr_positional[26607:26604], addr_6651_7);

wire[31:0] addr_6652_7;

Selector_2 s6652_7(wires_1663_6[0], addr_1663_6, addr_positional[26611:26608], addr_6652_7);

wire[31:0] addr_6653_7;

Selector_2 s6653_7(wires_1663_6[1], addr_1663_6, addr_positional[26615:26612], addr_6653_7);

wire[31:0] addr_6654_7;

Selector_2 s6654_7(wires_1663_6[2], addr_1663_6, addr_positional[26619:26616], addr_6654_7);

wire[31:0] addr_6655_7;

Selector_2 s6655_7(wires_1663_6[3], addr_1663_6, addr_positional[26623:26620], addr_6655_7);

wire[31:0] addr_6656_7;

Selector_2 s6656_7(wires_1664_6[0], addr_1664_6, addr_positional[26627:26624], addr_6656_7);

wire[31:0] addr_6657_7;

Selector_2 s6657_7(wires_1664_6[1], addr_1664_6, addr_positional[26631:26628], addr_6657_7);

wire[31:0] addr_6658_7;

Selector_2 s6658_7(wires_1664_6[2], addr_1664_6, addr_positional[26635:26632], addr_6658_7);

wire[31:0] addr_6659_7;

Selector_2 s6659_7(wires_1664_6[3], addr_1664_6, addr_positional[26639:26636], addr_6659_7);

wire[31:0] addr_6660_7;

Selector_2 s6660_7(wires_1665_6[0], addr_1665_6, addr_positional[26643:26640], addr_6660_7);

wire[31:0] addr_6661_7;

Selector_2 s6661_7(wires_1665_6[1], addr_1665_6, addr_positional[26647:26644], addr_6661_7);

wire[31:0] addr_6662_7;

Selector_2 s6662_7(wires_1665_6[2], addr_1665_6, addr_positional[26651:26648], addr_6662_7);

wire[31:0] addr_6663_7;

Selector_2 s6663_7(wires_1665_6[3], addr_1665_6, addr_positional[26655:26652], addr_6663_7);

wire[31:0] addr_6664_7;

Selector_2 s6664_7(wires_1666_6[0], addr_1666_6, addr_positional[26659:26656], addr_6664_7);

wire[31:0] addr_6665_7;

Selector_2 s6665_7(wires_1666_6[1], addr_1666_6, addr_positional[26663:26660], addr_6665_7);

wire[31:0] addr_6666_7;

Selector_2 s6666_7(wires_1666_6[2], addr_1666_6, addr_positional[26667:26664], addr_6666_7);

wire[31:0] addr_6667_7;

Selector_2 s6667_7(wires_1666_6[3], addr_1666_6, addr_positional[26671:26668], addr_6667_7);

wire[31:0] addr_6668_7;

Selector_2 s6668_7(wires_1667_6[0], addr_1667_6, addr_positional[26675:26672], addr_6668_7);

wire[31:0] addr_6669_7;

Selector_2 s6669_7(wires_1667_6[1], addr_1667_6, addr_positional[26679:26676], addr_6669_7);

wire[31:0] addr_6670_7;

Selector_2 s6670_7(wires_1667_6[2], addr_1667_6, addr_positional[26683:26680], addr_6670_7);

wire[31:0] addr_6671_7;

Selector_2 s6671_7(wires_1667_6[3], addr_1667_6, addr_positional[26687:26684], addr_6671_7);

wire[31:0] addr_6672_7;

Selector_2 s6672_7(wires_1668_6[0], addr_1668_6, addr_positional[26691:26688], addr_6672_7);

wire[31:0] addr_6673_7;

Selector_2 s6673_7(wires_1668_6[1], addr_1668_6, addr_positional[26695:26692], addr_6673_7);

wire[31:0] addr_6674_7;

Selector_2 s6674_7(wires_1668_6[2], addr_1668_6, addr_positional[26699:26696], addr_6674_7);

wire[31:0] addr_6675_7;

Selector_2 s6675_7(wires_1668_6[3], addr_1668_6, addr_positional[26703:26700], addr_6675_7);

wire[31:0] addr_6676_7;

Selector_2 s6676_7(wires_1669_6[0], addr_1669_6, addr_positional[26707:26704], addr_6676_7);

wire[31:0] addr_6677_7;

Selector_2 s6677_7(wires_1669_6[1], addr_1669_6, addr_positional[26711:26708], addr_6677_7);

wire[31:0] addr_6678_7;

Selector_2 s6678_7(wires_1669_6[2], addr_1669_6, addr_positional[26715:26712], addr_6678_7);

wire[31:0] addr_6679_7;

Selector_2 s6679_7(wires_1669_6[3], addr_1669_6, addr_positional[26719:26716], addr_6679_7);

wire[31:0] addr_6680_7;

Selector_2 s6680_7(wires_1670_6[0], addr_1670_6, addr_positional[26723:26720], addr_6680_7);

wire[31:0] addr_6681_7;

Selector_2 s6681_7(wires_1670_6[1], addr_1670_6, addr_positional[26727:26724], addr_6681_7);

wire[31:0] addr_6682_7;

Selector_2 s6682_7(wires_1670_6[2], addr_1670_6, addr_positional[26731:26728], addr_6682_7);

wire[31:0] addr_6683_7;

Selector_2 s6683_7(wires_1670_6[3], addr_1670_6, addr_positional[26735:26732], addr_6683_7);

wire[31:0] addr_6684_7;

Selector_2 s6684_7(wires_1671_6[0], addr_1671_6, addr_positional[26739:26736], addr_6684_7);

wire[31:0] addr_6685_7;

Selector_2 s6685_7(wires_1671_6[1], addr_1671_6, addr_positional[26743:26740], addr_6685_7);

wire[31:0] addr_6686_7;

Selector_2 s6686_7(wires_1671_6[2], addr_1671_6, addr_positional[26747:26744], addr_6686_7);

wire[31:0] addr_6687_7;

Selector_2 s6687_7(wires_1671_6[3], addr_1671_6, addr_positional[26751:26748], addr_6687_7);

wire[31:0] addr_6688_7;

Selector_2 s6688_7(wires_1672_6[0], addr_1672_6, addr_positional[26755:26752], addr_6688_7);

wire[31:0] addr_6689_7;

Selector_2 s6689_7(wires_1672_6[1], addr_1672_6, addr_positional[26759:26756], addr_6689_7);

wire[31:0] addr_6690_7;

Selector_2 s6690_7(wires_1672_6[2], addr_1672_6, addr_positional[26763:26760], addr_6690_7);

wire[31:0] addr_6691_7;

Selector_2 s6691_7(wires_1672_6[3], addr_1672_6, addr_positional[26767:26764], addr_6691_7);

wire[31:0] addr_6692_7;

Selector_2 s6692_7(wires_1673_6[0], addr_1673_6, addr_positional[26771:26768], addr_6692_7);

wire[31:0] addr_6693_7;

Selector_2 s6693_7(wires_1673_6[1], addr_1673_6, addr_positional[26775:26772], addr_6693_7);

wire[31:0] addr_6694_7;

Selector_2 s6694_7(wires_1673_6[2], addr_1673_6, addr_positional[26779:26776], addr_6694_7);

wire[31:0] addr_6695_7;

Selector_2 s6695_7(wires_1673_6[3], addr_1673_6, addr_positional[26783:26780], addr_6695_7);

wire[31:0] addr_6696_7;

Selector_2 s6696_7(wires_1674_6[0], addr_1674_6, addr_positional[26787:26784], addr_6696_7);

wire[31:0] addr_6697_7;

Selector_2 s6697_7(wires_1674_6[1], addr_1674_6, addr_positional[26791:26788], addr_6697_7);

wire[31:0] addr_6698_7;

Selector_2 s6698_7(wires_1674_6[2], addr_1674_6, addr_positional[26795:26792], addr_6698_7);

wire[31:0] addr_6699_7;

Selector_2 s6699_7(wires_1674_6[3], addr_1674_6, addr_positional[26799:26796], addr_6699_7);

wire[31:0] addr_6700_7;

Selector_2 s6700_7(wires_1675_6[0], addr_1675_6, addr_positional[26803:26800], addr_6700_7);

wire[31:0] addr_6701_7;

Selector_2 s6701_7(wires_1675_6[1], addr_1675_6, addr_positional[26807:26804], addr_6701_7);

wire[31:0] addr_6702_7;

Selector_2 s6702_7(wires_1675_6[2], addr_1675_6, addr_positional[26811:26808], addr_6702_7);

wire[31:0] addr_6703_7;

Selector_2 s6703_7(wires_1675_6[3], addr_1675_6, addr_positional[26815:26812], addr_6703_7);

wire[31:0] addr_6704_7;

Selector_2 s6704_7(wires_1676_6[0], addr_1676_6, addr_positional[26819:26816], addr_6704_7);

wire[31:0] addr_6705_7;

Selector_2 s6705_7(wires_1676_6[1], addr_1676_6, addr_positional[26823:26820], addr_6705_7);

wire[31:0] addr_6706_7;

Selector_2 s6706_7(wires_1676_6[2], addr_1676_6, addr_positional[26827:26824], addr_6706_7);

wire[31:0] addr_6707_7;

Selector_2 s6707_7(wires_1676_6[3], addr_1676_6, addr_positional[26831:26828], addr_6707_7);

wire[31:0] addr_6708_7;

Selector_2 s6708_7(wires_1677_6[0], addr_1677_6, addr_positional[26835:26832], addr_6708_7);

wire[31:0] addr_6709_7;

Selector_2 s6709_7(wires_1677_6[1], addr_1677_6, addr_positional[26839:26836], addr_6709_7);

wire[31:0] addr_6710_7;

Selector_2 s6710_7(wires_1677_6[2], addr_1677_6, addr_positional[26843:26840], addr_6710_7);

wire[31:0] addr_6711_7;

Selector_2 s6711_7(wires_1677_6[3], addr_1677_6, addr_positional[26847:26844], addr_6711_7);

wire[31:0] addr_6712_7;

Selector_2 s6712_7(wires_1678_6[0], addr_1678_6, addr_positional[26851:26848], addr_6712_7);

wire[31:0] addr_6713_7;

Selector_2 s6713_7(wires_1678_6[1], addr_1678_6, addr_positional[26855:26852], addr_6713_7);

wire[31:0] addr_6714_7;

Selector_2 s6714_7(wires_1678_6[2], addr_1678_6, addr_positional[26859:26856], addr_6714_7);

wire[31:0] addr_6715_7;

Selector_2 s6715_7(wires_1678_6[3], addr_1678_6, addr_positional[26863:26860], addr_6715_7);

wire[31:0] addr_6716_7;

Selector_2 s6716_7(wires_1679_6[0], addr_1679_6, addr_positional[26867:26864], addr_6716_7);

wire[31:0] addr_6717_7;

Selector_2 s6717_7(wires_1679_6[1], addr_1679_6, addr_positional[26871:26868], addr_6717_7);

wire[31:0] addr_6718_7;

Selector_2 s6718_7(wires_1679_6[2], addr_1679_6, addr_positional[26875:26872], addr_6718_7);

wire[31:0] addr_6719_7;

Selector_2 s6719_7(wires_1679_6[3], addr_1679_6, addr_positional[26879:26876], addr_6719_7);

wire[31:0] addr_6720_7;

Selector_2 s6720_7(wires_1680_6[0], addr_1680_6, addr_positional[26883:26880], addr_6720_7);

wire[31:0] addr_6721_7;

Selector_2 s6721_7(wires_1680_6[1], addr_1680_6, addr_positional[26887:26884], addr_6721_7);

wire[31:0] addr_6722_7;

Selector_2 s6722_7(wires_1680_6[2], addr_1680_6, addr_positional[26891:26888], addr_6722_7);

wire[31:0] addr_6723_7;

Selector_2 s6723_7(wires_1680_6[3], addr_1680_6, addr_positional[26895:26892], addr_6723_7);

wire[31:0] addr_6724_7;

Selector_2 s6724_7(wires_1681_6[0], addr_1681_6, addr_positional[26899:26896], addr_6724_7);

wire[31:0] addr_6725_7;

Selector_2 s6725_7(wires_1681_6[1], addr_1681_6, addr_positional[26903:26900], addr_6725_7);

wire[31:0] addr_6726_7;

Selector_2 s6726_7(wires_1681_6[2], addr_1681_6, addr_positional[26907:26904], addr_6726_7);

wire[31:0] addr_6727_7;

Selector_2 s6727_7(wires_1681_6[3], addr_1681_6, addr_positional[26911:26908], addr_6727_7);

wire[31:0] addr_6728_7;

Selector_2 s6728_7(wires_1682_6[0], addr_1682_6, addr_positional[26915:26912], addr_6728_7);

wire[31:0] addr_6729_7;

Selector_2 s6729_7(wires_1682_6[1], addr_1682_6, addr_positional[26919:26916], addr_6729_7);

wire[31:0] addr_6730_7;

Selector_2 s6730_7(wires_1682_6[2], addr_1682_6, addr_positional[26923:26920], addr_6730_7);

wire[31:0] addr_6731_7;

Selector_2 s6731_7(wires_1682_6[3], addr_1682_6, addr_positional[26927:26924], addr_6731_7);

wire[31:0] addr_6732_7;

Selector_2 s6732_7(wires_1683_6[0], addr_1683_6, addr_positional[26931:26928], addr_6732_7);

wire[31:0] addr_6733_7;

Selector_2 s6733_7(wires_1683_6[1], addr_1683_6, addr_positional[26935:26932], addr_6733_7);

wire[31:0] addr_6734_7;

Selector_2 s6734_7(wires_1683_6[2], addr_1683_6, addr_positional[26939:26936], addr_6734_7);

wire[31:0] addr_6735_7;

Selector_2 s6735_7(wires_1683_6[3], addr_1683_6, addr_positional[26943:26940], addr_6735_7);

wire[31:0] addr_6736_7;

Selector_2 s6736_7(wires_1684_6[0], addr_1684_6, addr_positional[26947:26944], addr_6736_7);

wire[31:0] addr_6737_7;

Selector_2 s6737_7(wires_1684_6[1], addr_1684_6, addr_positional[26951:26948], addr_6737_7);

wire[31:0] addr_6738_7;

Selector_2 s6738_7(wires_1684_6[2], addr_1684_6, addr_positional[26955:26952], addr_6738_7);

wire[31:0] addr_6739_7;

Selector_2 s6739_7(wires_1684_6[3], addr_1684_6, addr_positional[26959:26956], addr_6739_7);

wire[31:0] addr_6740_7;

Selector_2 s6740_7(wires_1685_6[0], addr_1685_6, addr_positional[26963:26960], addr_6740_7);

wire[31:0] addr_6741_7;

Selector_2 s6741_7(wires_1685_6[1], addr_1685_6, addr_positional[26967:26964], addr_6741_7);

wire[31:0] addr_6742_7;

Selector_2 s6742_7(wires_1685_6[2], addr_1685_6, addr_positional[26971:26968], addr_6742_7);

wire[31:0] addr_6743_7;

Selector_2 s6743_7(wires_1685_6[3], addr_1685_6, addr_positional[26975:26972], addr_6743_7);

wire[31:0] addr_6744_7;

Selector_2 s6744_7(wires_1686_6[0], addr_1686_6, addr_positional[26979:26976], addr_6744_7);

wire[31:0] addr_6745_7;

Selector_2 s6745_7(wires_1686_6[1], addr_1686_6, addr_positional[26983:26980], addr_6745_7);

wire[31:0] addr_6746_7;

Selector_2 s6746_7(wires_1686_6[2], addr_1686_6, addr_positional[26987:26984], addr_6746_7);

wire[31:0] addr_6747_7;

Selector_2 s6747_7(wires_1686_6[3], addr_1686_6, addr_positional[26991:26988], addr_6747_7);

wire[31:0] addr_6748_7;

Selector_2 s6748_7(wires_1687_6[0], addr_1687_6, addr_positional[26995:26992], addr_6748_7);

wire[31:0] addr_6749_7;

Selector_2 s6749_7(wires_1687_6[1], addr_1687_6, addr_positional[26999:26996], addr_6749_7);

wire[31:0] addr_6750_7;

Selector_2 s6750_7(wires_1687_6[2], addr_1687_6, addr_positional[27003:27000], addr_6750_7);

wire[31:0] addr_6751_7;

Selector_2 s6751_7(wires_1687_6[3], addr_1687_6, addr_positional[27007:27004], addr_6751_7);

wire[31:0] addr_6752_7;

Selector_2 s6752_7(wires_1688_6[0], addr_1688_6, addr_positional[27011:27008], addr_6752_7);

wire[31:0] addr_6753_7;

Selector_2 s6753_7(wires_1688_6[1], addr_1688_6, addr_positional[27015:27012], addr_6753_7);

wire[31:0] addr_6754_7;

Selector_2 s6754_7(wires_1688_6[2], addr_1688_6, addr_positional[27019:27016], addr_6754_7);

wire[31:0] addr_6755_7;

Selector_2 s6755_7(wires_1688_6[3], addr_1688_6, addr_positional[27023:27020], addr_6755_7);

wire[31:0] addr_6756_7;

Selector_2 s6756_7(wires_1689_6[0], addr_1689_6, addr_positional[27027:27024], addr_6756_7);

wire[31:0] addr_6757_7;

Selector_2 s6757_7(wires_1689_6[1], addr_1689_6, addr_positional[27031:27028], addr_6757_7);

wire[31:0] addr_6758_7;

Selector_2 s6758_7(wires_1689_6[2], addr_1689_6, addr_positional[27035:27032], addr_6758_7);

wire[31:0] addr_6759_7;

Selector_2 s6759_7(wires_1689_6[3], addr_1689_6, addr_positional[27039:27036], addr_6759_7);

wire[31:0] addr_6760_7;

Selector_2 s6760_7(wires_1690_6[0], addr_1690_6, addr_positional[27043:27040], addr_6760_7);

wire[31:0] addr_6761_7;

Selector_2 s6761_7(wires_1690_6[1], addr_1690_6, addr_positional[27047:27044], addr_6761_7);

wire[31:0] addr_6762_7;

Selector_2 s6762_7(wires_1690_6[2], addr_1690_6, addr_positional[27051:27048], addr_6762_7);

wire[31:0] addr_6763_7;

Selector_2 s6763_7(wires_1690_6[3], addr_1690_6, addr_positional[27055:27052], addr_6763_7);

wire[31:0] addr_6764_7;

Selector_2 s6764_7(wires_1691_6[0], addr_1691_6, addr_positional[27059:27056], addr_6764_7);

wire[31:0] addr_6765_7;

Selector_2 s6765_7(wires_1691_6[1], addr_1691_6, addr_positional[27063:27060], addr_6765_7);

wire[31:0] addr_6766_7;

Selector_2 s6766_7(wires_1691_6[2], addr_1691_6, addr_positional[27067:27064], addr_6766_7);

wire[31:0] addr_6767_7;

Selector_2 s6767_7(wires_1691_6[3], addr_1691_6, addr_positional[27071:27068], addr_6767_7);

wire[31:0] addr_6768_7;

Selector_2 s6768_7(wires_1692_6[0], addr_1692_6, addr_positional[27075:27072], addr_6768_7);

wire[31:0] addr_6769_7;

Selector_2 s6769_7(wires_1692_6[1], addr_1692_6, addr_positional[27079:27076], addr_6769_7);

wire[31:0] addr_6770_7;

Selector_2 s6770_7(wires_1692_6[2], addr_1692_6, addr_positional[27083:27080], addr_6770_7);

wire[31:0] addr_6771_7;

Selector_2 s6771_7(wires_1692_6[3], addr_1692_6, addr_positional[27087:27084], addr_6771_7);

wire[31:0] addr_6772_7;

Selector_2 s6772_7(wires_1693_6[0], addr_1693_6, addr_positional[27091:27088], addr_6772_7);

wire[31:0] addr_6773_7;

Selector_2 s6773_7(wires_1693_6[1], addr_1693_6, addr_positional[27095:27092], addr_6773_7);

wire[31:0] addr_6774_7;

Selector_2 s6774_7(wires_1693_6[2], addr_1693_6, addr_positional[27099:27096], addr_6774_7);

wire[31:0] addr_6775_7;

Selector_2 s6775_7(wires_1693_6[3], addr_1693_6, addr_positional[27103:27100], addr_6775_7);

wire[31:0] addr_6776_7;

Selector_2 s6776_7(wires_1694_6[0], addr_1694_6, addr_positional[27107:27104], addr_6776_7);

wire[31:0] addr_6777_7;

Selector_2 s6777_7(wires_1694_6[1], addr_1694_6, addr_positional[27111:27108], addr_6777_7);

wire[31:0] addr_6778_7;

Selector_2 s6778_7(wires_1694_6[2], addr_1694_6, addr_positional[27115:27112], addr_6778_7);

wire[31:0] addr_6779_7;

Selector_2 s6779_7(wires_1694_6[3], addr_1694_6, addr_positional[27119:27116], addr_6779_7);

wire[31:0] addr_6780_7;

Selector_2 s6780_7(wires_1695_6[0], addr_1695_6, addr_positional[27123:27120], addr_6780_7);

wire[31:0] addr_6781_7;

Selector_2 s6781_7(wires_1695_6[1], addr_1695_6, addr_positional[27127:27124], addr_6781_7);

wire[31:0] addr_6782_7;

Selector_2 s6782_7(wires_1695_6[2], addr_1695_6, addr_positional[27131:27128], addr_6782_7);

wire[31:0] addr_6783_7;

Selector_2 s6783_7(wires_1695_6[3], addr_1695_6, addr_positional[27135:27132], addr_6783_7);

wire[31:0] addr_6784_7;

Selector_2 s6784_7(wires_1696_6[0], addr_1696_6, addr_positional[27139:27136], addr_6784_7);

wire[31:0] addr_6785_7;

Selector_2 s6785_7(wires_1696_6[1], addr_1696_6, addr_positional[27143:27140], addr_6785_7);

wire[31:0] addr_6786_7;

Selector_2 s6786_7(wires_1696_6[2], addr_1696_6, addr_positional[27147:27144], addr_6786_7);

wire[31:0] addr_6787_7;

Selector_2 s6787_7(wires_1696_6[3], addr_1696_6, addr_positional[27151:27148], addr_6787_7);

wire[31:0] addr_6788_7;

Selector_2 s6788_7(wires_1697_6[0], addr_1697_6, addr_positional[27155:27152], addr_6788_7);

wire[31:0] addr_6789_7;

Selector_2 s6789_7(wires_1697_6[1], addr_1697_6, addr_positional[27159:27156], addr_6789_7);

wire[31:0] addr_6790_7;

Selector_2 s6790_7(wires_1697_6[2], addr_1697_6, addr_positional[27163:27160], addr_6790_7);

wire[31:0] addr_6791_7;

Selector_2 s6791_7(wires_1697_6[3], addr_1697_6, addr_positional[27167:27164], addr_6791_7);

wire[31:0] addr_6792_7;

Selector_2 s6792_7(wires_1698_6[0], addr_1698_6, addr_positional[27171:27168], addr_6792_7);

wire[31:0] addr_6793_7;

Selector_2 s6793_7(wires_1698_6[1], addr_1698_6, addr_positional[27175:27172], addr_6793_7);

wire[31:0] addr_6794_7;

Selector_2 s6794_7(wires_1698_6[2], addr_1698_6, addr_positional[27179:27176], addr_6794_7);

wire[31:0] addr_6795_7;

Selector_2 s6795_7(wires_1698_6[3], addr_1698_6, addr_positional[27183:27180], addr_6795_7);

wire[31:0] addr_6796_7;

Selector_2 s6796_7(wires_1699_6[0], addr_1699_6, addr_positional[27187:27184], addr_6796_7);

wire[31:0] addr_6797_7;

Selector_2 s6797_7(wires_1699_6[1], addr_1699_6, addr_positional[27191:27188], addr_6797_7);

wire[31:0] addr_6798_7;

Selector_2 s6798_7(wires_1699_6[2], addr_1699_6, addr_positional[27195:27192], addr_6798_7);

wire[31:0] addr_6799_7;

Selector_2 s6799_7(wires_1699_6[3], addr_1699_6, addr_positional[27199:27196], addr_6799_7);

wire[31:0] addr_6800_7;

Selector_2 s6800_7(wires_1700_6[0], addr_1700_6, addr_positional[27203:27200], addr_6800_7);

wire[31:0] addr_6801_7;

Selector_2 s6801_7(wires_1700_6[1], addr_1700_6, addr_positional[27207:27204], addr_6801_7);

wire[31:0] addr_6802_7;

Selector_2 s6802_7(wires_1700_6[2], addr_1700_6, addr_positional[27211:27208], addr_6802_7);

wire[31:0] addr_6803_7;

Selector_2 s6803_7(wires_1700_6[3], addr_1700_6, addr_positional[27215:27212], addr_6803_7);

wire[31:0] addr_6804_7;

Selector_2 s6804_7(wires_1701_6[0], addr_1701_6, addr_positional[27219:27216], addr_6804_7);

wire[31:0] addr_6805_7;

Selector_2 s6805_7(wires_1701_6[1], addr_1701_6, addr_positional[27223:27220], addr_6805_7);

wire[31:0] addr_6806_7;

Selector_2 s6806_7(wires_1701_6[2], addr_1701_6, addr_positional[27227:27224], addr_6806_7);

wire[31:0] addr_6807_7;

Selector_2 s6807_7(wires_1701_6[3], addr_1701_6, addr_positional[27231:27228], addr_6807_7);

wire[31:0] addr_6808_7;

Selector_2 s6808_7(wires_1702_6[0], addr_1702_6, addr_positional[27235:27232], addr_6808_7);

wire[31:0] addr_6809_7;

Selector_2 s6809_7(wires_1702_6[1], addr_1702_6, addr_positional[27239:27236], addr_6809_7);

wire[31:0] addr_6810_7;

Selector_2 s6810_7(wires_1702_6[2], addr_1702_6, addr_positional[27243:27240], addr_6810_7);

wire[31:0] addr_6811_7;

Selector_2 s6811_7(wires_1702_6[3], addr_1702_6, addr_positional[27247:27244], addr_6811_7);

wire[31:0] addr_6812_7;

Selector_2 s6812_7(wires_1703_6[0], addr_1703_6, addr_positional[27251:27248], addr_6812_7);

wire[31:0] addr_6813_7;

Selector_2 s6813_7(wires_1703_6[1], addr_1703_6, addr_positional[27255:27252], addr_6813_7);

wire[31:0] addr_6814_7;

Selector_2 s6814_7(wires_1703_6[2], addr_1703_6, addr_positional[27259:27256], addr_6814_7);

wire[31:0] addr_6815_7;

Selector_2 s6815_7(wires_1703_6[3], addr_1703_6, addr_positional[27263:27260], addr_6815_7);

wire[31:0] addr_6816_7;

Selector_2 s6816_7(wires_1704_6[0], addr_1704_6, addr_positional[27267:27264], addr_6816_7);

wire[31:0] addr_6817_7;

Selector_2 s6817_7(wires_1704_6[1], addr_1704_6, addr_positional[27271:27268], addr_6817_7);

wire[31:0] addr_6818_7;

Selector_2 s6818_7(wires_1704_6[2], addr_1704_6, addr_positional[27275:27272], addr_6818_7);

wire[31:0] addr_6819_7;

Selector_2 s6819_7(wires_1704_6[3], addr_1704_6, addr_positional[27279:27276], addr_6819_7);

wire[31:0] addr_6820_7;

Selector_2 s6820_7(wires_1705_6[0], addr_1705_6, addr_positional[27283:27280], addr_6820_7);

wire[31:0] addr_6821_7;

Selector_2 s6821_7(wires_1705_6[1], addr_1705_6, addr_positional[27287:27284], addr_6821_7);

wire[31:0] addr_6822_7;

Selector_2 s6822_7(wires_1705_6[2], addr_1705_6, addr_positional[27291:27288], addr_6822_7);

wire[31:0] addr_6823_7;

Selector_2 s6823_7(wires_1705_6[3], addr_1705_6, addr_positional[27295:27292], addr_6823_7);

wire[31:0] addr_6824_7;

Selector_2 s6824_7(wires_1706_6[0], addr_1706_6, addr_positional[27299:27296], addr_6824_7);

wire[31:0] addr_6825_7;

Selector_2 s6825_7(wires_1706_6[1], addr_1706_6, addr_positional[27303:27300], addr_6825_7);

wire[31:0] addr_6826_7;

Selector_2 s6826_7(wires_1706_6[2], addr_1706_6, addr_positional[27307:27304], addr_6826_7);

wire[31:0] addr_6827_7;

Selector_2 s6827_7(wires_1706_6[3], addr_1706_6, addr_positional[27311:27308], addr_6827_7);

wire[31:0] addr_6828_7;

Selector_2 s6828_7(wires_1707_6[0], addr_1707_6, addr_positional[27315:27312], addr_6828_7);

wire[31:0] addr_6829_7;

Selector_2 s6829_7(wires_1707_6[1], addr_1707_6, addr_positional[27319:27316], addr_6829_7);

wire[31:0] addr_6830_7;

Selector_2 s6830_7(wires_1707_6[2], addr_1707_6, addr_positional[27323:27320], addr_6830_7);

wire[31:0] addr_6831_7;

Selector_2 s6831_7(wires_1707_6[3], addr_1707_6, addr_positional[27327:27324], addr_6831_7);

wire[31:0] addr_6832_7;

Selector_2 s6832_7(wires_1708_6[0], addr_1708_6, addr_positional[27331:27328], addr_6832_7);

wire[31:0] addr_6833_7;

Selector_2 s6833_7(wires_1708_6[1], addr_1708_6, addr_positional[27335:27332], addr_6833_7);

wire[31:0] addr_6834_7;

Selector_2 s6834_7(wires_1708_6[2], addr_1708_6, addr_positional[27339:27336], addr_6834_7);

wire[31:0] addr_6835_7;

Selector_2 s6835_7(wires_1708_6[3], addr_1708_6, addr_positional[27343:27340], addr_6835_7);

wire[31:0] addr_6836_7;

Selector_2 s6836_7(wires_1709_6[0], addr_1709_6, addr_positional[27347:27344], addr_6836_7);

wire[31:0] addr_6837_7;

Selector_2 s6837_7(wires_1709_6[1], addr_1709_6, addr_positional[27351:27348], addr_6837_7);

wire[31:0] addr_6838_7;

Selector_2 s6838_7(wires_1709_6[2], addr_1709_6, addr_positional[27355:27352], addr_6838_7);

wire[31:0] addr_6839_7;

Selector_2 s6839_7(wires_1709_6[3], addr_1709_6, addr_positional[27359:27356], addr_6839_7);

wire[31:0] addr_6840_7;

Selector_2 s6840_7(wires_1710_6[0], addr_1710_6, addr_positional[27363:27360], addr_6840_7);

wire[31:0] addr_6841_7;

Selector_2 s6841_7(wires_1710_6[1], addr_1710_6, addr_positional[27367:27364], addr_6841_7);

wire[31:0] addr_6842_7;

Selector_2 s6842_7(wires_1710_6[2], addr_1710_6, addr_positional[27371:27368], addr_6842_7);

wire[31:0] addr_6843_7;

Selector_2 s6843_7(wires_1710_6[3], addr_1710_6, addr_positional[27375:27372], addr_6843_7);

wire[31:0] addr_6844_7;

Selector_2 s6844_7(wires_1711_6[0], addr_1711_6, addr_positional[27379:27376], addr_6844_7);

wire[31:0] addr_6845_7;

Selector_2 s6845_7(wires_1711_6[1], addr_1711_6, addr_positional[27383:27380], addr_6845_7);

wire[31:0] addr_6846_7;

Selector_2 s6846_7(wires_1711_6[2], addr_1711_6, addr_positional[27387:27384], addr_6846_7);

wire[31:0] addr_6847_7;

Selector_2 s6847_7(wires_1711_6[3], addr_1711_6, addr_positional[27391:27388], addr_6847_7);

wire[31:0] addr_6848_7;

Selector_2 s6848_7(wires_1712_6[0], addr_1712_6, addr_positional[27395:27392], addr_6848_7);

wire[31:0] addr_6849_7;

Selector_2 s6849_7(wires_1712_6[1], addr_1712_6, addr_positional[27399:27396], addr_6849_7);

wire[31:0] addr_6850_7;

Selector_2 s6850_7(wires_1712_6[2], addr_1712_6, addr_positional[27403:27400], addr_6850_7);

wire[31:0] addr_6851_7;

Selector_2 s6851_7(wires_1712_6[3], addr_1712_6, addr_positional[27407:27404], addr_6851_7);

wire[31:0] addr_6852_7;

Selector_2 s6852_7(wires_1713_6[0], addr_1713_6, addr_positional[27411:27408], addr_6852_7);

wire[31:0] addr_6853_7;

Selector_2 s6853_7(wires_1713_6[1], addr_1713_6, addr_positional[27415:27412], addr_6853_7);

wire[31:0] addr_6854_7;

Selector_2 s6854_7(wires_1713_6[2], addr_1713_6, addr_positional[27419:27416], addr_6854_7);

wire[31:0] addr_6855_7;

Selector_2 s6855_7(wires_1713_6[3], addr_1713_6, addr_positional[27423:27420], addr_6855_7);

wire[31:0] addr_6856_7;

Selector_2 s6856_7(wires_1714_6[0], addr_1714_6, addr_positional[27427:27424], addr_6856_7);

wire[31:0] addr_6857_7;

Selector_2 s6857_7(wires_1714_6[1], addr_1714_6, addr_positional[27431:27428], addr_6857_7);

wire[31:0] addr_6858_7;

Selector_2 s6858_7(wires_1714_6[2], addr_1714_6, addr_positional[27435:27432], addr_6858_7);

wire[31:0] addr_6859_7;

Selector_2 s6859_7(wires_1714_6[3], addr_1714_6, addr_positional[27439:27436], addr_6859_7);

wire[31:0] addr_6860_7;

Selector_2 s6860_7(wires_1715_6[0], addr_1715_6, addr_positional[27443:27440], addr_6860_7);

wire[31:0] addr_6861_7;

Selector_2 s6861_7(wires_1715_6[1], addr_1715_6, addr_positional[27447:27444], addr_6861_7);

wire[31:0] addr_6862_7;

Selector_2 s6862_7(wires_1715_6[2], addr_1715_6, addr_positional[27451:27448], addr_6862_7);

wire[31:0] addr_6863_7;

Selector_2 s6863_7(wires_1715_6[3], addr_1715_6, addr_positional[27455:27452], addr_6863_7);

wire[31:0] addr_6864_7;

Selector_2 s6864_7(wires_1716_6[0], addr_1716_6, addr_positional[27459:27456], addr_6864_7);

wire[31:0] addr_6865_7;

Selector_2 s6865_7(wires_1716_6[1], addr_1716_6, addr_positional[27463:27460], addr_6865_7);

wire[31:0] addr_6866_7;

Selector_2 s6866_7(wires_1716_6[2], addr_1716_6, addr_positional[27467:27464], addr_6866_7);

wire[31:0] addr_6867_7;

Selector_2 s6867_7(wires_1716_6[3], addr_1716_6, addr_positional[27471:27468], addr_6867_7);

wire[31:0] addr_6868_7;

Selector_2 s6868_7(wires_1717_6[0], addr_1717_6, addr_positional[27475:27472], addr_6868_7);

wire[31:0] addr_6869_7;

Selector_2 s6869_7(wires_1717_6[1], addr_1717_6, addr_positional[27479:27476], addr_6869_7);

wire[31:0] addr_6870_7;

Selector_2 s6870_7(wires_1717_6[2], addr_1717_6, addr_positional[27483:27480], addr_6870_7);

wire[31:0] addr_6871_7;

Selector_2 s6871_7(wires_1717_6[3], addr_1717_6, addr_positional[27487:27484], addr_6871_7);

wire[31:0] addr_6872_7;

Selector_2 s6872_7(wires_1718_6[0], addr_1718_6, addr_positional[27491:27488], addr_6872_7);

wire[31:0] addr_6873_7;

Selector_2 s6873_7(wires_1718_6[1], addr_1718_6, addr_positional[27495:27492], addr_6873_7);

wire[31:0] addr_6874_7;

Selector_2 s6874_7(wires_1718_6[2], addr_1718_6, addr_positional[27499:27496], addr_6874_7);

wire[31:0] addr_6875_7;

Selector_2 s6875_7(wires_1718_6[3], addr_1718_6, addr_positional[27503:27500], addr_6875_7);

wire[31:0] addr_6876_7;

Selector_2 s6876_7(wires_1719_6[0], addr_1719_6, addr_positional[27507:27504], addr_6876_7);

wire[31:0] addr_6877_7;

Selector_2 s6877_7(wires_1719_6[1], addr_1719_6, addr_positional[27511:27508], addr_6877_7);

wire[31:0] addr_6878_7;

Selector_2 s6878_7(wires_1719_6[2], addr_1719_6, addr_positional[27515:27512], addr_6878_7);

wire[31:0] addr_6879_7;

Selector_2 s6879_7(wires_1719_6[3], addr_1719_6, addr_positional[27519:27516], addr_6879_7);

wire[31:0] addr_6880_7;

Selector_2 s6880_7(wires_1720_6[0], addr_1720_6, addr_positional[27523:27520], addr_6880_7);

wire[31:0] addr_6881_7;

Selector_2 s6881_7(wires_1720_6[1], addr_1720_6, addr_positional[27527:27524], addr_6881_7);

wire[31:0] addr_6882_7;

Selector_2 s6882_7(wires_1720_6[2], addr_1720_6, addr_positional[27531:27528], addr_6882_7);

wire[31:0] addr_6883_7;

Selector_2 s6883_7(wires_1720_6[3], addr_1720_6, addr_positional[27535:27532], addr_6883_7);

wire[31:0] addr_6884_7;

Selector_2 s6884_7(wires_1721_6[0], addr_1721_6, addr_positional[27539:27536], addr_6884_7);

wire[31:0] addr_6885_7;

Selector_2 s6885_7(wires_1721_6[1], addr_1721_6, addr_positional[27543:27540], addr_6885_7);

wire[31:0] addr_6886_7;

Selector_2 s6886_7(wires_1721_6[2], addr_1721_6, addr_positional[27547:27544], addr_6886_7);

wire[31:0] addr_6887_7;

Selector_2 s6887_7(wires_1721_6[3], addr_1721_6, addr_positional[27551:27548], addr_6887_7);

wire[31:0] addr_6888_7;

Selector_2 s6888_7(wires_1722_6[0], addr_1722_6, addr_positional[27555:27552], addr_6888_7);

wire[31:0] addr_6889_7;

Selector_2 s6889_7(wires_1722_6[1], addr_1722_6, addr_positional[27559:27556], addr_6889_7);

wire[31:0] addr_6890_7;

Selector_2 s6890_7(wires_1722_6[2], addr_1722_6, addr_positional[27563:27560], addr_6890_7);

wire[31:0] addr_6891_7;

Selector_2 s6891_7(wires_1722_6[3], addr_1722_6, addr_positional[27567:27564], addr_6891_7);

wire[31:0] addr_6892_7;

Selector_2 s6892_7(wires_1723_6[0], addr_1723_6, addr_positional[27571:27568], addr_6892_7);

wire[31:0] addr_6893_7;

Selector_2 s6893_7(wires_1723_6[1], addr_1723_6, addr_positional[27575:27572], addr_6893_7);

wire[31:0] addr_6894_7;

Selector_2 s6894_7(wires_1723_6[2], addr_1723_6, addr_positional[27579:27576], addr_6894_7);

wire[31:0] addr_6895_7;

Selector_2 s6895_7(wires_1723_6[3], addr_1723_6, addr_positional[27583:27580], addr_6895_7);

wire[31:0] addr_6896_7;

Selector_2 s6896_7(wires_1724_6[0], addr_1724_6, addr_positional[27587:27584], addr_6896_7);

wire[31:0] addr_6897_7;

Selector_2 s6897_7(wires_1724_6[1], addr_1724_6, addr_positional[27591:27588], addr_6897_7);

wire[31:0] addr_6898_7;

Selector_2 s6898_7(wires_1724_6[2], addr_1724_6, addr_positional[27595:27592], addr_6898_7);

wire[31:0] addr_6899_7;

Selector_2 s6899_7(wires_1724_6[3], addr_1724_6, addr_positional[27599:27596], addr_6899_7);

wire[31:0] addr_6900_7;

Selector_2 s6900_7(wires_1725_6[0], addr_1725_6, addr_positional[27603:27600], addr_6900_7);

wire[31:0] addr_6901_7;

Selector_2 s6901_7(wires_1725_6[1], addr_1725_6, addr_positional[27607:27604], addr_6901_7);

wire[31:0] addr_6902_7;

Selector_2 s6902_7(wires_1725_6[2], addr_1725_6, addr_positional[27611:27608], addr_6902_7);

wire[31:0] addr_6903_7;

Selector_2 s6903_7(wires_1725_6[3], addr_1725_6, addr_positional[27615:27612], addr_6903_7);

wire[31:0] addr_6904_7;

Selector_2 s6904_7(wires_1726_6[0], addr_1726_6, addr_positional[27619:27616], addr_6904_7);

wire[31:0] addr_6905_7;

Selector_2 s6905_7(wires_1726_6[1], addr_1726_6, addr_positional[27623:27620], addr_6905_7);

wire[31:0] addr_6906_7;

Selector_2 s6906_7(wires_1726_6[2], addr_1726_6, addr_positional[27627:27624], addr_6906_7);

wire[31:0] addr_6907_7;

Selector_2 s6907_7(wires_1726_6[3], addr_1726_6, addr_positional[27631:27628], addr_6907_7);

wire[31:0] addr_6908_7;

Selector_2 s6908_7(wires_1727_6[0], addr_1727_6, addr_positional[27635:27632], addr_6908_7);

wire[31:0] addr_6909_7;

Selector_2 s6909_7(wires_1727_6[1], addr_1727_6, addr_positional[27639:27636], addr_6909_7);

wire[31:0] addr_6910_7;

Selector_2 s6910_7(wires_1727_6[2], addr_1727_6, addr_positional[27643:27640], addr_6910_7);

wire[31:0] addr_6911_7;

Selector_2 s6911_7(wires_1727_6[3], addr_1727_6, addr_positional[27647:27644], addr_6911_7);

wire[31:0] addr_6912_7;

Selector_2 s6912_7(wires_1728_6[0], addr_1728_6, addr_positional[27651:27648], addr_6912_7);

wire[31:0] addr_6913_7;

Selector_2 s6913_7(wires_1728_6[1], addr_1728_6, addr_positional[27655:27652], addr_6913_7);

wire[31:0] addr_6914_7;

Selector_2 s6914_7(wires_1728_6[2], addr_1728_6, addr_positional[27659:27656], addr_6914_7);

wire[31:0] addr_6915_7;

Selector_2 s6915_7(wires_1728_6[3], addr_1728_6, addr_positional[27663:27660], addr_6915_7);

wire[31:0] addr_6916_7;

Selector_2 s6916_7(wires_1729_6[0], addr_1729_6, addr_positional[27667:27664], addr_6916_7);

wire[31:0] addr_6917_7;

Selector_2 s6917_7(wires_1729_6[1], addr_1729_6, addr_positional[27671:27668], addr_6917_7);

wire[31:0] addr_6918_7;

Selector_2 s6918_7(wires_1729_6[2], addr_1729_6, addr_positional[27675:27672], addr_6918_7);

wire[31:0] addr_6919_7;

Selector_2 s6919_7(wires_1729_6[3], addr_1729_6, addr_positional[27679:27676], addr_6919_7);

wire[31:0] addr_6920_7;

Selector_2 s6920_7(wires_1730_6[0], addr_1730_6, addr_positional[27683:27680], addr_6920_7);

wire[31:0] addr_6921_7;

Selector_2 s6921_7(wires_1730_6[1], addr_1730_6, addr_positional[27687:27684], addr_6921_7);

wire[31:0] addr_6922_7;

Selector_2 s6922_7(wires_1730_6[2], addr_1730_6, addr_positional[27691:27688], addr_6922_7);

wire[31:0] addr_6923_7;

Selector_2 s6923_7(wires_1730_6[3], addr_1730_6, addr_positional[27695:27692], addr_6923_7);

wire[31:0] addr_6924_7;

Selector_2 s6924_7(wires_1731_6[0], addr_1731_6, addr_positional[27699:27696], addr_6924_7);

wire[31:0] addr_6925_7;

Selector_2 s6925_7(wires_1731_6[1], addr_1731_6, addr_positional[27703:27700], addr_6925_7);

wire[31:0] addr_6926_7;

Selector_2 s6926_7(wires_1731_6[2], addr_1731_6, addr_positional[27707:27704], addr_6926_7);

wire[31:0] addr_6927_7;

Selector_2 s6927_7(wires_1731_6[3], addr_1731_6, addr_positional[27711:27708], addr_6927_7);

wire[31:0] addr_6928_7;

Selector_2 s6928_7(wires_1732_6[0], addr_1732_6, addr_positional[27715:27712], addr_6928_7);

wire[31:0] addr_6929_7;

Selector_2 s6929_7(wires_1732_6[1], addr_1732_6, addr_positional[27719:27716], addr_6929_7);

wire[31:0] addr_6930_7;

Selector_2 s6930_7(wires_1732_6[2], addr_1732_6, addr_positional[27723:27720], addr_6930_7);

wire[31:0] addr_6931_7;

Selector_2 s6931_7(wires_1732_6[3], addr_1732_6, addr_positional[27727:27724], addr_6931_7);

wire[31:0] addr_6932_7;

Selector_2 s6932_7(wires_1733_6[0], addr_1733_6, addr_positional[27731:27728], addr_6932_7);

wire[31:0] addr_6933_7;

Selector_2 s6933_7(wires_1733_6[1], addr_1733_6, addr_positional[27735:27732], addr_6933_7);

wire[31:0] addr_6934_7;

Selector_2 s6934_7(wires_1733_6[2], addr_1733_6, addr_positional[27739:27736], addr_6934_7);

wire[31:0] addr_6935_7;

Selector_2 s6935_7(wires_1733_6[3], addr_1733_6, addr_positional[27743:27740], addr_6935_7);

wire[31:0] addr_6936_7;

Selector_2 s6936_7(wires_1734_6[0], addr_1734_6, addr_positional[27747:27744], addr_6936_7);

wire[31:0] addr_6937_7;

Selector_2 s6937_7(wires_1734_6[1], addr_1734_6, addr_positional[27751:27748], addr_6937_7);

wire[31:0] addr_6938_7;

Selector_2 s6938_7(wires_1734_6[2], addr_1734_6, addr_positional[27755:27752], addr_6938_7);

wire[31:0] addr_6939_7;

Selector_2 s6939_7(wires_1734_6[3], addr_1734_6, addr_positional[27759:27756], addr_6939_7);

wire[31:0] addr_6940_7;

Selector_2 s6940_7(wires_1735_6[0], addr_1735_6, addr_positional[27763:27760], addr_6940_7);

wire[31:0] addr_6941_7;

Selector_2 s6941_7(wires_1735_6[1], addr_1735_6, addr_positional[27767:27764], addr_6941_7);

wire[31:0] addr_6942_7;

Selector_2 s6942_7(wires_1735_6[2], addr_1735_6, addr_positional[27771:27768], addr_6942_7);

wire[31:0] addr_6943_7;

Selector_2 s6943_7(wires_1735_6[3], addr_1735_6, addr_positional[27775:27772], addr_6943_7);

wire[31:0] addr_6944_7;

Selector_2 s6944_7(wires_1736_6[0], addr_1736_6, addr_positional[27779:27776], addr_6944_7);

wire[31:0] addr_6945_7;

Selector_2 s6945_7(wires_1736_6[1], addr_1736_6, addr_positional[27783:27780], addr_6945_7);

wire[31:0] addr_6946_7;

Selector_2 s6946_7(wires_1736_6[2], addr_1736_6, addr_positional[27787:27784], addr_6946_7);

wire[31:0] addr_6947_7;

Selector_2 s6947_7(wires_1736_6[3], addr_1736_6, addr_positional[27791:27788], addr_6947_7);

wire[31:0] addr_6948_7;

Selector_2 s6948_7(wires_1737_6[0], addr_1737_6, addr_positional[27795:27792], addr_6948_7);

wire[31:0] addr_6949_7;

Selector_2 s6949_7(wires_1737_6[1], addr_1737_6, addr_positional[27799:27796], addr_6949_7);

wire[31:0] addr_6950_7;

Selector_2 s6950_7(wires_1737_6[2], addr_1737_6, addr_positional[27803:27800], addr_6950_7);

wire[31:0] addr_6951_7;

Selector_2 s6951_7(wires_1737_6[3], addr_1737_6, addr_positional[27807:27804], addr_6951_7);

wire[31:0] addr_6952_7;

Selector_2 s6952_7(wires_1738_6[0], addr_1738_6, addr_positional[27811:27808], addr_6952_7);

wire[31:0] addr_6953_7;

Selector_2 s6953_7(wires_1738_6[1], addr_1738_6, addr_positional[27815:27812], addr_6953_7);

wire[31:0] addr_6954_7;

Selector_2 s6954_7(wires_1738_6[2], addr_1738_6, addr_positional[27819:27816], addr_6954_7);

wire[31:0] addr_6955_7;

Selector_2 s6955_7(wires_1738_6[3], addr_1738_6, addr_positional[27823:27820], addr_6955_7);

wire[31:0] addr_6956_7;

Selector_2 s6956_7(wires_1739_6[0], addr_1739_6, addr_positional[27827:27824], addr_6956_7);

wire[31:0] addr_6957_7;

Selector_2 s6957_7(wires_1739_6[1], addr_1739_6, addr_positional[27831:27828], addr_6957_7);

wire[31:0] addr_6958_7;

Selector_2 s6958_7(wires_1739_6[2], addr_1739_6, addr_positional[27835:27832], addr_6958_7);

wire[31:0] addr_6959_7;

Selector_2 s6959_7(wires_1739_6[3], addr_1739_6, addr_positional[27839:27836], addr_6959_7);

wire[31:0] addr_6960_7;

Selector_2 s6960_7(wires_1740_6[0], addr_1740_6, addr_positional[27843:27840], addr_6960_7);

wire[31:0] addr_6961_7;

Selector_2 s6961_7(wires_1740_6[1], addr_1740_6, addr_positional[27847:27844], addr_6961_7);

wire[31:0] addr_6962_7;

Selector_2 s6962_7(wires_1740_6[2], addr_1740_6, addr_positional[27851:27848], addr_6962_7);

wire[31:0] addr_6963_7;

Selector_2 s6963_7(wires_1740_6[3], addr_1740_6, addr_positional[27855:27852], addr_6963_7);

wire[31:0] addr_6964_7;

Selector_2 s6964_7(wires_1741_6[0], addr_1741_6, addr_positional[27859:27856], addr_6964_7);

wire[31:0] addr_6965_7;

Selector_2 s6965_7(wires_1741_6[1], addr_1741_6, addr_positional[27863:27860], addr_6965_7);

wire[31:0] addr_6966_7;

Selector_2 s6966_7(wires_1741_6[2], addr_1741_6, addr_positional[27867:27864], addr_6966_7);

wire[31:0] addr_6967_7;

Selector_2 s6967_7(wires_1741_6[3], addr_1741_6, addr_positional[27871:27868], addr_6967_7);

wire[31:0] addr_6968_7;

Selector_2 s6968_7(wires_1742_6[0], addr_1742_6, addr_positional[27875:27872], addr_6968_7);

wire[31:0] addr_6969_7;

Selector_2 s6969_7(wires_1742_6[1], addr_1742_6, addr_positional[27879:27876], addr_6969_7);

wire[31:0] addr_6970_7;

Selector_2 s6970_7(wires_1742_6[2], addr_1742_6, addr_positional[27883:27880], addr_6970_7);

wire[31:0] addr_6971_7;

Selector_2 s6971_7(wires_1742_6[3], addr_1742_6, addr_positional[27887:27884], addr_6971_7);

wire[31:0] addr_6972_7;

Selector_2 s6972_7(wires_1743_6[0], addr_1743_6, addr_positional[27891:27888], addr_6972_7);

wire[31:0] addr_6973_7;

Selector_2 s6973_7(wires_1743_6[1], addr_1743_6, addr_positional[27895:27892], addr_6973_7);

wire[31:0] addr_6974_7;

Selector_2 s6974_7(wires_1743_6[2], addr_1743_6, addr_positional[27899:27896], addr_6974_7);

wire[31:0] addr_6975_7;

Selector_2 s6975_7(wires_1743_6[3], addr_1743_6, addr_positional[27903:27900], addr_6975_7);

wire[31:0] addr_6976_7;

Selector_2 s6976_7(wires_1744_6[0], addr_1744_6, addr_positional[27907:27904], addr_6976_7);

wire[31:0] addr_6977_7;

Selector_2 s6977_7(wires_1744_6[1], addr_1744_6, addr_positional[27911:27908], addr_6977_7);

wire[31:0] addr_6978_7;

Selector_2 s6978_7(wires_1744_6[2], addr_1744_6, addr_positional[27915:27912], addr_6978_7);

wire[31:0] addr_6979_7;

Selector_2 s6979_7(wires_1744_6[3], addr_1744_6, addr_positional[27919:27916], addr_6979_7);

wire[31:0] addr_6980_7;

Selector_2 s6980_7(wires_1745_6[0], addr_1745_6, addr_positional[27923:27920], addr_6980_7);

wire[31:0] addr_6981_7;

Selector_2 s6981_7(wires_1745_6[1], addr_1745_6, addr_positional[27927:27924], addr_6981_7);

wire[31:0] addr_6982_7;

Selector_2 s6982_7(wires_1745_6[2], addr_1745_6, addr_positional[27931:27928], addr_6982_7);

wire[31:0] addr_6983_7;

Selector_2 s6983_7(wires_1745_6[3], addr_1745_6, addr_positional[27935:27932], addr_6983_7);

wire[31:0] addr_6984_7;

Selector_2 s6984_7(wires_1746_6[0], addr_1746_6, addr_positional[27939:27936], addr_6984_7);

wire[31:0] addr_6985_7;

Selector_2 s6985_7(wires_1746_6[1], addr_1746_6, addr_positional[27943:27940], addr_6985_7);

wire[31:0] addr_6986_7;

Selector_2 s6986_7(wires_1746_6[2], addr_1746_6, addr_positional[27947:27944], addr_6986_7);

wire[31:0] addr_6987_7;

Selector_2 s6987_7(wires_1746_6[3], addr_1746_6, addr_positional[27951:27948], addr_6987_7);

wire[31:0] addr_6988_7;

Selector_2 s6988_7(wires_1747_6[0], addr_1747_6, addr_positional[27955:27952], addr_6988_7);

wire[31:0] addr_6989_7;

Selector_2 s6989_7(wires_1747_6[1], addr_1747_6, addr_positional[27959:27956], addr_6989_7);

wire[31:0] addr_6990_7;

Selector_2 s6990_7(wires_1747_6[2], addr_1747_6, addr_positional[27963:27960], addr_6990_7);

wire[31:0] addr_6991_7;

Selector_2 s6991_7(wires_1747_6[3], addr_1747_6, addr_positional[27967:27964], addr_6991_7);

wire[31:0] addr_6992_7;

Selector_2 s6992_7(wires_1748_6[0], addr_1748_6, addr_positional[27971:27968], addr_6992_7);

wire[31:0] addr_6993_7;

Selector_2 s6993_7(wires_1748_6[1], addr_1748_6, addr_positional[27975:27972], addr_6993_7);

wire[31:0] addr_6994_7;

Selector_2 s6994_7(wires_1748_6[2], addr_1748_6, addr_positional[27979:27976], addr_6994_7);

wire[31:0] addr_6995_7;

Selector_2 s6995_7(wires_1748_6[3], addr_1748_6, addr_positional[27983:27980], addr_6995_7);

wire[31:0] addr_6996_7;

Selector_2 s6996_7(wires_1749_6[0], addr_1749_6, addr_positional[27987:27984], addr_6996_7);

wire[31:0] addr_6997_7;

Selector_2 s6997_7(wires_1749_6[1], addr_1749_6, addr_positional[27991:27988], addr_6997_7);

wire[31:0] addr_6998_7;

Selector_2 s6998_7(wires_1749_6[2], addr_1749_6, addr_positional[27995:27992], addr_6998_7);

wire[31:0] addr_6999_7;

Selector_2 s6999_7(wires_1749_6[3], addr_1749_6, addr_positional[27999:27996], addr_6999_7);

wire[31:0] addr_7000_7;

Selector_2 s7000_7(wires_1750_6[0], addr_1750_6, addr_positional[28003:28000], addr_7000_7);

wire[31:0] addr_7001_7;

Selector_2 s7001_7(wires_1750_6[1], addr_1750_6, addr_positional[28007:28004], addr_7001_7);

wire[31:0] addr_7002_7;

Selector_2 s7002_7(wires_1750_6[2], addr_1750_6, addr_positional[28011:28008], addr_7002_7);

wire[31:0] addr_7003_7;

Selector_2 s7003_7(wires_1750_6[3], addr_1750_6, addr_positional[28015:28012], addr_7003_7);

wire[31:0] addr_7004_7;

Selector_2 s7004_7(wires_1751_6[0], addr_1751_6, addr_positional[28019:28016], addr_7004_7);

wire[31:0] addr_7005_7;

Selector_2 s7005_7(wires_1751_6[1], addr_1751_6, addr_positional[28023:28020], addr_7005_7);

wire[31:0] addr_7006_7;

Selector_2 s7006_7(wires_1751_6[2], addr_1751_6, addr_positional[28027:28024], addr_7006_7);

wire[31:0] addr_7007_7;

Selector_2 s7007_7(wires_1751_6[3], addr_1751_6, addr_positional[28031:28028], addr_7007_7);

wire[31:0] addr_7008_7;

Selector_2 s7008_7(wires_1752_6[0], addr_1752_6, addr_positional[28035:28032], addr_7008_7);

wire[31:0] addr_7009_7;

Selector_2 s7009_7(wires_1752_6[1], addr_1752_6, addr_positional[28039:28036], addr_7009_7);

wire[31:0] addr_7010_7;

Selector_2 s7010_7(wires_1752_6[2], addr_1752_6, addr_positional[28043:28040], addr_7010_7);

wire[31:0] addr_7011_7;

Selector_2 s7011_7(wires_1752_6[3], addr_1752_6, addr_positional[28047:28044], addr_7011_7);

wire[31:0] addr_7012_7;

Selector_2 s7012_7(wires_1753_6[0], addr_1753_6, addr_positional[28051:28048], addr_7012_7);

wire[31:0] addr_7013_7;

Selector_2 s7013_7(wires_1753_6[1], addr_1753_6, addr_positional[28055:28052], addr_7013_7);

wire[31:0] addr_7014_7;

Selector_2 s7014_7(wires_1753_6[2], addr_1753_6, addr_positional[28059:28056], addr_7014_7);

wire[31:0] addr_7015_7;

Selector_2 s7015_7(wires_1753_6[3], addr_1753_6, addr_positional[28063:28060], addr_7015_7);

wire[31:0] addr_7016_7;

Selector_2 s7016_7(wires_1754_6[0], addr_1754_6, addr_positional[28067:28064], addr_7016_7);

wire[31:0] addr_7017_7;

Selector_2 s7017_7(wires_1754_6[1], addr_1754_6, addr_positional[28071:28068], addr_7017_7);

wire[31:0] addr_7018_7;

Selector_2 s7018_7(wires_1754_6[2], addr_1754_6, addr_positional[28075:28072], addr_7018_7);

wire[31:0] addr_7019_7;

Selector_2 s7019_7(wires_1754_6[3], addr_1754_6, addr_positional[28079:28076], addr_7019_7);

wire[31:0] addr_7020_7;

Selector_2 s7020_7(wires_1755_6[0], addr_1755_6, addr_positional[28083:28080], addr_7020_7);

wire[31:0] addr_7021_7;

Selector_2 s7021_7(wires_1755_6[1], addr_1755_6, addr_positional[28087:28084], addr_7021_7);

wire[31:0] addr_7022_7;

Selector_2 s7022_7(wires_1755_6[2], addr_1755_6, addr_positional[28091:28088], addr_7022_7);

wire[31:0] addr_7023_7;

Selector_2 s7023_7(wires_1755_6[3], addr_1755_6, addr_positional[28095:28092], addr_7023_7);

wire[31:0] addr_7024_7;

Selector_2 s7024_7(wires_1756_6[0], addr_1756_6, addr_positional[28099:28096], addr_7024_7);

wire[31:0] addr_7025_7;

Selector_2 s7025_7(wires_1756_6[1], addr_1756_6, addr_positional[28103:28100], addr_7025_7);

wire[31:0] addr_7026_7;

Selector_2 s7026_7(wires_1756_6[2], addr_1756_6, addr_positional[28107:28104], addr_7026_7);

wire[31:0] addr_7027_7;

Selector_2 s7027_7(wires_1756_6[3], addr_1756_6, addr_positional[28111:28108], addr_7027_7);

wire[31:0] addr_7028_7;

Selector_2 s7028_7(wires_1757_6[0], addr_1757_6, addr_positional[28115:28112], addr_7028_7);

wire[31:0] addr_7029_7;

Selector_2 s7029_7(wires_1757_6[1], addr_1757_6, addr_positional[28119:28116], addr_7029_7);

wire[31:0] addr_7030_7;

Selector_2 s7030_7(wires_1757_6[2], addr_1757_6, addr_positional[28123:28120], addr_7030_7);

wire[31:0] addr_7031_7;

Selector_2 s7031_7(wires_1757_6[3], addr_1757_6, addr_positional[28127:28124], addr_7031_7);

wire[31:0] addr_7032_7;

Selector_2 s7032_7(wires_1758_6[0], addr_1758_6, addr_positional[28131:28128], addr_7032_7);

wire[31:0] addr_7033_7;

Selector_2 s7033_7(wires_1758_6[1], addr_1758_6, addr_positional[28135:28132], addr_7033_7);

wire[31:0] addr_7034_7;

Selector_2 s7034_7(wires_1758_6[2], addr_1758_6, addr_positional[28139:28136], addr_7034_7);

wire[31:0] addr_7035_7;

Selector_2 s7035_7(wires_1758_6[3], addr_1758_6, addr_positional[28143:28140], addr_7035_7);

wire[31:0] addr_7036_7;

Selector_2 s7036_7(wires_1759_6[0], addr_1759_6, addr_positional[28147:28144], addr_7036_7);

wire[31:0] addr_7037_7;

Selector_2 s7037_7(wires_1759_6[1], addr_1759_6, addr_positional[28151:28148], addr_7037_7);

wire[31:0] addr_7038_7;

Selector_2 s7038_7(wires_1759_6[2], addr_1759_6, addr_positional[28155:28152], addr_7038_7);

wire[31:0] addr_7039_7;

Selector_2 s7039_7(wires_1759_6[3], addr_1759_6, addr_positional[28159:28156], addr_7039_7);

wire[31:0] addr_7040_7;

Selector_2 s7040_7(wires_1760_6[0], addr_1760_6, addr_positional[28163:28160], addr_7040_7);

wire[31:0] addr_7041_7;

Selector_2 s7041_7(wires_1760_6[1], addr_1760_6, addr_positional[28167:28164], addr_7041_7);

wire[31:0] addr_7042_7;

Selector_2 s7042_7(wires_1760_6[2], addr_1760_6, addr_positional[28171:28168], addr_7042_7);

wire[31:0] addr_7043_7;

Selector_2 s7043_7(wires_1760_6[3], addr_1760_6, addr_positional[28175:28172], addr_7043_7);

wire[31:0] addr_7044_7;

Selector_2 s7044_7(wires_1761_6[0], addr_1761_6, addr_positional[28179:28176], addr_7044_7);

wire[31:0] addr_7045_7;

Selector_2 s7045_7(wires_1761_6[1], addr_1761_6, addr_positional[28183:28180], addr_7045_7);

wire[31:0] addr_7046_7;

Selector_2 s7046_7(wires_1761_6[2], addr_1761_6, addr_positional[28187:28184], addr_7046_7);

wire[31:0] addr_7047_7;

Selector_2 s7047_7(wires_1761_6[3], addr_1761_6, addr_positional[28191:28188], addr_7047_7);

wire[31:0] addr_7048_7;

Selector_2 s7048_7(wires_1762_6[0], addr_1762_6, addr_positional[28195:28192], addr_7048_7);

wire[31:0] addr_7049_7;

Selector_2 s7049_7(wires_1762_6[1], addr_1762_6, addr_positional[28199:28196], addr_7049_7);

wire[31:0] addr_7050_7;

Selector_2 s7050_7(wires_1762_6[2], addr_1762_6, addr_positional[28203:28200], addr_7050_7);

wire[31:0] addr_7051_7;

Selector_2 s7051_7(wires_1762_6[3], addr_1762_6, addr_positional[28207:28204], addr_7051_7);

wire[31:0] addr_7052_7;

Selector_2 s7052_7(wires_1763_6[0], addr_1763_6, addr_positional[28211:28208], addr_7052_7);

wire[31:0] addr_7053_7;

Selector_2 s7053_7(wires_1763_6[1], addr_1763_6, addr_positional[28215:28212], addr_7053_7);

wire[31:0] addr_7054_7;

Selector_2 s7054_7(wires_1763_6[2], addr_1763_6, addr_positional[28219:28216], addr_7054_7);

wire[31:0] addr_7055_7;

Selector_2 s7055_7(wires_1763_6[3], addr_1763_6, addr_positional[28223:28220], addr_7055_7);

wire[31:0] addr_7056_7;

Selector_2 s7056_7(wires_1764_6[0], addr_1764_6, addr_positional[28227:28224], addr_7056_7);

wire[31:0] addr_7057_7;

Selector_2 s7057_7(wires_1764_6[1], addr_1764_6, addr_positional[28231:28228], addr_7057_7);

wire[31:0] addr_7058_7;

Selector_2 s7058_7(wires_1764_6[2], addr_1764_6, addr_positional[28235:28232], addr_7058_7);

wire[31:0] addr_7059_7;

Selector_2 s7059_7(wires_1764_6[3], addr_1764_6, addr_positional[28239:28236], addr_7059_7);

wire[31:0] addr_7060_7;

Selector_2 s7060_7(wires_1765_6[0], addr_1765_6, addr_positional[28243:28240], addr_7060_7);

wire[31:0] addr_7061_7;

Selector_2 s7061_7(wires_1765_6[1], addr_1765_6, addr_positional[28247:28244], addr_7061_7);

wire[31:0] addr_7062_7;

Selector_2 s7062_7(wires_1765_6[2], addr_1765_6, addr_positional[28251:28248], addr_7062_7);

wire[31:0] addr_7063_7;

Selector_2 s7063_7(wires_1765_6[3], addr_1765_6, addr_positional[28255:28252], addr_7063_7);

wire[31:0] addr_7064_7;

Selector_2 s7064_7(wires_1766_6[0], addr_1766_6, addr_positional[28259:28256], addr_7064_7);

wire[31:0] addr_7065_7;

Selector_2 s7065_7(wires_1766_6[1], addr_1766_6, addr_positional[28263:28260], addr_7065_7);

wire[31:0] addr_7066_7;

Selector_2 s7066_7(wires_1766_6[2], addr_1766_6, addr_positional[28267:28264], addr_7066_7);

wire[31:0] addr_7067_7;

Selector_2 s7067_7(wires_1766_6[3], addr_1766_6, addr_positional[28271:28268], addr_7067_7);

wire[31:0] addr_7068_7;

Selector_2 s7068_7(wires_1767_6[0], addr_1767_6, addr_positional[28275:28272], addr_7068_7);

wire[31:0] addr_7069_7;

Selector_2 s7069_7(wires_1767_6[1], addr_1767_6, addr_positional[28279:28276], addr_7069_7);

wire[31:0] addr_7070_7;

Selector_2 s7070_7(wires_1767_6[2], addr_1767_6, addr_positional[28283:28280], addr_7070_7);

wire[31:0] addr_7071_7;

Selector_2 s7071_7(wires_1767_6[3], addr_1767_6, addr_positional[28287:28284], addr_7071_7);

wire[31:0] addr_7072_7;

Selector_2 s7072_7(wires_1768_6[0], addr_1768_6, addr_positional[28291:28288], addr_7072_7);

wire[31:0] addr_7073_7;

Selector_2 s7073_7(wires_1768_6[1], addr_1768_6, addr_positional[28295:28292], addr_7073_7);

wire[31:0] addr_7074_7;

Selector_2 s7074_7(wires_1768_6[2], addr_1768_6, addr_positional[28299:28296], addr_7074_7);

wire[31:0] addr_7075_7;

Selector_2 s7075_7(wires_1768_6[3], addr_1768_6, addr_positional[28303:28300], addr_7075_7);

wire[31:0] addr_7076_7;

Selector_2 s7076_7(wires_1769_6[0], addr_1769_6, addr_positional[28307:28304], addr_7076_7);

wire[31:0] addr_7077_7;

Selector_2 s7077_7(wires_1769_6[1], addr_1769_6, addr_positional[28311:28308], addr_7077_7);

wire[31:0] addr_7078_7;

Selector_2 s7078_7(wires_1769_6[2], addr_1769_6, addr_positional[28315:28312], addr_7078_7);

wire[31:0] addr_7079_7;

Selector_2 s7079_7(wires_1769_6[3], addr_1769_6, addr_positional[28319:28316], addr_7079_7);

wire[31:0] addr_7080_7;

Selector_2 s7080_7(wires_1770_6[0], addr_1770_6, addr_positional[28323:28320], addr_7080_7);

wire[31:0] addr_7081_7;

Selector_2 s7081_7(wires_1770_6[1], addr_1770_6, addr_positional[28327:28324], addr_7081_7);

wire[31:0] addr_7082_7;

Selector_2 s7082_7(wires_1770_6[2], addr_1770_6, addr_positional[28331:28328], addr_7082_7);

wire[31:0] addr_7083_7;

Selector_2 s7083_7(wires_1770_6[3], addr_1770_6, addr_positional[28335:28332], addr_7083_7);

wire[31:0] addr_7084_7;

Selector_2 s7084_7(wires_1771_6[0], addr_1771_6, addr_positional[28339:28336], addr_7084_7);

wire[31:0] addr_7085_7;

Selector_2 s7085_7(wires_1771_6[1], addr_1771_6, addr_positional[28343:28340], addr_7085_7);

wire[31:0] addr_7086_7;

Selector_2 s7086_7(wires_1771_6[2], addr_1771_6, addr_positional[28347:28344], addr_7086_7);

wire[31:0] addr_7087_7;

Selector_2 s7087_7(wires_1771_6[3], addr_1771_6, addr_positional[28351:28348], addr_7087_7);

wire[31:0] addr_7088_7;

Selector_2 s7088_7(wires_1772_6[0], addr_1772_6, addr_positional[28355:28352], addr_7088_7);

wire[31:0] addr_7089_7;

Selector_2 s7089_7(wires_1772_6[1], addr_1772_6, addr_positional[28359:28356], addr_7089_7);

wire[31:0] addr_7090_7;

Selector_2 s7090_7(wires_1772_6[2], addr_1772_6, addr_positional[28363:28360], addr_7090_7);

wire[31:0] addr_7091_7;

Selector_2 s7091_7(wires_1772_6[3], addr_1772_6, addr_positional[28367:28364], addr_7091_7);

wire[31:0] addr_7092_7;

Selector_2 s7092_7(wires_1773_6[0], addr_1773_6, addr_positional[28371:28368], addr_7092_7);

wire[31:0] addr_7093_7;

Selector_2 s7093_7(wires_1773_6[1], addr_1773_6, addr_positional[28375:28372], addr_7093_7);

wire[31:0] addr_7094_7;

Selector_2 s7094_7(wires_1773_6[2], addr_1773_6, addr_positional[28379:28376], addr_7094_7);

wire[31:0] addr_7095_7;

Selector_2 s7095_7(wires_1773_6[3], addr_1773_6, addr_positional[28383:28380], addr_7095_7);

wire[31:0] addr_7096_7;

Selector_2 s7096_7(wires_1774_6[0], addr_1774_6, addr_positional[28387:28384], addr_7096_7);

wire[31:0] addr_7097_7;

Selector_2 s7097_7(wires_1774_6[1], addr_1774_6, addr_positional[28391:28388], addr_7097_7);

wire[31:0] addr_7098_7;

Selector_2 s7098_7(wires_1774_6[2], addr_1774_6, addr_positional[28395:28392], addr_7098_7);

wire[31:0] addr_7099_7;

Selector_2 s7099_7(wires_1774_6[3], addr_1774_6, addr_positional[28399:28396], addr_7099_7);

wire[31:0] addr_7100_7;

Selector_2 s7100_7(wires_1775_6[0], addr_1775_6, addr_positional[28403:28400], addr_7100_7);

wire[31:0] addr_7101_7;

Selector_2 s7101_7(wires_1775_6[1], addr_1775_6, addr_positional[28407:28404], addr_7101_7);

wire[31:0] addr_7102_7;

Selector_2 s7102_7(wires_1775_6[2], addr_1775_6, addr_positional[28411:28408], addr_7102_7);

wire[31:0] addr_7103_7;

Selector_2 s7103_7(wires_1775_6[3], addr_1775_6, addr_positional[28415:28412], addr_7103_7);

wire[31:0] addr_7104_7;

Selector_2 s7104_7(wires_1776_6[0], addr_1776_6, addr_positional[28419:28416], addr_7104_7);

wire[31:0] addr_7105_7;

Selector_2 s7105_7(wires_1776_6[1], addr_1776_6, addr_positional[28423:28420], addr_7105_7);

wire[31:0] addr_7106_7;

Selector_2 s7106_7(wires_1776_6[2], addr_1776_6, addr_positional[28427:28424], addr_7106_7);

wire[31:0] addr_7107_7;

Selector_2 s7107_7(wires_1776_6[3], addr_1776_6, addr_positional[28431:28428], addr_7107_7);

wire[31:0] addr_7108_7;

Selector_2 s7108_7(wires_1777_6[0], addr_1777_6, addr_positional[28435:28432], addr_7108_7);

wire[31:0] addr_7109_7;

Selector_2 s7109_7(wires_1777_6[1], addr_1777_6, addr_positional[28439:28436], addr_7109_7);

wire[31:0] addr_7110_7;

Selector_2 s7110_7(wires_1777_6[2], addr_1777_6, addr_positional[28443:28440], addr_7110_7);

wire[31:0] addr_7111_7;

Selector_2 s7111_7(wires_1777_6[3], addr_1777_6, addr_positional[28447:28444], addr_7111_7);

wire[31:0] addr_7112_7;

Selector_2 s7112_7(wires_1778_6[0], addr_1778_6, addr_positional[28451:28448], addr_7112_7);

wire[31:0] addr_7113_7;

Selector_2 s7113_7(wires_1778_6[1], addr_1778_6, addr_positional[28455:28452], addr_7113_7);

wire[31:0] addr_7114_7;

Selector_2 s7114_7(wires_1778_6[2], addr_1778_6, addr_positional[28459:28456], addr_7114_7);

wire[31:0] addr_7115_7;

Selector_2 s7115_7(wires_1778_6[3], addr_1778_6, addr_positional[28463:28460], addr_7115_7);

wire[31:0] addr_7116_7;

Selector_2 s7116_7(wires_1779_6[0], addr_1779_6, addr_positional[28467:28464], addr_7116_7);

wire[31:0] addr_7117_7;

Selector_2 s7117_7(wires_1779_6[1], addr_1779_6, addr_positional[28471:28468], addr_7117_7);

wire[31:0] addr_7118_7;

Selector_2 s7118_7(wires_1779_6[2], addr_1779_6, addr_positional[28475:28472], addr_7118_7);

wire[31:0] addr_7119_7;

Selector_2 s7119_7(wires_1779_6[3], addr_1779_6, addr_positional[28479:28476], addr_7119_7);

wire[31:0] addr_7120_7;

Selector_2 s7120_7(wires_1780_6[0], addr_1780_6, addr_positional[28483:28480], addr_7120_7);

wire[31:0] addr_7121_7;

Selector_2 s7121_7(wires_1780_6[1], addr_1780_6, addr_positional[28487:28484], addr_7121_7);

wire[31:0] addr_7122_7;

Selector_2 s7122_7(wires_1780_6[2], addr_1780_6, addr_positional[28491:28488], addr_7122_7);

wire[31:0] addr_7123_7;

Selector_2 s7123_7(wires_1780_6[3], addr_1780_6, addr_positional[28495:28492], addr_7123_7);

wire[31:0] addr_7124_7;

Selector_2 s7124_7(wires_1781_6[0], addr_1781_6, addr_positional[28499:28496], addr_7124_7);

wire[31:0] addr_7125_7;

Selector_2 s7125_7(wires_1781_6[1], addr_1781_6, addr_positional[28503:28500], addr_7125_7);

wire[31:0] addr_7126_7;

Selector_2 s7126_7(wires_1781_6[2], addr_1781_6, addr_positional[28507:28504], addr_7126_7);

wire[31:0] addr_7127_7;

Selector_2 s7127_7(wires_1781_6[3], addr_1781_6, addr_positional[28511:28508], addr_7127_7);

wire[31:0] addr_7128_7;

Selector_2 s7128_7(wires_1782_6[0], addr_1782_6, addr_positional[28515:28512], addr_7128_7);

wire[31:0] addr_7129_7;

Selector_2 s7129_7(wires_1782_6[1], addr_1782_6, addr_positional[28519:28516], addr_7129_7);

wire[31:0] addr_7130_7;

Selector_2 s7130_7(wires_1782_6[2], addr_1782_6, addr_positional[28523:28520], addr_7130_7);

wire[31:0] addr_7131_7;

Selector_2 s7131_7(wires_1782_6[3], addr_1782_6, addr_positional[28527:28524], addr_7131_7);

wire[31:0] addr_7132_7;

Selector_2 s7132_7(wires_1783_6[0], addr_1783_6, addr_positional[28531:28528], addr_7132_7);

wire[31:0] addr_7133_7;

Selector_2 s7133_7(wires_1783_6[1], addr_1783_6, addr_positional[28535:28532], addr_7133_7);

wire[31:0] addr_7134_7;

Selector_2 s7134_7(wires_1783_6[2], addr_1783_6, addr_positional[28539:28536], addr_7134_7);

wire[31:0] addr_7135_7;

Selector_2 s7135_7(wires_1783_6[3], addr_1783_6, addr_positional[28543:28540], addr_7135_7);

wire[31:0] addr_7136_7;

Selector_2 s7136_7(wires_1784_6[0], addr_1784_6, addr_positional[28547:28544], addr_7136_7);

wire[31:0] addr_7137_7;

Selector_2 s7137_7(wires_1784_6[1], addr_1784_6, addr_positional[28551:28548], addr_7137_7);

wire[31:0] addr_7138_7;

Selector_2 s7138_7(wires_1784_6[2], addr_1784_6, addr_positional[28555:28552], addr_7138_7);

wire[31:0] addr_7139_7;

Selector_2 s7139_7(wires_1784_6[3], addr_1784_6, addr_positional[28559:28556], addr_7139_7);

wire[31:0] addr_7140_7;

Selector_2 s7140_7(wires_1785_6[0], addr_1785_6, addr_positional[28563:28560], addr_7140_7);

wire[31:0] addr_7141_7;

Selector_2 s7141_7(wires_1785_6[1], addr_1785_6, addr_positional[28567:28564], addr_7141_7);

wire[31:0] addr_7142_7;

Selector_2 s7142_7(wires_1785_6[2], addr_1785_6, addr_positional[28571:28568], addr_7142_7);

wire[31:0] addr_7143_7;

Selector_2 s7143_7(wires_1785_6[3], addr_1785_6, addr_positional[28575:28572], addr_7143_7);

wire[31:0] addr_7144_7;

Selector_2 s7144_7(wires_1786_6[0], addr_1786_6, addr_positional[28579:28576], addr_7144_7);

wire[31:0] addr_7145_7;

Selector_2 s7145_7(wires_1786_6[1], addr_1786_6, addr_positional[28583:28580], addr_7145_7);

wire[31:0] addr_7146_7;

Selector_2 s7146_7(wires_1786_6[2], addr_1786_6, addr_positional[28587:28584], addr_7146_7);

wire[31:0] addr_7147_7;

Selector_2 s7147_7(wires_1786_6[3], addr_1786_6, addr_positional[28591:28588], addr_7147_7);

wire[31:0] addr_7148_7;

Selector_2 s7148_7(wires_1787_6[0], addr_1787_6, addr_positional[28595:28592], addr_7148_7);

wire[31:0] addr_7149_7;

Selector_2 s7149_7(wires_1787_6[1], addr_1787_6, addr_positional[28599:28596], addr_7149_7);

wire[31:0] addr_7150_7;

Selector_2 s7150_7(wires_1787_6[2], addr_1787_6, addr_positional[28603:28600], addr_7150_7);

wire[31:0] addr_7151_7;

Selector_2 s7151_7(wires_1787_6[3], addr_1787_6, addr_positional[28607:28604], addr_7151_7);

wire[31:0] addr_7152_7;

Selector_2 s7152_7(wires_1788_6[0], addr_1788_6, addr_positional[28611:28608], addr_7152_7);

wire[31:0] addr_7153_7;

Selector_2 s7153_7(wires_1788_6[1], addr_1788_6, addr_positional[28615:28612], addr_7153_7);

wire[31:0] addr_7154_7;

Selector_2 s7154_7(wires_1788_6[2], addr_1788_6, addr_positional[28619:28616], addr_7154_7);

wire[31:0] addr_7155_7;

Selector_2 s7155_7(wires_1788_6[3], addr_1788_6, addr_positional[28623:28620], addr_7155_7);

wire[31:0] addr_7156_7;

Selector_2 s7156_7(wires_1789_6[0], addr_1789_6, addr_positional[28627:28624], addr_7156_7);

wire[31:0] addr_7157_7;

Selector_2 s7157_7(wires_1789_6[1], addr_1789_6, addr_positional[28631:28628], addr_7157_7);

wire[31:0] addr_7158_7;

Selector_2 s7158_7(wires_1789_6[2], addr_1789_6, addr_positional[28635:28632], addr_7158_7);

wire[31:0] addr_7159_7;

Selector_2 s7159_7(wires_1789_6[3], addr_1789_6, addr_positional[28639:28636], addr_7159_7);

wire[31:0] addr_7160_7;

Selector_2 s7160_7(wires_1790_6[0], addr_1790_6, addr_positional[28643:28640], addr_7160_7);

wire[31:0] addr_7161_7;

Selector_2 s7161_7(wires_1790_6[1], addr_1790_6, addr_positional[28647:28644], addr_7161_7);

wire[31:0] addr_7162_7;

Selector_2 s7162_7(wires_1790_6[2], addr_1790_6, addr_positional[28651:28648], addr_7162_7);

wire[31:0] addr_7163_7;

Selector_2 s7163_7(wires_1790_6[3], addr_1790_6, addr_positional[28655:28652], addr_7163_7);

wire[31:0] addr_7164_7;

Selector_2 s7164_7(wires_1791_6[0], addr_1791_6, addr_positional[28659:28656], addr_7164_7);

wire[31:0] addr_7165_7;

Selector_2 s7165_7(wires_1791_6[1], addr_1791_6, addr_positional[28663:28660], addr_7165_7);

wire[31:0] addr_7166_7;

Selector_2 s7166_7(wires_1791_6[2], addr_1791_6, addr_positional[28667:28664], addr_7166_7);

wire[31:0] addr_7167_7;

Selector_2 s7167_7(wires_1791_6[3], addr_1791_6, addr_positional[28671:28668], addr_7167_7);

wire[31:0] addr_7168_7;

Selector_2 s7168_7(wires_1792_6[0], addr_1792_6, addr_positional[28675:28672], addr_7168_7);

wire[31:0] addr_7169_7;

Selector_2 s7169_7(wires_1792_6[1], addr_1792_6, addr_positional[28679:28676], addr_7169_7);

wire[31:0] addr_7170_7;

Selector_2 s7170_7(wires_1792_6[2], addr_1792_6, addr_positional[28683:28680], addr_7170_7);

wire[31:0] addr_7171_7;

Selector_2 s7171_7(wires_1792_6[3], addr_1792_6, addr_positional[28687:28684], addr_7171_7);

wire[31:0] addr_7172_7;

Selector_2 s7172_7(wires_1793_6[0], addr_1793_6, addr_positional[28691:28688], addr_7172_7);

wire[31:0] addr_7173_7;

Selector_2 s7173_7(wires_1793_6[1], addr_1793_6, addr_positional[28695:28692], addr_7173_7);

wire[31:0] addr_7174_7;

Selector_2 s7174_7(wires_1793_6[2], addr_1793_6, addr_positional[28699:28696], addr_7174_7);

wire[31:0] addr_7175_7;

Selector_2 s7175_7(wires_1793_6[3], addr_1793_6, addr_positional[28703:28700], addr_7175_7);

wire[31:0] addr_7176_7;

Selector_2 s7176_7(wires_1794_6[0], addr_1794_6, addr_positional[28707:28704], addr_7176_7);

wire[31:0] addr_7177_7;

Selector_2 s7177_7(wires_1794_6[1], addr_1794_6, addr_positional[28711:28708], addr_7177_7);

wire[31:0] addr_7178_7;

Selector_2 s7178_7(wires_1794_6[2], addr_1794_6, addr_positional[28715:28712], addr_7178_7);

wire[31:0] addr_7179_7;

Selector_2 s7179_7(wires_1794_6[3], addr_1794_6, addr_positional[28719:28716], addr_7179_7);

wire[31:0] addr_7180_7;

Selector_2 s7180_7(wires_1795_6[0], addr_1795_6, addr_positional[28723:28720], addr_7180_7);

wire[31:0] addr_7181_7;

Selector_2 s7181_7(wires_1795_6[1], addr_1795_6, addr_positional[28727:28724], addr_7181_7);

wire[31:0] addr_7182_7;

Selector_2 s7182_7(wires_1795_6[2], addr_1795_6, addr_positional[28731:28728], addr_7182_7);

wire[31:0] addr_7183_7;

Selector_2 s7183_7(wires_1795_6[3], addr_1795_6, addr_positional[28735:28732], addr_7183_7);

wire[31:0] addr_7184_7;

Selector_2 s7184_7(wires_1796_6[0], addr_1796_6, addr_positional[28739:28736], addr_7184_7);

wire[31:0] addr_7185_7;

Selector_2 s7185_7(wires_1796_6[1], addr_1796_6, addr_positional[28743:28740], addr_7185_7);

wire[31:0] addr_7186_7;

Selector_2 s7186_7(wires_1796_6[2], addr_1796_6, addr_positional[28747:28744], addr_7186_7);

wire[31:0] addr_7187_7;

Selector_2 s7187_7(wires_1796_6[3], addr_1796_6, addr_positional[28751:28748], addr_7187_7);

wire[31:0] addr_7188_7;

Selector_2 s7188_7(wires_1797_6[0], addr_1797_6, addr_positional[28755:28752], addr_7188_7);

wire[31:0] addr_7189_7;

Selector_2 s7189_7(wires_1797_6[1], addr_1797_6, addr_positional[28759:28756], addr_7189_7);

wire[31:0] addr_7190_7;

Selector_2 s7190_7(wires_1797_6[2], addr_1797_6, addr_positional[28763:28760], addr_7190_7);

wire[31:0] addr_7191_7;

Selector_2 s7191_7(wires_1797_6[3], addr_1797_6, addr_positional[28767:28764], addr_7191_7);

wire[31:0] addr_7192_7;

Selector_2 s7192_7(wires_1798_6[0], addr_1798_6, addr_positional[28771:28768], addr_7192_7);

wire[31:0] addr_7193_7;

Selector_2 s7193_7(wires_1798_6[1], addr_1798_6, addr_positional[28775:28772], addr_7193_7);

wire[31:0] addr_7194_7;

Selector_2 s7194_7(wires_1798_6[2], addr_1798_6, addr_positional[28779:28776], addr_7194_7);

wire[31:0] addr_7195_7;

Selector_2 s7195_7(wires_1798_6[3], addr_1798_6, addr_positional[28783:28780], addr_7195_7);

wire[31:0] addr_7196_7;

Selector_2 s7196_7(wires_1799_6[0], addr_1799_6, addr_positional[28787:28784], addr_7196_7);

wire[31:0] addr_7197_7;

Selector_2 s7197_7(wires_1799_6[1], addr_1799_6, addr_positional[28791:28788], addr_7197_7);

wire[31:0] addr_7198_7;

Selector_2 s7198_7(wires_1799_6[2], addr_1799_6, addr_positional[28795:28792], addr_7198_7);

wire[31:0] addr_7199_7;

Selector_2 s7199_7(wires_1799_6[3], addr_1799_6, addr_positional[28799:28796], addr_7199_7);

wire[31:0] addr_7200_7;

Selector_2 s7200_7(wires_1800_6[0], addr_1800_6, addr_positional[28803:28800], addr_7200_7);

wire[31:0] addr_7201_7;

Selector_2 s7201_7(wires_1800_6[1], addr_1800_6, addr_positional[28807:28804], addr_7201_7);

wire[31:0] addr_7202_7;

Selector_2 s7202_7(wires_1800_6[2], addr_1800_6, addr_positional[28811:28808], addr_7202_7);

wire[31:0] addr_7203_7;

Selector_2 s7203_7(wires_1800_6[3], addr_1800_6, addr_positional[28815:28812], addr_7203_7);

wire[31:0] addr_7204_7;

Selector_2 s7204_7(wires_1801_6[0], addr_1801_6, addr_positional[28819:28816], addr_7204_7);

wire[31:0] addr_7205_7;

Selector_2 s7205_7(wires_1801_6[1], addr_1801_6, addr_positional[28823:28820], addr_7205_7);

wire[31:0] addr_7206_7;

Selector_2 s7206_7(wires_1801_6[2], addr_1801_6, addr_positional[28827:28824], addr_7206_7);

wire[31:0] addr_7207_7;

Selector_2 s7207_7(wires_1801_6[3], addr_1801_6, addr_positional[28831:28828], addr_7207_7);

wire[31:0] addr_7208_7;

Selector_2 s7208_7(wires_1802_6[0], addr_1802_6, addr_positional[28835:28832], addr_7208_7);

wire[31:0] addr_7209_7;

Selector_2 s7209_7(wires_1802_6[1], addr_1802_6, addr_positional[28839:28836], addr_7209_7);

wire[31:0] addr_7210_7;

Selector_2 s7210_7(wires_1802_6[2], addr_1802_6, addr_positional[28843:28840], addr_7210_7);

wire[31:0] addr_7211_7;

Selector_2 s7211_7(wires_1802_6[3], addr_1802_6, addr_positional[28847:28844], addr_7211_7);

wire[31:0] addr_7212_7;

Selector_2 s7212_7(wires_1803_6[0], addr_1803_6, addr_positional[28851:28848], addr_7212_7);

wire[31:0] addr_7213_7;

Selector_2 s7213_7(wires_1803_6[1], addr_1803_6, addr_positional[28855:28852], addr_7213_7);

wire[31:0] addr_7214_7;

Selector_2 s7214_7(wires_1803_6[2], addr_1803_6, addr_positional[28859:28856], addr_7214_7);

wire[31:0] addr_7215_7;

Selector_2 s7215_7(wires_1803_6[3], addr_1803_6, addr_positional[28863:28860], addr_7215_7);

wire[31:0] addr_7216_7;

Selector_2 s7216_7(wires_1804_6[0], addr_1804_6, addr_positional[28867:28864], addr_7216_7);

wire[31:0] addr_7217_7;

Selector_2 s7217_7(wires_1804_6[1], addr_1804_6, addr_positional[28871:28868], addr_7217_7);

wire[31:0] addr_7218_7;

Selector_2 s7218_7(wires_1804_6[2], addr_1804_6, addr_positional[28875:28872], addr_7218_7);

wire[31:0] addr_7219_7;

Selector_2 s7219_7(wires_1804_6[3], addr_1804_6, addr_positional[28879:28876], addr_7219_7);

wire[31:0] addr_7220_7;

Selector_2 s7220_7(wires_1805_6[0], addr_1805_6, addr_positional[28883:28880], addr_7220_7);

wire[31:0] addr_7221_7;

Selector_2 s7221_7(wires_1805_6[1], addr_1805_6, addr_positional[28887:28884], addr_7221_7);

wire[31:0] addr_7222_7;

Selector_2 s7222_7(wires_1805_6[2], addr_1805_6, addr_positional[28891:28888], addr_7222_7);

wire[31:0] addr_7223_7;

Selector_2 s7223_7(wires_1805_6[3], addr_1805_6, addr_positional[28895:28892], addr_7223_7);

wire[31:0] addr_7224_7;

Selector_2 s7224_7(wires_1806_6[0], addr_1806_6, addr_positional[28899:28896], addr_7224_7);

wire[31:0] addr_7225_7;

Selector_2 s7225_7(wires_1806_6[1], addr_1806_6, addr_positional[28903:28900], addr_7225_7);

wire[31:0] addr_7226_7;

Selector_2 s7226_7(wires_1806_6[2], addr_1806_6, addr_positional[28907:28904], addr_7226_7);

wire[31:0] addr_7227_7;

Selector_2 s7227_7(wires_1806_6[3], addr_1806_6, addr_positional[28911:28908], addr_7227_7);

wire[31:0] addr_7228_7;

Selector_2 s7228_7(wires_1807_6[0], addr_1807_6, addr_positional[28915:28912], addr_7228_7);

wire[31:0] addr_7229_7;

Selector_2 s7229_7(wires_1807_6[1], addr_1807_6, addr_positional[28919:28916], addr_7229_7);

wire[31:0] addr_7230_7;

Selector_2 s7230_7(wires_1807_6[2], addr_1807_6, addr_positional[28923:28920], addr_7230_7);

wire[31:0] addr_7231_7;

Selector_2 s7231_7(wires_1807_6[3], addr_1807_6, addr_positional[28927:28924], addr_7231_7);

wire[31:0] addr_7232_7;

Selector_2 s7232_7(wires_1808_6[0], addr_1808_6, addr_positional[28931:28928], addr_7232_7);

wire[31:0] addr_7233_7;

Selector_2 s7233_7(wires_1808_6[1], addr_1808_6, addr_positional[28935:28932], addr_7233_7);

wire[31:0] addr_7234_7;

Selector_2 s7234_7(wires_1808_6[2], addr_1808_6, addr_positional[28939:28936], addr_7234_7);

wire[31:0] addr_7235_7;

Selector_2 s7235_7(wires_1808_6[3], addr_1808_6, addr_positional[28943:28940], addr_7235_7);

wire[31:0] addr_7236_7;

Selector_2 s7236_7(wires_1809_6[0], addr_1809_6, addr_positional[28947:28944], addr_7236_7);

wire[31:0] addr_7237_7;

Selector_2 s7237_7(wires_1809_6[1], addr_1809_6, addr_positional[28951:28948], addr_7237_7);

wire[31:0] addr_7238_7;

Selector_2 s7238_7(wires_1809_6[2], addr_1809_6, addr_positional[28955:28952], addr_7238_7);

wire[31:0] addr_7239_7;

Selector_2 s7239_7(wires_1809_6[3], addr_1809_6, addr_positional[28959:28956], addr_7239_7);

wire[31:0] addr_7240_7;

Selector_2 s7240_7(wires_1810_6[0], addr_1810_6, addr_positional[28963:28960], addr_7240_7);

wire[31:0] addr_7241_7;

Selector_2 s7241_7(wires_1810_6[1], addr_1810_6, addr_positional[28967:28964], addr_7241_7);

wire[31:0] addr_7242_7;

Selector_2 s7242_7(wires_1810_6[2], addr_1810_6, addr_positional[28971:28968], addr_7242_7);

wire[31:0] addr_7243_7;

Selector_2 s7243_7(wires_1810_6[3], addr_1810_6, addr_positional[28975:28972], addr_7243_7);

wire[31:0] addr_7244_7;

Selector_2 s7244_7(wires_1811_6[0], addr_1811_6, addr_positional[28979:28976], addr_7244_7);

wire[31:0] addr_7245_7;

Selector_2 s7245_7(wires_1811_6[1], addr_1811_6, addr_positional[28983:28980], addr_7245_7);

wire[31:0] addr_7246_7;

Selector_2 s7246_7(wires_1811_6[2], addr_1811_6, addr_positional[28987:28984], addr_7246_7);

wire[31:0] addr_7247_7;

Selector_2 s7247_7(wires_1811_6[3], addr_1811_6, addr_positional[28991:28988], addr_7247_7);

wire[31:0] addr_7248_7;

Selector_2 s7248_7(wires_1812_6[0], addr_1812_6, addr_positional[28995:28992], addr_7248_7);

wire[31:0] addr_7249_7;

Selector_2 s7249_7(wires_1812_6[1], addr_1812_6, addr_positional[28999:28996], addr_7249_7);

wire[31:0] addr_7250_7;

Selector_2 s7250_7(wires_1812_6[2], addr_1812_6, addr_positional[29003:29000], addr_7250_7);

wire[31:0] addr_7251_7;

Selector_2 s7251_7(wires_1812_6[3], addr_1812_6, addr_positional[29007:29004], addr_7251_7);

wire[31:0] addr_7252_7;

Selector_2 s7252_7(wires_1813_6[0], addr_1813_6, addr_positional[29011:29008], addr_7252_7);

wire[31:0] addr_7253_7;

Selector_2 s7253_7(wires_1813_6[1], addr_1813_6, addr_positional[29015:29012], addr_7253_7);

wire[31:0] addr_7254_7;

Selector_2 s7254_7(wires_1813_6[2], addr_1813_6, addr_positional[29019:29016], addr_7254_7);

wire[31:0] addr_7255_7;

Selector_2 s7255_7(wires_1813_6[3], addr_1813_6, addr_positional[29023:29020], addr_7255_7);

wire[31:0] addr_7256_7;

Selector_2 s7256_7(wires_1814_6[0], addr_1814_6, addr_positional[29027:29024], addr_7256_7);

wire[31:0] addr_7257_7;

Selector_2 s7257_7(wires_1814_6[1], addr_1814_6, addr_positional[29031:29028], addr_7257_7);

wire[31:0] addr_7258_7;

Selector_2 s7258_7(wires_1814_6[2], addr_1814_6, addr_positional[29035:29032], addr_7258_7);

wire[31:0] addr_7259_7;

Selector_2 s7259_7(wires_1814_6[3], addr_1814_6, addr_positional[29039:29036], addr_7259_7);

wire[31:0] addr_7260_7;

Selector_2 s7260_7(wires_1815_6[0], addr_1815_6, addr_positional[29043:29040], addr_7260_7);

wire[31:0] addr_7261_7;

Selector_2 s7261_7(wires_1815_6[1], addr_1815_6, addr_positional[29047:29044], addr_7261_7);

wire[31:0] addr_7262_7;

Selector_2 s7262_7(wires_1815_6[2], addr_1815_6, addr_positional[29051:29048], addr_7262_7);

wire[31:0] addr_7263_7;

Selector_2 s7263_7(wires_1815_6[3], addr_1815_6, addr_positional[29055:29052], addr_7263_7);

wire[31:0] addr_7264_7;

Selector_2 s7264_7(wires_1816_6[0], addr_1816_6, addr_positional[29059:29056], addr_7264_7);

wire[31:0] addr_7265_7;

Selector_2 s7265_7(wires_1816_6[1], addr_1816_6, addr_positional[29063:29060], addr_7265_7);

wire[31:0] addr_7266_7;

Selector_2 s7266_7(wires_1816_6[2], addr_1816_6, addr_positional[29067:29064], addr_7266_7);

wire[31:0] addr_7267_7;

Selector_2 s7267_7(wires_1816_6[3], addr_1816_6, addr_positional[29071:29068], addr_7267_7);

wire[31:0] addr_7268_7;

Selector_2 s7268_7(wires_1817_6[0], addr_1817_6, addr_positional[29075:29072], addr_7268_7);

wire[31:0] addr_7269_7;

Selector_2 s7269_7(wires_1817_6[1], addr_1817_6, addr_positional[29079:29076], addr_7269_7);

wire[31:0] addr_7270_7;

Selector_2 s7270_7(wires_1817_6[2], addr_1817_6, addr_positional[29083:29080], addr_7270_7);

wire[31:0] addr_7271_7;

Selector_2 s7271_7(wires_1817_6[3], addr_1817_6, addr_positional[29087:29084], addr_7271_7);

wire[31:0] addr_7272_7;

Selector_2 s7272_7(wires_1818_6[0], addr_1818_6, addr_positional[29091:29088], addr_7272_7);

wire[31:0] addr_7273_7;

Selector_2 s7273_7(wires_1818_6[1], addr_1818_6, addr_positional[29095:29092], addr_7273_7);

wire[31:0] addr_7274_7;

Selector_2 s7274_7(wires_1818_6[2], addr_1818_6, addr_positional[29099:29096], addr_7274_7);

wire[31:0] addr_7275_7;

Selector_2 s7275_7(wires_1818_6[3], addr_1818_6, addr_positional[29103:29100], addr_7275_7);

wire[31:0] addr_7276_7;

Selector_2 s7276_7(wires_1819_6[0], addr_1819_6, addr_positional[29107:29104], addr_7276_7);

wire[31:0] addr_7277_7;

Selector_2 s7277_7(wires_1819_6[1], addr_1819_6, addr_positional[29111:29108], addr_7277_7);

wire[31:0] addr_7278_7;

Selector_2 s7278_7(wires_1819_6[2], addr_1819_6, addr_positional[29115:29112], addr_7278_7);

wire[31:0] addr_7279_7;

Selector_2 s7279_7(wires_1819_6[3], addr_1819_6, addr_positional[29119:29116], addr_7279_7);

wire[31:0] addr_7280_7;

Selector_2 s7280_7(wires_1820_6[0], addr_1820_6, addr_positional[29123:29120], addr_7280_7);

wire[31:0] addr_7281_7;

Selector_2 s7281_7(wires_1820_6[1], addr_1820_6, addr_positional[29127:29124], addr_7281_7);

wire[31:0] addr_7282_7;

Selector_2 s7282_7(wires_1820_6[2], addr_1820_6, addr_positional[29131:29128], addr_7282_7);

wire[31:0] addr_7283_7;

Selector_2 s7283_7(wires_1820_6[3], addr_1820_6, addr_positional[29135:29132], addr_7283_7);

wire[31:0] addr_7284_7;

Selector_2 s7284_7(wires_1821_6[0], addr_1821_6, addr_positional[29139:29136], addr_7284_7);

wire[31:0] addr_7285_7;

Selector_2 s7285_7(wires_1821_6[1], addr_1821_6, addr_positional[29143:29140], addr_7285_7);

wire[31:0] addr_7286_7;

Selector_2 s7286_7(wires_1821_6[2], addr_1821_6, addr_positional[29147:29144], addr_7286_7);

wire[31:0] addr_7287_7;

Selector_2 s7287_7(wires_1821_6[3], addr_1821_6, addr_positional[29151:29148], addr_7287_7);

wire[31:0] addr_7288_7;

Selector_2 s7288_7(wires_1822_6[0], addr_1822_6, addr_positional[29155:29152], addr_7288_7);

wire[31:0] addr_7289_7;

Selector_2 s7289_7(wires_1822_6[1], addr_1822_6, addr_positional[29159:29156], addr_7289_7);

wire[31:0] addr_7290_7;

Selector_2 s7290_7(wires_1822_6[2], addr_1822_6, addr_positional[29163:29160], addr_7290_7);

wire[31:0] addr_7291_7;

Selector_2 s7291_7(wires_1822_6[3], addr_1822_6, addr_positional[29167:29164], addr_7291_7);

wire[31:0] addr_7292_7;

Selector_2 s7292_7(wires_1823_6[0], addr_1823_6, addr_positional[29171:29168], addr_7292_7);

wire[31:0] addr_7293_7;

Selector_2 s7293_7(wires_1823_6[1], addr_1823_6, addr_positional[29175:29172], addr_7293_7);

wire[31:0] addr_7294_7;

Selector_2 s7294_7(wires_1823_6[2], addr_1823_6, addr_positional[29179:29176], addr_7294_7);

wire[31:0] addr_7295_7;

Selector_2 s7295_7(wires_1823_6[3], addr_1823_6, addr_positional[29183:29180], addr_7295_7);

wire[31:0] addr_7296_7;

Selector_2 s7296_7(wires_1824_6[0], addr_1824_6, addr_positional[29187:29184], addr_7296_7);

wire[31:0] addr_7297_7;

Selector_2 s7297_7(wires_1824_6[1], addr_1824_6, addr_positional[29191:29188], addr_7297_7);

wire[31:0] addr_7298_7;

Selector_2 s7298_7(wires_1824_6[2], addr_1824_6, addr_positional[29195:29192], addr_7298_7);

wire[31:0] addr_7299_7;

Selector_2 s7299_7(wires_1824_6[3], addr_1824_6, addr_positional[29199:29196], addr_7299_7);

wire[31:0] addr_7300_7;

Selector_2 s7300_7(wires_1825_6[0], addr_1825_6, addr_positional[29203:29200], addr_7300_7);

wire[31:0] addr_7301_7;

Selector_2 s7301_7(wires_1825_6[1], addr_1825_6, addr_positional[29207:29204], addr_7301_7);

wire[31:0] addr_7302_7;

Selector_2 s7302_7(wires_1825_6[2], addr_1825_6, addr_positional[29211:29208], addr_7302_7);

wire[31:0] addr_7303_7;

Selector_2 s7303_7(wires_1825_6[3], addr_1825_6, addr_positional[29215:29212], addr_7303_7);

wire[31:0] addr_7304_7;

Selector_2 s7304_7(wires_1826_6[0], addr_1826_6, addr_positional[29219:29216], addr_7304_7);

wire[31:0] addr_7305_7;

Selector_2 s7305_7(wires_1826_6[1], addr_1826_6, addr_positional[29223:29220], addr_7305_7);

wire[31:0] addr_7306_7;

Selector_2 s7306_7(wires_1826_6[2], addr_1826_6, addr_positional[29227:29224], addr_7306_7);

wire[31:0] addr_7307_7;

Selector_2 s7307_7(wires_1826_6[3], addr_1826_6, addr_positional[29231:29228], addr_7307_7);

wire[31:0] addr_7308_7;

Selector_2 s7308_7(wires_1827_6[0], addr_1827_6, addr_positional[29235:29232], addr_7308_7);

wire[31:0] addr_7309_7;

Selector_2 s7309_7(wires_1827_6[1], addr_1827_6, addr_positional[29239:29236], addr_7309_7);

wire[31:0] addr_7310_7;

Selector_2 s7310_7(wires_1827_6[2], addr_1827_6, addr_positional[29243:29240], addr_7310_7);

wire[31:0] addr_7311_7;

Selector_2 s7311_7(wires_1827_6[3], addr_1827_6, addr_positional[29247:29244], addr_7311_7);

wire[31:0] addr_7312_7;

Selector_2 s7312_7(wires_1828_6[0], addr_1828_6, addr_positional[29251:29248], addr_7312_7);

wire[31:0] addr_7313_7;

Selector_2 s7313_7(wires_1828_6[1], addr_1828_6, addr_positional[29255:29252], addr_7313_7);

wire[31:0] addr_7314_7;

Selector_2 s7314_7(wires_1828_6[2], addr_1828_6, addr_positional[29259:29256], addr_7314_7);

wire[31:0] addr_7315_7;

Selector_2 s7315_7(wires_1828_6[3], addr_1828_6, addr_positional[29263:29260], addr_7315_7);

wire[31:0] addr_7316_7;

Selector_2 s7316_7(wires_1829_6[0], addr_1829_6, addr_positional[29267:29264], addr_7316_7);

wire[31:0] addr_7317_7;

Selector_2 s7317_7(wires_1829_6[1], addr_1829_6, addr_positional[29271:29268], addr_7317_7);

wire[31:0] addr_7318_7;

Selector_2 s7318_7(wires_1829_6[2], addr_1829_6, addr_positional[29275:29272], addr_7318_7);

wire[31:0] addr_7319_7;

Selector_2 s7319_7(wires_1829_6[3], addr_1829_6, addr_positional[29279:29276], addr_7319_7);

wire[31:0] addr_7320_7;

Selector_2 s7320_7(wires_1830_6[0], addr_1830_6, addr_positional[29283:29280], addr_7320_7);

wire[31:0] addr_7321_7;

Selector_2 s7321_7(wires_1830_6[1], addr_1830_6, addr_positional[29287:29284], addr_7321_7);

wire[31:0] addr_7322_7;

Selector_2 s7322_7(wires_1830_6[2], addr_1830_6, addr_positional[29291:29288], addr_7322_7);

wire[31:0] addr_7323_7;

Selector_2 s7323_7(wires_1830_6[3], addr_1830_6, addr_positional[29295:29292], addr_7323_7);

wire[31:0] addr_7324_7;

Selector_2 s7324_7(wires_1831_6[0], addr_1831_6, addr_positional[29299:29296], addr_7324_7);

wire[31:0] addr_7325_7;

Selector_2 s7325_7(wires_1831_6[1], addr_1831_6, addr_positional[29303:29300], addr_7325_7);

wire[31:0] addr_7326_7;

Selector_2 s7326_7(wires_1831_6[2], addr_1831_6, addr_positional[29307:29304], addr_7326_7);

wire[31:0] addr_7327_7;

Selector_2 s7327_7(wires_1831_6[3], addr_1831_6, addr_positional[29311:29308], addr_7327_7);

wire[31:0] addr_7328_7;

Selector_2 s7328_7(wires_1832_6[0], addr_1832_6, addr_positional[29315:29312], addr_7328_7);

wire[31:0] addr_7329_7;

Selector_2 s7329_7(wires_1832_6[1], addr_1832_6, addr_positional[29319:29316], addr_7329_7);

wire[31:0] addr_7330_7;

Selector_2 s7330_7(wires_1832_6[2], addr_1832_6, addr_positional[29323:29320], addr_7330_7);

wire[31:0] addr_7331_7;

Selector_2 s7331_7(wires_1832_6[3], addr_1832_6, addr_positional[29327:29324], addr_7331_7);

wire[31:0] addr_7332_7;

Selector_2 s7332_7(wires_1833_6[0], addr_1833_6, addr_positional[29331:29328], addr_7332_7);

wire[31:0] addr_7333_7;

Selector_2 s7333_7(wires_1833_6[1], addr_1833_6, addr_positional[29335:29332], addr_7333_7);

wire[31:0] addr_7334_7;

Selector_2 s7334_7(wires_1833_6[2], addr_1833_6, addr_positional[29339:29336], addr_7334_7);

wire[31:0] addr_7335_7;

Selector_2 s7335_7(wires_1833_6[3], addr_1833_6, addr_positional[29343:29340], addr_7335_7);

wire[31:0] addr_7336_7;

Selector_2 s7336_7(wires_1834_6[0], addr_1834_6, addr_positional[29347:29344], addr_7336_7);

wire[31:0] addr_7337_7;

Selector_2 s7337_7(wires_1834_6[1], addr_1834_6, addr_positional[29351:29348], addr_7337_7);

wire[31:0] addr_7338_7;

Selector_2 s7338_7(wires_1834_6[2], addr_1834_6, addr_positional[29355:29352], addr_7338_7);

wire[31:0] addr_7339_7;

Selector_2 s7339_7(wires_1834_6[3], addr_1834_6, addr_positional[29359:29356], addr_7339_7);

wire[31:0] addr_7340_7;

Selector_2 s7340_7(wires_1835_6[0], addr_1835_6, addr_positional[29363:29360], addr_7340_7);

wire[31:0] addr_7341_7;

Selector_2 s7341_7(wires_1835_6[1], addr_1835_6, addr_positional[29367:29364], addr_7341_7);

wire[31:0] addr_7342_7;

Selector_2 s7342_7(wires_1835_6[2], addr_1835_6, addr_positional[29371:29368], addr_7342_7);

wire[31:0] addr_7343_7;

Selector_2 s7343_7(wires_1835_6[3], addr_1835_6, addr_positional[29375:29372], addr_7343_7);

wire[31:0] addr_7344_7;

Selector_2 s7344_7(wires_1836_6[0], addr_1836_6, addr_positional[29379:29376], addr_7344_7);

wire[31:0] addr_7345_7;

Selector_2 s7345_7(wires_1836_6[1], addr_1836_6, addr_positional[29383:29380], addr_7345_7);

wire[31:0] addr_7346_7;

Selector_2 s7346_7(wires_1836_6[2], addr_1836_6, addr_positional[29387:29384], addr_7346_7);

wire[31:0] addr_7347_7;

Selector_2 s7347_7(wires_1836_6[3], addr_1836_6, addr_positional[29391:29388], addr_7347_7);

wire[31:0] addr_7348_7;

Selector_2 s7348_7(wires_1837_6[0], addr_1837_6, addr_positional[29395:29392], addr_7348_7);

wire[31:0] addr_7349_7;

Selector_2 s7349_7(wires_1837_6[1], addr_1837_6, addr_positional[29399:29396], addr_7349_7);

wire[31:0] addr_7350_7;

Selector_2 s7350_7(wires_1837_6[2], addr_1837_6, addr_positional[29403:29400], addr_7350_7);

wire[31:0] addr_7351_7;

Selector_2 s7351_7(wires_1837_6[3], addr_1837_6, addr_positional[29407:29404], addr_7351_7);

wire[31:0] addr_7352_7;

Selector_2 s7352_7(wires_1838_6[0], addr_1838_6, addr_positional[29411:29408], addr_7352_7);

wire[31:0] addr_7353_7;

Selector_2 s7353_7(wires_1838_6[1], addr_1838_6, addr_positional[29415:29412], addr_7353_7);

wire[31:0] addr_7354_7;

Selector_2 s7354_7(wires_1838_6[2], addr_1838_6, addr_positional[29419:29416], addr_7354_7);

wire[31:0] addr_7355_7;

Selector_2 s7355_7(wires_1838_6[3], addr_1838_6, addr_positional[29423:29420], addr_7355_7);

wire[31:0] addr_7356_7;

Selector_2 s7356_7(wires_1839_6[0], addr_1839_6, addr_positional[29427:29424], addr_7356_7);

wire[31:0] addr_7357_7;

Selector_2 s7357_7(wires_1839_6[1], addr_1839_6, addr_positional[29431:29428], addr_7357_7);

wire[31:0] addr_7358_7;

Selector_2 s7358_7(wires_1839_6[2], addr_1839_6, addr_positional[29435:29432], addr_7358_7);

wire[31:0] addr_7359_7;

Selector_2 s7359_7(wires_1839_6[3], addr_1839_6, addr_positional[29439:29436], addr_7359_7);

wire[31:0] addr_7360_7;

Selector_2 s7360_7(wires_1840_6[0], addr_1840_6, addr_positional[29443:29440], addr_7360_7);

wire[31:0] addr_7361_7;

Selector_2 s7361_7(wires_1840_6[1], addr_1840_6, addr_positional[29447:29444], addr_7361_7);

wire[31:0] addr_7362_7;

Selector_2 s7362_7(wires_1840_6[2], addr_1840_6, addr_positional[29451:29448], addr_7362_7);

wire[31:0] addr_7363_7;

Selector_2 s7363_7(wires_1840_6[3], addr_1840_6, addr_positional[29455:29452], addr_7363_7);

wire[31:0] addr_7364_7;

Selector_2 s7364_7(wires_1841_6[0], addr_1841_6, addr_positional[29459:29456], addr_7364_7);

wire[31:0] addr_7365_7;

Selector_2 s7365_7(wires_1841_6[1], addr_1841_6, addr_positional[29463:29460], addr_7365_7);

wire[31:0] addr_7366_7;

Selector_2 s7366_7(wires_1841_6[2], addr_1841_6, addr_positional[29467:29464], addr_7366_7);

wire[31:0] addr_7367_7;

Selector_2 s7367_7(wires_1841_6[3], addr_1841_6, addr_positional[29471:29468], addr_7367_7);

wire[31:0] addr_7368_7;

Selector_2 s7368_7(wires_1842_6[0], addr_1842_6, addr_positional[29475:29472], addr_7368_7);

wire[31:0] addr_7369_7;

Selector_2 s7369_7(wires_1842_6[1], addr_1842_6, addr_positional[29479:29476], addr_7369_7);

wire[31:0] addr_7370_7;

Selector_2 s7370_7(wires_1842_6[2], addr_1842_6, addr_positional[29483:29480], addr_7370_7);

wire[31:0] addr_7371_7;

Selector_2 s7371_7(wires_1842_6[3], addr_1842_6, addr_positional[29487:29484], addr_7371_7);

wire[31:0] addr_7372_7;

Selector_2 s7372_7(wires_1843_6[0], addr_1843_6, addr_positional[29491:29488], addr_7372_7);

wire[31:0] addr_7373_7;

Selector_2 s7373_7(wires_1843_6[1], addr_1843_6, addr_positional[29495:29492], addr_7373_7);

wire[31:0] addr_7374_7;

Selector_2 s7374_7(wires_1843_6[2], addr_1843_6, addr_positional[29499:29496], addr_7374_7);

wire[31:0] addr_7375_7;

Selector_2 s7375_7(wires_1843_6[3], addr_1843_6, addr_positional[29503:29500], addr_7375_7);

wire[31:0] addr_7376_7;

Selector_2 s7376_7(wires_1844_6[0], addr_1844_6, addr_positional[29507:29504], addr_7376_7);

wire[31:0] addr_7377_7;

Selector_2 s7377_7(wires_1844_6[1], addr_1844_6, addr_positional[29511:29508], addr_7377_7);

wire[31:0] addr_7378_7;

Selector_2 s7378_7(wires_1844_6[2], addr_1844_6, addr_positional[29515:29512], addr_7378_7);

wire[31:0] addr_7379_7;

Selector_2 s7379_7(wires_1844_6[3], addr_1844_6, addr_positional[29519:29516], addr_7379_7);

wire[31:0] addr_7380_7;

Selector_2 s7380_7(wires_1845_6[0], addr_1845_6, addr_positional[29523:29520], addr_7380_7);

wire[31:0] addr_7381_7;

Selector_2 s7381_7(wires_1845_6[1], addr_1845_6, addr_positional[29527:29524], addr_7381_7);

wire[31:0] addr_7382_7;

Selector_2 s7382_7(wires_1845_6[2], addr_1845_6, addr_positional[29531:29528], addr_7382_7);

wire[31:0] addr_7383_7;

Selector_2 s7383_7(wires_1845_6[3], addr_1845_6, addr_positional[29535:29532], addr_7383_7);

wire[31:0] addr_7384_7;

Selector_2 s7384_7(wires_1846_6[0], addr_1846_6, addr_positional[29539:29536], addr_7384_7);

wire[31:0] addr_7385_7;

Selector_2 s7385_7(wires_1846_6[1], addr_1846_6, addr_positional[29543:29540], addr_7385_7);

wire[31:0] addr_7386_7;

Selector_2 s7386_7(wires_1846_6[2], addr_1846_6, addr_positional[29547:29544], addr_7386_7);

wire[31:0] addr_7387_7;

Selector_2 s7387_7(wires_1846_6[3], addr_1846_6, addr_positional[29551:29548], addr_7387_7);

wire[31:0] addr_7388_7;

Selector_2 s7388_7(wires_1847_6[0], addr_1847_6, addr_positional[29555:29552], addr_7388_7);

wire[31:0] addr_7389_7;

Selector_2 s7389_7(wires_1847_6[1], addr_1847_6, addr_positional[29559:29556], addr_7389_7);

wire[31:0] addr_7390_7;

Selector_2 s7390_7(wires_1847_6[2], addr_1847_6, addr_positional[29563:29560], addr_7390_7);

wire[31:0] addr_7391_7;

Selector_2 s7391_7(wires_1847_6[3], addr_1847_6, addr_positional[29567:29564], addr_7391_7);

wire[31:0] addr_7392_7;

Selector_2 s7392_7(wires_1848_6[0], addr_1848_6, addr_positional[29571:29568], addr_7392_7);

wire[31:0] addr_7393_7;

Selector_2 s7393_7(wires_1848_6[1], addr_1848_6, addr_positional[29575:29572], addr_7393_7);

wire[31:0] addr_7394_7;

Selector_2 s7394_7(wires_1848_6[2], addr_1848_6, addr_positional[29579:29576], addr_7394_7);

wire[31:0] addr_7395_7;

Selector_2 s7395_7(wires_1848_6[3], addr_1848_6, addr_positional[29583:29580], addr_7395_7);

wire[31:0] addr_7396_7;

Selector_2 s7396_7(wires_1849_6[0], addr_1849_6, addr_positional[29587:29584], addr_7396_7);

wire[31:0] addr_7397_7;

Selector_2 s7397_7(wires_1849_6[1], addr_1849_6, addr_positional[29591:29588], addr_7397_7);

wire[31:0] addr_7398_7;

Selector_2 s7398_7(wires_1849_6[2], addr_1849_6, addr_positional[29595:29592], addr_7398_7);

wire[31:0] addr_7399_7;

Selector_2 s7399_7(wires_1849_6[3], addr_1849_6, addr_positional[29599:29596], addr_7399_7);

wire[31:0] addr_7400_7;

Selector_2 s7400_7(wires_1850_6[0], addr_1850_6, addr_positional[29603:29600], addr_7400_7);

wire[31:0] addr_7401_7;

Selector_2 s7401_7(wires_1850_6[1], addr_1850_6, addr_positional[29607:29604], addr_7401_7);

wire[31:0] addr_7402_7;

Selector_2 s7402_7(wires_1850_6[2], addr_1850_6, addr_positional[29611:29608], addr_7402_7);

wire[31:0] addr_7403_7;

Selector_2 s7403_7(wires_1850_6[3], addr_1850_6, addr_positional[29615:29612], addr_7403_7);

wire[31:0] addr_7404_7;

Selector_2 s7404_7(wires_1851_6[0], addr_1851_6, addr_positional[29619:29616], addr_7404_7);

wire[31:0] addr_7405_7;

Selector_2 s7405_7(wires_1851_6[1], addr_1851_6, addr_positional[29623:29620], addr_7405_7);

wire[31:0] addr_7406_7;

Selector_2 s7406_7(wires_1851_6[2], addr_1851_6, addr_positional[29627:29624], addr_7406_7);

wire[31:0] addr_7407_7;

Selector_2 s7407_7(wires_1851_6[3], addr_1851_6, addr_positional[29631:29628], addr_7407_7);

wire[31:0] addr_7408_7;

Selector_2 s7408_7(wires_1852_6[0], addr_1852_6, addr_positional[29635:29632], addr_7408_7);

wire[31:0] addr_7409_7;

Selector_2 s7409_7(wires_1852_6[1], addr_1852_6, addr_positional[29639:29636], addr_7409_7);

wire[31:0] addr_7410_7;

Selector_2 s7410_7(wires_1852_6[2], addr_1852_6, addr_positional[29643:29640], addr_7410_7);

wire[31:0] addr_7411_7;

Selector_2 s7411_7(wires_1852_6[3], addr_1852_6, addr_positional[29647:29644], addr_7411_7);

wire[31:0] addr_7412_7;

Selector_2 s7412_7(wires_1853_6[0], addr_1853_6, addr_positional[29651:29648], addr_7412_7);

wire[31:0] addr_7413_7;

Selector_2 s7413_7(wires_1853_6[1], addr_1853_6, addr_positional[29655:29652], addr_7413_7);

wire[31:0] addr_7414_7;

Selector_2 s7414_7(wires_1853_6[2], addr_1853_6, addr_positional[29659:29656], addr_7414_7);

wire[31:0] addr_7415_7;

Selector_2 s7415_7(wires_1853_6[3], addr_1853_6, addr_positional[29663:29660], addr_7415_7);

wire[31:0] addr_7416_7;

Selector_2 s7416_7(wires_1854_6[0], addr_1854_6, addr_positional[29667:29664], addr_7416_7);

wire[31:0] addr_7417_7;

Selector_2 s7417_7(wires_1854_6[1], addr_1854_6, addr_positional[29671:29668], addr_7417_7);

wire[31:0] addr_7418_7;

Selector_2 s7418_7(wires_1854_6[2], addr_1854_6, addr_positional[29675:29672], addr_7418_7);

wire[31:0] addr_7419_7;

Selector_2 s7419_7(wires_1854_6[3], addr_1854_6, addr_positional[29679:29676], addr_7419_7);

wire[31:0] addr_7420_7;

Selector_2 s7420_7(wires_1855_6[0], addr_1855_6, addr_positional[29683:29680], addr_7420_7);

wire[31:0] addr_7421_7;

Selector_2 s7421_7(wires_1855_6[1], addr_1855_6, addr_positional[29687:29684], addr_7421_7);

wire[31:0] addr_7422_7;

Selector_2 s7422_7(wires_1855_6[2], addr_1855_6, addr_positional[29691:29688], addr_7422_7);

wire[31:0] addr_7423_7;

Selector_2 s7423_7(wires_1855_6[3], addr_1855_6, addr_positional[29695:29692], addr_7423_7);

wire[31:0] addr_7424_7;

Selector_2 s7424_7(wires_1856_6[0], addr_1856_6, addr_positional[29699:29696], addr_7424_7);

wire[31:0] addr_7425_7;

Selector_2 s7425_7(wires_1856_6[1], addr_1856_6, addr_positional[29703:29700], addr_7425_7);

wire[31:0] addr_7426_7;

Selector_2 s7426_7(wires_1856_6[2], addr_1856_6, addr_positional[29707:29704], addr_7426_7);

wire[31:0] addr_7427_7;

Selector_2 s7427_7(wires_1856_6[3], addr_1856_6, addr_positional[29711:29708], addr_7427_7);

wire[31:0] addr_7428_7;

Selector_2 s7428_7(wires_1857_6[0], addr_1857_6, addr_positional[29715:29712], addr_7428_7);

wire[31:0] addr_7429_7;

Selector_2 s7429_7(wires_1857_6[1], addr_1857_6, addr_positional[29719:29716], addr_7429_7);

wire[31:0] addr_7430_7;

Selector_2 s7430_7(wires_1857_6[2], addr_1857_6, addr_positional[29723:29720], addr_7430_7);

wire[31:0] addr_7431_7;

Selector_2 s7431_7(wires_1857_6[3], addr_1857_6, addr_positional[29727:29724], addr_7431_7);

wire[31:0] addr_7432_7;

Selector_2 s7432_7(wires_1858_6[0], addr_1858_6, addr_positional[29731:29728], addr_7432_7);

wire[31:0] addr_7433_7;

Selector_2 s7433_7(wires_1858_6[1], addr_1858_6, addr_positional[29735:29732], addr_7433_7);

wire[31:0] addr_7434_7;

Selector_2 s7434_7(wires_1858_6[2], addr_1858_6, addr_positional[29739:29736], addr_7434_7);

wire[31:0] addr_7435_7;

Selector_2 s7435_7(wires_1858_6[3], addr_1858_6, addr_positional[29743:29740], addr_7435_7);

wire[31:0] addr_7436_7;

Selector_2 s7436_7(wires_1859_6[0], addr_1859_6, addr_positional[29747:29744], addr_7436_7);

wire[31:0] addr_7437_7;

Selector_2 s7437_7(wires_1859_6[1], addr_1859_6, addr_positional[29751:29748], addr_7437_7);

wire[31:0] addr_7438_7;

Selector_2 s7438_7(wires_1859_6[2], addr_1859_6, addr_positional[29755:29752], addr_7438_7);

wire[31:0] addr_7439_7;

Selector_2 s7439_7(wires_1859_6[3], addr_1859_6, addr_positional[29759:29756], addr_7439_7);

wire[31:0] addr_7440_7;

Selector_2 s7440_7(wires_1860_6[0], addr_1860_6, addr_positional[29763:29760], addr_7440_7);

wire[31:0] addr_7441_7;

Selector_2 s7441_7(wires_1860_6[1], addr_1860_6, addr_positional[29767:29764], addr_7441_7);

wire[31:0] addr_7442_7;

Selector_2 s7442_7(wires_1860_6[2], addr_1860_6, addr_positional[29771:29768], addr_7442_7);

wire[31:0] addr_7443_7;

Selector_2 s7443_7(wires_1860_6[3], addr_1860_6, addr_positional[29775:29772], addr_7443_7);

wire[31:0] addr_7444_7;

Selector_2 s7444_7(wires_1861_6[0], addr_1861_6, addr_positional[29779:29776], addr_7444_7);

wire[31:0] addr_7445_7;

Selector_2 s7445_7(wires_1861_6[1], addr_1861_6, addr_positional[29783:29780], addr_7445_7);

wire[31:0] addr_7446_7;

Selector_2 s7446_7(wires_1861_6[2], addr_1861_6, addr_positional[29787:29784], addr_7446_7);

wire[31:0] addr_7447_7;

Selector_2 s7447_7(wires_1861_6[3], addr_1861_6, addr_positional[29791:29788], addr_7447_7);

wire[31:0] addr_7448_7;

Selector_2 s7448_7(wires_1862_6[0], addr_1862_6, addr_positional[29795:29792], addr_7448_7);

wire[31:0] addr_7449_7;

Selector_2 s7449_7(wires_1862_6[1], addr_1862_6, addr_positional[29799:29796], addr_7449_7);

wire[31:0] addr_7450_7;

Selector_2 s7450_7(wires_1862_6[2], addr_1862_6, addr_positional[29803:29800], addr_7450_7);

wire[31:0] addr_7451_7;

Selector_2 s7451_7(wires_1862_6[3], addr_1862_6, addr_positional[29807:29804], addr_7451_7);

wire[31:0] addr_7452_7;

Selector_2 s7452_7(wires_1863_6[0], addr_1863_6, addr_positional[29811:29808], addr_7452_7);

wire[31:0] addr_7453_7;

Selector_2 s7453_7(wires_1863_6[1], addr_1863_6, addr_positional[29815:29812], addr_7453_7);

wire[31:0] addr_7454_7;

Selector_2 s7454_7(wires_1863_6[2], addr_1863_6, addr_positional[29819:29816], addr_7454_7);

wire[31:0] addr_7455_7;

Selector_2 s7455_7(wires_1863_6[3], addr_1863_6, addr_positional[29823:29820], addr_7455_7);

wire[31:0] addr_7456_7;

Selector_2 s7456_7(wires_1864_6[0], addr_1864_6, addr_positional[29827:29824], addr_7456_7);

wire[31:0] addr_7457_7;

Selector_2 s7457_7(wires_1864_6[1], addr_1864_6, addr_positional[29831:29828], addr_7457_7);

wire[31:0] addr_7458_7;

Selector_2 s7458_7(wires_1864_6[2], addr_1864_6, addr_positional[29835:29832], addr_7458_7);

wire[31:0] addr_7459_7;

Selector_2 s7459_7(wires_1864_6[3], addr_1864_6, addr_positional[29839:29836], addr_7459_7);

wire[31:0] addr_7460_7;

Selector_2 s7460_7(wires_1865_6[0], addr_1865_6, addr_positional[29843:29840], addr_7460_7);

wire[31:0] addr_7461_7;

Selector_2 s7461_7(wires_1865_6[1], addr_1865_6, addr_positional[29847:29844], addr_7461_7);

wire[31:0] addr_7462_7;

Selector_2 s7462_7(wires_1865_6[2], addr_1865_6, addr_positional[29851:29848], addr_7462_7);

wire[31:0] addr_7463_7;

Selector_2 s7463_7(wires_1865_6[3], addr_1865_6, addr_positional[29855:29852], addr_7463_7);

wire[31:0] addr_7464_7;

Selector_2 s7464_7(wires_1866_6[0], addr_1866_6, addr_positional[29859:29856], addr_7464_7);

wire[31:0] addr_7465_7;

Selector_2 s7465_7(wires_1866_6[1], addr_1866_6, addr_positional[29863:29860], addr_7465_7);

wire[31:0] addr_7466_7;

Selector_2 s7466_7(wires_1866_6[2], addr_1866_6, addr_positional[29867:29864], addr_7466_7);

wire[31:0] addr_7467_7;

Selector_2 s7467_7(wires_1866_6[3], addr_1866_6, addr_positional[29871:29868], addr_7467_7);

wire[31:0] addr_7468_7;

Selector_2 s7468_7(wires_1867_6[0], addr_1867_6, addr_positional[29875:29872], addr_7468_7);

wire[31:0] addr_7469_7;

Selector_2 s7469_7(wires_1867_6[1], addr_1867_6, addr_positional[29879:29876], addr_7469_7);

wire[31:0] addr_7470_7;

Selector_2 s7470_7(wires_1867_6[2], addr_1867_6, addr_positional[29883:29880], addr_7470_7);

wire[31:0] addr_7471_7;

Selector_2 s7471_7(wires_1867_6[3], addr_1867_6, addr_positional[29887:29884], addr_7471_7);

wire[31:0] addr_7472_7;

Selector_2 s7472_7(wires_1868_6[0], addr_1868_6, addr_positional[29891:29888], addr_7472_7);

wire[31:0] addr_7473_7;

Selector_2 s7473_7(wires_1868_6[1], addr_1868_6, addr_positional[29895:29892], addr_7473_7);

wire[31:0] addr_7474_7;

Selector_2 s7474_7(wires_1868_6[2], addr_1868_6, addr_positional[29899:29896], addr_7474_7);

wire[31:0] addr_7475_7;

Selector_2 s7475_7(wires_1868_6[3], addr_1868_6, addr_positional[29903:29900], addr_7475_7);

wire[31:0] addr_7476_7;

Selector_2 s7476_7(wires_1869_6[0], addr_1869_6, addr_positional[29907:29904], addr_7476_7);

wire[31:0] addr_7477_7;

Selector_2 s7477_7(wires_1869_6[1], addr_1869_6, addr_positional[29911:29908], addr_7477_7);

wire[31:0] addr_7478_7;

Selector_2 s7478_7(wires_1869_6[2], addr_1869_6, addr_positional[29915:29912], addr_7478_7);

wire[31:0] addr_7479_7;

Selector_2 s7479_7(wires_1869_6[3], addr_1869_6, addr_positional[29919:29916], addr_7479_7);

wire[31:0] addr_7480_7;

Selector_2 s7480_7(wires_1870_6[0], addr_1870_6, addr_positional[29923:29920], addr_7480_7);

wire[31:0] addr_7481_7;

Selector_2 s7481_7(wires_1870_6[1], addr_1870_6, addr_positional[29927:29924], addr_7481_7);

wire[31:0] addr_7482_7;

Selector_2 s7482_7(wires_1870_6[2], addr_1870_6, addr_positional[29931:29928], addr_7482_7);

wire[31:0] addr_7483_7;

Selector_2 s7483_7(wires_1870_6[3], addr_1870_6, addr_positional[29935:29932], addr_7483_7);

wire[31:0] addr_7484_7;

Selector_2 s7484_7(wires_1871_6[0], addr_1871_6, addr_positional[29939:29936], addr_7484_7);

wire[31:0] addr_7485_7;

Selector_2 s7485_7(wires_1871_6[1], addr_1871_6, addr_positional[29943:29940], addr_7485_7);

wire[31:0] addr_7486_7;

Selector_2 s7486_7(wires_1871_6[2], addr_1871_6, addr_positional[29947:29944], addr_7486_7);

wire[31:0] addr_7487_7;

Selector_2 s7487_7(wires_1871_6[3], addr_1871_6, addr_positional[29951:29948], addr_7487_7);

wire[31:0] addr_7488_7;

Selector_2 s7488_7(wires_1872_6[0], addr_1872_6, addr_positional[29955:29952], addr_7488_7);

wire[31:0] addr_7489_7;

Selector_2 s7489_7(wires_1872_6[1], addr_1872_6, addr_positional[29959:29956], addr_7489_7);

wire[31:0] addr_7490_7;

Selector_2 s7490_7(wires_1872_6[2], addr_1872_6, addr_positional[29963:29960], addr_7490_7);

wire[31:0] addr_7491_7;

Selector_2 s7491_7(wires_1872_6[3], addr_1872_6, addr_positional[29967:29964], addr_7491_7);

wire[31:0] addr_7492_7;

Selector_2 s7492_7(wires_1873_6[0], addr_1873_6, addr_positional[29971:29968], addr_7492_7);

wire[31:0] addr_7493_7;

Selector_2 s7493_7(wires_1873_6[1], addr_1873_6, addr_positional[29975:29972], addr_7493_7);

wire[31:0] addr_7494_7;

Selector_2 s7494_7(wires_1873_6[2], addr_1873_6, addr_positional[29979:29976], addr_7494_7);

wire[31:0] addr_7495_7;

Selector_2 s7495_7(wires_1873_6[3], addr_1873_6, addr_positional[29983:29980], addr_7495_7);

wire[31:0] addr_7496_7;

Selector_2 s7496_7(wires_1874_6[0], addr_1874_6, addr_positional[29987:29984], addr_7496_7);

wire[31:0] addr_7497_7;

Selector_2 s7497_7(wires_1874_6[1], addr_1874_6, addr_positional[29991:29988], addr_7497_7);

wire[31:0] addr_7498_7;

Selector_2 s7498_7(wires_1874_6[2], addr_1874_6, addr_positional[29995:29992], addr_7498_7);

wire[31:0] addr_7499_7;

Selector_2 s7499_7(wires_1874_6[3], addr_1874_6, addr_positional[29999:29996], addr_7499_7);

wire[31:0] addr_7500_7;

Selector_2 s7500_7(wires_1875_6[0], addr_1875_6, addr_positional[30003:30000], addr_7500_7);

wire[31:0] addr_7501_7;

Selector_2 s7501_7(wires_1875_6[1], addr_1875_6, addr_positional[30007:30004], addr_7501_7);

wire[31:0] addr_7502_7;

Selector_2 s7502_7(wires_1875_6[2], addr_1875_6, addr_positional[30011:30008], addr_7502_7);

wire[31:0] addr_7503_7;

Selector_2 s7503_7(wires_1875_6[3], addr_1875_6, addr_positional[30015:30012], addr_7503_7);

wire[31:0] addr_7504_7;

Selector_2 s7504_7(wires_1876_6[0], addr_1876_6, addr_positional[30019:30016], addr_7504_7);

wire[31:0] addr_7505_7;

Selector_2 s7505_7(wires_1876_6[1], addr_1876_6, addr_positional[30023:30020], addr_7505_7);

wire[31:0] addr_7506_7;

Selector_2 s7506_7(wires_1876_6[2], addr_1876_6, addr_positional[30027:30024], addr_7506_7);

wire[31:0] addr_7507_7;

Selector_2 s7507_7(wires_1876_6[3], addr_1876_6, addr_positional[30031:30028], addr_7507_7);

wire[31:0] addr_7508_7;

Selector_2 s7508_7(wires_1877_6[0], addr_1877_6, addr_positional[30035:30032], addr_7508_7);

wire[31:0] addr_7509_7;

Selector_2 s7509_7(wires_1877_6[1], addr_1877_6, addr_positional[30039:30036], addr_7509_7);

wire[31:0] addr_7510_7;

Selector_2 s7510_7(wires_1877_6[2], addr_1877_6, addr_positional[30043:30040], addr_7510_7);

wire[31:0] addr_7511_7;

Selector_2 s7511_7(wires_1877_6[3], addr_1877_6, addr_positional[30047:30044], addr_7511_7);

wire[31:0] addr_7512_7;

Selector_2 s7512_7(wires_1878_6[0], addr_1878_6, addr_positional[30051:30048], addr_7512_7);

wire[31:0] addr_7513_7;

Selector_2 s7513_7(wires_1878_6[1], addr_1878_6, addr_positional[30055:30052], addr_7513_7);

wire[31:0] addr_7514_7;

Selector_2 s7514_7(wires_1878_6[2], addr_1878_6, addr_positional[30059:30056], addr_7514_7);

wire[31:0] addr_7515_7;

Selector_2 s7515_7(wires_1878_6[3], addr_1878_6, addr_positional[30063:30060], addr_7515_7);

wire[31:0] addr_7516_7;

Selector_2 s7516_7(wires_1879_6[0], addr_1879_6, addr_positional[30067:30064], addr_7516_7);

wire[31:0] addr_7517_7;

Selector_2 s7517_7(wires_1879_6[1], addr_1879_6, addr_positional[30071:30068], addr_7517_7);

wire[31:0] addr_7518_7;

Selector_2 s7518_7(wires_1879_6[2], addr_1879_6, addr_positional[30075:30072], addr_7518_7);

wire[31:0] addr_7519_7;

Selector_2 s7519_7(wires_1879_6[3], addr_1879_6, addr_positional[30079:30076], addr_7519_7);

wire[31:0] addr_7520_7;

Selector_2 s7520_7(wires_1880_6[0], addr_1880_6, addr_positional[30083:30080], addr_7520_7);

wire[31:0] addr_7521_7;

Selector_2 s7521_7(wires_1880_6[1], addr_1880_6, addr_positional[30087:30084], addr_7521_7);

wire[31:0] addr_7522_7;

Selector_2 s7522_7(wires_1880_6[2], addr_1880_6, addr_positional[30091:30088], addr_7522_7);

wire[31:0] addr_7523_7;

Selector_2 s7523_7(wires_1880_6[3], addr_1880_6, addr_positional[30095:30092], addr_7523_7);

wire[31:0] addr_7524_7;

Selector_2 s7524_7(wires_1881_6[0], addr_1881_6, addr_positional[30099:30096], addr_7524_7);

wire[31:0] addr_7525_7;

Selector_2 s7525_7(wires_1881_6[1], addr_1881_6, addr_positional[30103:30100], addr_7525_7);

wire[31:0] addr_7526_7;

Selector_2 s7526_7(wires_1881_6[2], addr_1881_6, addr_positional[30107:30104], addr_7526_7);

wire[31:0] addr_7527_7;

Selector_2 s7527_7(wires_1881_6[3], addr_1881_6, addr_positional[30111:30108], addr_7527_7);

wire[31:0] addr_7528_7;

Selector_2 s7528_7(wires_1882_6[0], addr_1882_6, addr_positional[30115:30112], addr_7528_7);

wire[31:0] addr_7529_7;

Selector_2 s7529_7(wires_1882_6[1], addr_1882_6, addr_positional[30119:30116], addr_7529_7);

wire[31:0] addr_7530_7;

Selector_2 s7530_7(wires_1882_6[2], addr_1882_6, addr_positional[30123:30120], addr_7530_7);

wire[31:0] addr_7531_7;

Selector_2 s7531_7(wires_1882_6[3], addr_1882_6, addr_positional[30127:30124], addr_7531_7);

wire[31:0] addr_7532_7;

Selector_2 s7532_7(wires_1883_6[0], addr_1883_6, addr_positional[30131:30128], addr_7532_7);

wire[31:0] addr_7533_7;

Selector_2 s7533_7(wires_1883_6[1], addr_1883_6, addr_positional[30135:30132], addr_7533_7);

wire[31:0] addr_7534_7;

Selector_2 s7534_7(wires_1883_6[2], addr_1883_6, addr_positional[30139:30136], addr_7534_7);

wire[31:0] addr_7535_7;

Selector_2 s7535_7(wires_1883_6[3], addr_1883_6, addr_positional[30143:30140], addr_7535_7);

wire[31:0] addr_7536_7;

Selector_2 s7536_7(wires_1884_6[0], addr_1884_6, addr_positional[30147:30144], addr_7536_7);

wire[31:0] addr_7537_7;

Selector_2 s7537_7(wires_1884_6[1], addr_1884_6, addr_positional[30151:30148], addr_7537_7);

wire[31:0] addr_7538_7;

Selector_2 s7538_7(wires_1884_6[2], addr_1884_6, addr_positional[30155:30152], addr_7538_7);

wire[31:0] addr_7539_7;

Selector_2 s7539_7(wires_1884_6[3], addr_1884_6, addr_positional[30159:30156], addr_7539_7);

wire[31:0] addr_7540_7;

Selector_2 s7540_7(wires_1885_6[0], addr_1885_6, addr_positional[30163:30160], addr_7540_7);

wire[31:0] addr_7541_7;

Selector_2 s7541_7(wires_1885_6[1], addr_1885_6, addr_positional[30167:30164], addr_7541_7);

wire[31:0] addr_7542_7;

Selector_2 s7542_7(wires_1885_6[2], addr_1885_6, addr_positional[30171:30168], addr_7542_7);

wire[31:0] addr_7543_7;

Selector_2 s7543_7(wires_1885_6[3], addr_1885_6, addr_positional[30175:30172], addr_7543_7);

wire[31:0] addr_7544_7;

Selector_2 s7544_7(wires_1886_6[0], addr_1886_6, addr_positional[30179:30176], addr_7544_7);

wire[31:0] addr_7545_7;

Selector_2 s7545_7(wires_1886_6[1], addr_1886_6, addr_positional[30183:30180], addr_7545_7);

wire[31:0] addr_7546_7;

Selector_2 s7546_7(wires_1886_6[2], addr_1886_6, addr_positional[30187:30184], addr_7546_7);

wire[31:0] addr_7547_7;

Selector_2 s7547_7(wires_1886_6[3], addr_1886_6, addr_positional[30191:30188], addr_7547_7);

wire[31:0] addr_7548_7;

Selector_2 s7548_7(wires_1887_6[0], addr_1887_6, addr_positional[30195:30192], addr_7548_7);

wire[31:0] addr_7549_7;

Selector_2 s7549_7(wires_1887_6[1], addr_1887_6, addr_positional[30199:30196], addr_7549_7);

wire[31:0] addr_7550_7;

Selector_2 s7550_7(wires_1887_6[2], addr_1887_6, addr_positional[30203:30200], addr_7550_7);

wire[31:0] addr_7551_7;

Selector_2 s7551_7(wires_1887_6[3], addr_1887_6, addr_positional[30207:30204], addr_7551_7);

wire[31:0] addr_7552_7;

Selector_2 s7552_7(wires_1888_6[0], addr_1888_6, addr_positional[30211:30208], addr_7552_7);

wire[31:0] addr_7553_7;

Selector_2 s7553_7(wires_1888_6[1], addr_1888_6, addr_positional[30215:30212], addr_7553_7);

wire[31:0] addr_7554_7;

Selector_2 s7554_7(wires_1888_6[2], addr_1888_6, addr_positional[30219:30216], addr_7554_7);

wire[31:0] addr_7555_7;

Selector_2 s7555_7(wires_1888_6[3], addr_1888_6, addr_positional[30223:30220], addr_7555_7);

wire[31:0] addr_7556_7;

Selector_2 s7556_7(wires_1889_6[0], addr_1889_6, addr_positional[30227:30224], addr_7556_7);

wire[31:0] addr_7557_7;

Selector_2 s7557_7(wires_1889_6[1], addr_1889_6, addr_positional[30231:30228], addr_7557_7);

wire[31:0] addr_7558_7;

Selector_2 s7558_7(wires_1889_6[2], addr_1889_6, addr_positional[30235:30232], addr_7558_7);

wire[31:0] addr_7559_7;

Selector_2 s7559_7(wires_1889_6[3], addr_1889_6, addr_positional[30239:30236], addr_7559_7);

wire[31:0] addr_7560_7;

Selector_2 s7560_7(wires_1890_6[0], addr_1890_6, addr_positional[30243:30240], addr_7560_7);

wire[31:0] addr_7561_7;

Selector_2 s7561_7(wires_1890_6[1], addr_1890_6, addr_positional[30247:30244], addr_7561_7);

wire[31:0] addr_7562_7;

Selector_2 s7562_7(wires_1890_6[2], addr_1890_6, addr_positional[30251:30248], addr_7562_7);

wire[31:0] addr_7563_7;

Selector_2 s7563_7(wires_1890_6[3], addr_1890_6, addr_positional[30255:30252], addr_7563_7);

wire[31:0] addr_7564_7;

Selector_2 s7564_7(wires_1891_6[0], addr_1891_6, addr_positional[30259:30256], addr_7564_7);

wire[31:0] addr_7565_7;

Selector_2 s7565_7(wires_1891_6[1], addr_1891_6, addr_positional[30263:30260], addr_7565_7);

wire[31:0] addr_7566_7;

Selector_2 s7566_7(wires_1891_6[2], addr_1891_6, addr_positional[30267:30264], addr_7566_7);

wire[31:0] addr_7567_7;

Selector_2 s7567_7(wires_1891_6[3], addr_1891_6, addr_positional[30271:30268], addr_7567_7);

wire[31:0] addr_7568_7;

Selector_2 s7568_7(wires_1892_6[0], addr_1892_6, addr_positional[30275:30272], addr_7568_7);

wire[31:0] addr_7569_7;

Selector_2 s7569_7(wires_1892_6[1], addr_1892_6, addr_positional[30279:30276], addr_7569_7);

wire[31:0] addr_7570_7;

Selector_2 s7570_7(wires_1892_6[2], addr_1892_6, addr_positional[30283:30280], addr_7570_7);

wire[31:0] addr_7571_7;

Selector_2 s7571_7(wires_1892_6[3], addr_1892_6, addr_positional[30287:30284], addr_7571_7);

wire[31:0] addr_7572_7;

Selector_2 s7572_7(wires_1893_6[0], addr_1893_6, addr_positional[30291:30288], addr_7572_7);

wire[31:0] addr_7573_7;

Selector_2 s7573_7(wires_1893_6[1], addr_1893_6, addr_positional[30295:30292], addr_7573_7);

wire[31:0] addr_7574_7;

Selector_2 s7574_7(wires_1893_6[2], addr_1893_6, addr_positional[30299:30296], addr_7574_7);

wire[31:0] addr_7575_7;

Selector_2 s7575_7(wires_1893_6[3], addr_1893_6, addr_positional[30303:30300], addr_7575_7);

wire[31:0] addr_7576_7;

Selector_2 s7576_7(wires_1894_6[0], addr_1894_6, addr_positional[30307:30304], addr_7576_7);

wire[31:0] addr_7577_7;

Selector_2 s7577_7(wires_1894_6[1], addr_1894_6, addr_positional[30311:30308], addr_7577_7);

wire[31:0] addr_7578_7;

Selector_2 s7578_7(wires_1894_6[2], addr_1894_6, addr_positional[30315:30312], addr_7578_7);

wire[31:0] addr_7579_7;

Selector_2 s7579_7(wires_1894_6[3], addr_1894_6, addr_positional[30319:30316], addr_7579_7);

wire[31:0] addr_7580_7;

Selector_2 s7580_7(wires_1895_6[0], addr_1895_6, addr_positional[30323:30320], addr_7580_7);

wire[31:0] addr_7581_7;

Selector_2 s7581_7(wires_1895_6[1], addr_1895_6, addr_positional[30327:30324], addr_7581_7);

wire[31:0] addr_7582_7;

Selector_2 s7582_7(wires_1895_6[2], addr_1895_6, addr_positional[30331:30328], addr_7582_7);

wire[31:0] addr_7583_7;

Selector_2 s7583_7(wires_1895_6[3], addr_1895_6, addr_positional[30335:30332], addr_7583_7);

wire[31:0] addr_7584_7;

Selector_2 s7584_7(wires_1896_6[0], addr_1896_6, addr_positional[30339:30336], addr_7584_7);

wire[31:0] addr_7585_7;

Selector_2 s7585_7(wires_1896_6[1], addr_1896_6, addr_positional[30343:30340], addr_7585_7);

wire[31:0] addr_7586_7;

Selector_2 s7586_7(wires_1896_6[2], addr_1896_6, addr_positional[30347:30344], addr_7586_7);

wire[31:0] addr_7587_7;

Selector_2 s7587_7(wires_1896_6[3], addr_1896_6, addr_positional[30351:30348], addr_7587_7);

wire[31:0] addr_7588_7;

Selector_2 s7588_7(wires_1897_6[0], addr_1897_6, addr_positional[30355:30352], addr_7588_7);

wire[31:0] addr_7589_7;

Selector_2 s7589_7(wires_1897_6[1], addr_1897_6, addr_positional[30359:30356], addr_7589_7);

wire[31:0] addr_7590_7;

Selector_2 s7590_7(wires_1897_6[2], addr_1897_6, addr_positional[30363:30360], addr_7590_7);

wire[31:0] addr_7591_7;

Selector_2 s7591_7(wires_1897_6[3], addr_1897_6, addr_positional[30367:30364], addr_7591_7);

wire[31:0] addr_7592_7;

Selector_2 s7592_7(wires_1898_6[0], addr_1898_6, addr_positional[30371:30368], addr_7592_7);

wire[31:0] addr_7593_7;

Selector_2 s7593_7(wires_1898_6[1], addr_1898_6, addr_positional[30375:30372], addr_7593_7);

wire[31:0] addr_7594_7;

Selector_2 s7594_7(wires_1898_6[2], addr_1898_6, addr_positional[30379:30376], addr_7594_7);

wire[31:0] addr_7595_7;

Selector_2 s7595_7(wires_1898_6[3], addr_1898_6, addr_positional[30383:30380], addr_7595_7);

wire[31:0] addr_7596_7;

Selector_2 s7596_7(wires_1899_6[0], addr_1899_6, addr_positional[30387:30384], addr_7596_7);

wire[31:0] addr_7597_7;

Selector_2 s7597_7(wires_1899_6[1], addr_1899_6, addr_positional[30391:30388], addr_7597_7);

wire[31:0] addr_7598_7;

Selector_2 s7598_7(wires_1899_6[2], addr_1899_6, addr_positional[30395:30392], addr_7598_7);

wire[31:0] addr_7599_7;

Selector_2 s7599_7(wires_1899_6[3], addr_1899_6, addr_positional[30399:30396], addr_7599_7);

wire[31:0] addr_7600_7;

Selector_2 s7600_7(wires_1900_6[0], addr_1900_6, addr_positional[30403:30400], addr_7600_7);

wire[31:0] addr_7601_7;

Selector_2 s7601_7(wires_1900_6[1], addr_1900_6, addr_positional[30407:30404], addr_7601_7);

wire[31:0] addr_7602_7;

Selector_2 s7602_7(wires_1900_6[2], addr_1900_6, addr_positional[30411:30408], addr_7602_7);

wire[31:0] addr_7603_7;

Selector_2 s7603_7(wires_1900_6[3], addr_1900_6, addr_positional[30415:30412], addr_7603_7);

wire[31:0] addr_7604_7;

Selector_2 s7604_7(wires_1901_6[0], addr_1901_6, addr_positional[30419:30416], addr_7604_7);

wire[31:0] addr_7605_7;

Selector_2 s7605_7(wires_1901_6[1], addr_1901_6, addr_positional[30423:30420], addr_7605_7);

wire[31:0] addr_7606_7;

Selector_2 s7606_7(wires_1901_6[2], addr_1901_6, addr_positional[30427:30424], addr_7606_7);

wire[31:0] addr_7607_7;

Selector_2 s7607_7(wires_1901_6[3], addr_1901_6, addr_positional[30431:30428], addr_7607_7);

wire[31:0] addr_7608_7;

Selector_2 s7608_7(wires_1902_6[0], addr_1902_6, addr_positional[30435:30432], addr_7608_7);

wire[31:0] addr_7609_7;

Selector_2 s7609_7(wires_1902_6[1], addr_1902_6, addr_positional[30439:30436], addr_7609_7);

wire[31:0] addr_7610_7;

Selector_2 s7610_7(wires_1902_6[2], addr_1902_6, addr_positional[30443:30440], addr_7610_7);

wire[31:0] addr_7611_7;

Selector_2 s7611_7(wires_1902_6[3], addr_1902_6, addr_positional[30447:30444], addr_7611_7);

wire[31:0] addr_7612_7;

Selector_2 s7612_7(wires_1903_6[0], addr_1903_6, addr_positional[30451:30448], addr_7612_7);

wire[31:0] addr_7613_7;

Selector_2 s7613_7(wires_1903_6[1], addr_1903_6, addr_positional[30455:30452], addr_7613_7);

wire[31:0] addr_7614_7;

Selector_2 s7614_7(wires_1903_6[2], addr_1903_6, addr_positional[30459:30456], addr_7614_7);

wire[31:0] addr_7615_7;

Selector_2 s7615_7(wires_1903_6[3], addr_1903_6, addr_positional[30463:30460], addr_7615_7);

wire[31:0] addr_7616_7;

Selector_2 s7616_7(wires_1904_6[0], addr_1904_6, addr_positional[30467:30464], addr_7616_7);

wire[31:0] addr_7617_7;

Selector_2 s7617_7(wires_1904_6[1], addr_1904_6, addr_positional[30471:30468], addr_7617_7);

wire[31:0] addr_7618_7;

Selector_2 s7618_7(wires_1904_6[2], addr_1904_6, addr_positional[30475:30472], addr_7618_7);

wire[31:0] addr_7619_7;

Selector_2 s7619_7(wires_1904_6[3], addr_1904_6, addr_positional[30479:30476], addr_7619_7);

wire[31:0] addr_7620_7;

Selector_2 s7620_7(wires_1905_6[0], addr_1905_6, addr_positional[30483:30480], addr_7620_7);

wire[31:0] addr_7621_7;

Selector_2 s7621_7(wires_1905_6[1], addr_1905_6, addr_positional[30487:30484], addr_7621_7);

wire[31:0] addr_7622_7;

Selector_2 s7622_7(wires_1905_6[2], addr_1905_6, addr_positional[30491:30488], addr_7622_7);

wire[31:0] addr_7623_7;

Selector_2 s7623_7(wires_1905_6[3], addr_1905_6, addr_positional[30495:30492], addr_7623_7);

wire[31:0] addr_7624_7;

Selector_2 s7624_7(wires_1906_6[0], addr_1906_6, addr_positional[30499:30496], addr_7624_7);

wire[31:0] addr_7625_7;

Selector_2 s7625_7(wires_1906_6[1], addr_1906_6, addr_positional[30503:30500], addr_7625_7);

wire[31:0] addr_7626_7;

Selector_2 s7626_7(wires_1906_6[2], addr_1906_6, addr_positional[30507:30504], addr_7626_7);

wire[31:0] addr_7627_7;

Selector_2 s7627_7(wires_1906_6[3], addr_1906_6, addr_positional[30511:30508], addr_7627_7);

wire[31:0] addr_7628_7;

Selector_2 s7628_7(wires_1907_6[0], addr_1907_6, addr_positional[30515:30512], addr_7628_7);

wire[31:0] addr_7629_7;

Selector_2 s7629_7(wires_1907_6[1], addr_1907_6, addr_positional[30519:30516], addr_7629_7);

wire[31:0] addr_7630_7;

Selector_2 s7630_7(wires_1907_6[2], addr_1907_6, addr_positional[30523:30520], addr_7630_7);

wire[31:0] addr_7631_7;

Selector_2 s7631_7(wires_1907_6[3], addr_1907_6, addr_positional[30527:30524], addr_7631_7);

wire[31:0] addr_7632_7;

Selector_2 s7632_7(wires_1908_6[0], addr_1908_6, addr_positional[30531:30528], addr_7632_7);

wire[31:0] addr_7633_7;

Selector_2 s7633_7(wires_1908_6[1], addr_1908_6, addr_positional[30535:30532], addr_7633_7);

wire[31:0] addr_7634_7;

Selector_2 s7634_7(wires_1908_6[2], addr_1908_6, addr_positional[30539:30536], addr_7634_7);

wire[31:0] addr_7635_7;

Selector_2 s7635_7(wires_1908_6[3], addr_1908_6, addr_positional[30543:30540], addr_7635_7);

wire[31:0] addr_7636_7;

Selector_2 s7636_7(wires_1909_6[0], addr_1909_6, addr_positional[30547:30544], addr_7636_7);

wire[31:0] addr_7637_7;

Selector_2 s7637_7(wires_1909_6[1], addr_1909_6, addr_positional[30551:30548], addr_7637_7);

wire[31:0] addr_7638_7;

Selector_2 s7638_7(wires_1909_6[2], addr_1909_6, addr_positional[30555:30552], addr_7638_7);

wire[31:0] addr_7639_7;

Selector_2 s7639_7(wires_1909_6[3], addr_1909_6, addr_positional[30559:30556], addr_7639_7);

wire[31:0] addr_7640_7;

Selector_2 s7640_7(wires_1910_6[0], addr_1910_6, addr_positional[30563:30560], addr_7640_7);

wire[31:0] addr_7641_7;

Selector_2 s7641_7(wires_1910_6[1], addr_1910_6, addr_positional[30567:30564], addr_7641_7);

wire[31:0] addr_7642_7;

Selector_2 s7642_7(wires_1910_6[2], addr_1910_6, addr_positional[30571:30568], addr_7642_7);

wire[31:0] addr_7643_7;

Selector_2 s7643_7(wires_1910_6[3], addr_1910_6, addr_positional[30575:30572], addr_7643_7);

wire[31:0] addr_7644_7;

Selector_2 s7644_7(wires_1911_6[0], addr_1911_6, addr_positional[30579:30576], addr_7644_7);

wire[31:0] addr_7645_7;

Selector_2 s7645_7(wires_1911_6[1], addr_1911_6, addr_positional[30583:30580], addr_7645_7);

wire[31:0] addr_7646_7;

Selector_2 s7646_7(wires_1911_6[2], addr_1911_6, addr_positional[30587:30584], addr_7646_7);

wire[31:0] addr_7647_7;

Selector_2 s7647_7(wires_1911_6[3], addr_1911_6, addr_positional[30591:30588], addr_7647_7);

wire[31:0] addr_7648_7;

Selector_2 s7648_7(wires_1912_6[0], addr_1912_6, addr_positional[30595:30592], addr_7648_7);

wire[31:0] addr_7649_7;

Selector_2 s7649_7(wires_1912_6[1], addr_1912_6, addr_positional[30599:30596], addr_7649_7);

wire[31:0] addr_7650_7;

Selector_2 s7650_7(wires_1912_6[2], addr_1912_6, addr_positional[30603:30600], addr_7650_7);

wire[31:0] addr_7651_7;

Selector_2 s7651_7(wires_1912_6[3], addr_1912_6, addr_positional[30607:30604], addr_7651_7);

wire[31:0] addr_7652_7;

Selector_2 s7652_7(wires_1913_6[0], addr_1913_6, addr_positional[30611:30608], addr_7652_7);

wire[31:0] addr_7653_7;

Selector_2 s7653_7(wires_1913_6[1], addr_1913_6, addr_positional[30615:30612], addr_7653_7);

wire[31:0] addr_7654_7;

Selector_2 s7654_7(wires_1913_6[2], addr_1913_6, addr_positional[30619:30616], addr_7654_7);

wire[31:0] addr_7655_7;

Selector_2 s7655_7(wires_1913_6[3], addr_1913_6, addr_positional[30623:30620], addr_7655_7);

wire[31:0] addr_7656_7;

Selector_2 s7656_7(wires_1914_6[0], addr_1914_6, addr_positional[30627:30624], addr_7656_7);

wire[31:0] addr_7657_7;

Selector_2 s7657_7(wires_1914_6[1], addr_1914_6, addr_positional[30631:30628], addr_7657_7);

wire[31:0] addr_7658_7;

Selector_2 s7658_7(wires_1914_6[2], addr_1914_6, addr_positional[30635:30632], addr_7658_7);

wire[31:0] addr_7659_7;

Selector_2 s7659_7(wires_1914_6[3], addr_1914_6, addr_positional[30639:30636], addr_7659_7);

wire[31:0] addr_7660_7;

Selector_2 s7660_7(wires_1915_6[0], addr_1915_6, addr_positional[30643:30640], addr_7660_7);

wire[31:0] addr_7661_7;

Selector_2 s7661_7(wires_1915_6[1], addr_1915_6, addr_positional[30647:30644], addr_7661_7);

wire[31:0] addr_7662_7;

Selector_2 s7662_7(wires_1915_6[2], addr_1915_6, addr_positional[30651:30648], addr_7662_7);

wire[31:0] addr_7663_7;

Selector_2 s7663_7(wires_1915_6[3], addr_1915_6, addr_positional[30655:30652], addr_7663_7);

wire[31:0] addr_7664_7;

Selector_2 s7664_7(wires_1916_6[0], addr_1916_6, addr_positional[30659:30656], addr_7664_7);

wire[31:0] addr_7665_7;

Selector_2 s7665_7(wires_1916_6[1], addr_1916_6, addr_positional[30663:30660], addr_7665_7);

wire[31:0] addr_7666_7;

Selector_2 s7666_7(wires_1916_6[2], addr_1916_6, addr_positional[30667:30664], addr_7666_7);

wire[31:0] addr_7667_7;

Selector_2 s7667_7(wires_1916_6[3], addr_1916_6, addr_positional[30671:30668], addr_7667_7);

wire[31:0] addr_7668_7;

Selector_2 s7668_7(wires_1917_6[0], addr_1917_6, addr_positional[30675:30672], addr_7668_7);

wire[31:0] addr_7669_7;

Selector_2 s7669_7(wires_1917_6[1], addr_1917_6, addr_positional[30679:30676], addr_7669_7);

wire[31:0] addr_7670_7;

Selector_2 s7670_7(wires_1917_6[2], addr_1917_6, addr_positional[30683:30680], addr_7670_7);

wire[31:0] addr_7671_7;

Selector_2 s7671_7(wires_1917_6[3], addr_1917_6, addr_positional[30687:30684], addr_7671_7);

wire[31:0] addr_7672_7;

Selector_2 s7672_7(wires_1918_6[0], addr_1918_6, addr_positional[30691:30688], addr_7672_7);

wire[31:0] addr_7673_7;

Selector_2 s7673_7(wires_1918_6[1], addr_1918_6, addr_positional[30695:30692], addr_7673_7);

wire[31:0] addr_7674_7;

Selector_2 s7674_7(wires_1918_6[2], addr_1918_6, addr_positional[30699:30696], addr_7674_7);

wire[31:0] addr_7675_7;

Selector_2 s7675_7(wires_1918_6[3], addr_1918_6, addr_positional[30703:30700], addr_7675_7);

wire[31:0] addr_7676_7;

Selector_2 s7676_7(wires_1919_6[0], addr_1919_6, addr_positional[30707:30704], addr_7676_7);

wire[31:0] addr_7677_7;

Selector_2 s7677_7(wires_1919_6[1], addr_1919_6, addr_positional[30711:30708], addr_7677_7);

wire[31:0] addr_7678_7;

Selector_2 s7678_7(wires_1919_6[2], addr_1919_6, addr_positional[30715:30712], addr_7678_7);

wire[31:0] addr_7679_7;

Selector_2 s7679_7(wires_1919_6[3], addr_1919_6, addr_positional[30719:30716], addr_7679_7);

wire[31:0] addr_7680_7;

Selector_2 s7680_7(wires_1920_6[0], addr_1920_6, addr_positional[30723:30720], addr_7680_7);

wire[31:0] addr_7681_7;

Selector_2 s7681_7(wires_1920_6[1], addr_1920_6, addr_positional[30727:30724], addr_7681_7);

wire[31:0] addr_7682_7;

Selector_2 s7682_7(wires_1920_6[2], addr_1920_6, addr_positional[30731:30728], addr_7682_7);

wire[31:0] addr_7683_7;

Selector_2 s7683_7(wires_1920_6[3], addr_1920_6, addr_positional[30735:30732], addr_7683_7);

wire[31:0] addr_7684_7;

Selector_2 s7684_7(wires_1921_6[0], addr_1921_6, addr_positional[30739:30736], addr_7684_7);

wire[31:0] addr_7685_7;

Selector_2 s7685_7(wires_1921_6[1], addr_1921_6, addr_positional[30743:30740], addr_7685_7);

wire[31:0] addr_7686_7;

Selector_2 s7686_7(wires_1921_6[2], addr_1921_6, addr_positional[30747:30744], addr_7686_7);

wire[31:0] addr_7687_7;

Selector_2 s7687_7(wires_1921_6[3], addr_1921_6, addr_positional[30751:30748], addr_7687_7);

wire[31:0] addr_7688_7;

Selector_2 s7688_7(wires_1922_6[0], addr_1922_6, addr_positional[30755:30752], addr_7688_7);

wire[31:0] addr_7689_7;

Selector_2 s7689_7(wires_1922_6[1], addr_1922_6, addr_positional[30759:30756], addr_7689_7);

wire[31:0] addr_7690_7;

Selector_2 s7690_7(wires_1922_6[2], addr_1922_6, addr_positional[30763:30760], addr_7690_7);

wire[31:0] addr_7691_7;

Selector_2 s7691_7(wires_1922_6[3], addr_1922_6, addr_positional[30767:30764], addr_7691_7);

wire[31:0] addr_7692_7;

Selector_2 s7692_7(wires_1923_6[0], addr_1923_6, addr_positional[30771:30768], addr_7692_7);

wire[31:0] addr_7693_7;

Selector_2 s7693_7(wires_1923_6[1], addr_1923_6, addr_positional[30775:30772], addr_7693_7);

wire[31:0] addr_7694_7;

Selector_2 s7694_7(wires_1923_6[2], addr_1923_6, addr_positional[30779:30776], addr_7694_7);

wire[31:0] addr_7695_7;

Selector_2 s7695_7(wires_1923_6[3], addr_1923_6, addr_positional[30783:30780], addr_7695_7);

wire[31:0] addr_7696_7;

Selector_2 s7696_7(wires_1924_6[0], addr_1924_6, addr_positional[30787:30784], addr_7696_7);

wire[31:0] addr_7697_7;

Selector_2 s7697_7(wires_1924_6[1], addr_1924_6, addr_positional[30791:30788], addr_7697_7);

wire[31:0] addr_7698_7;

Selector_2 s7698_7(wires_1924_6[2], addr_1924_6, addr_positional[30795:30792], addr_7698_7);

wire[31:0] addr_7699_7;

Selector_2 s7699_7(wires_1924_6[3], addr_1924_6, addr_positional[30799:30796], addr_7699_7);

wire[31:0] addr_7700_7;

Selector_2 s7700_7(wires_1925_6[0], addr_1925_6, addr_positional[30803:30800], addr_7700_7);

wire[31:0] addr_7701_7;

Selector_2 s7701_7(wires_1925_6[1], addr_1925_6, addr_positional[30807:30804], addr_7701_7);

wire[31:0] addr_7702_7;

Selector_2 s7702_7(wires_1925_6[2], addr_1925_6, addr_positional[30811:30808], addr_7702_7);

wire[31:0] addr_7703_7;

Selector_2 s7703_7(wires_1925_6[3], addr_1925_6, addr_positional[30815:30812], addr_7703_7);

wire[31:0] addr_7704_7;

Selector_2 s7704_7(wires_1926_6[0], addr_1926_6, addr_positional[30819:30816], addr_7704_7);

wire[31:0] addr_7705_7;

Selector_2 s7705_7(wires_1926_6[1], addr_1926_6, addr_positional[30823:30820], addr_7705_7);

wire[31:0] addr_7706_7;

Selector_2 s7706_7(wires_1926_6[2], addr_1926_6, addr_positional[30827:30824], addr_7706_7);

wire[31:0] addr_7707_7;

Selector_2 s7707_7(wires_1926_6[3], addr_1926_6, addr_positional[30831:30828], addr_7707_7);

wire[31:0] addr_7708_7;

Selector_2 s7708_7(wires_1927_6[0], addr_1927_6, addr_positional[30835:30832], addr_7708_7);

wire[31:0] addr_7709_7;

Selector_2 s7709_7(wires_1927_6[1], addr_1927_6, addr_positional[30839:30836], addr_7709_7);

wire[31:0] addr_7710_7;

Selector_2 s7710_7(wires_1927_6[2], addr_1927_6, addr_positional[30843:30840], addr_7710_7);

wire[31:0] addr_7711_7;

Selector_2 s7711_7(wires_1927_6[3], addr_1927_6, addr_positional[30847:30844], addr_7711_7);

wire[31:0] addr_7712_7;

Selector_2 s7712_7(wires_1928_6[0], addr_1928_6, addr_positional[30851:30848], addr_7712_7);

wire[31:0] addr_7713_7;

Selector_2 s7713_7(wires_1928_6[1], addr_1928_6, addr_positional[30855:30852], addr_7713_7);

wire[31:0] addr_7714_7;

Selector_2 s7714_7(wires_1928_6[2], addr_1928_6, addr_positional[30859:30856], addr_7714_7);

wire[31:0] addr_7715_7;

Selector_2 s7715_7(wires_1928_6[3], addr_1928_6, addr_positional[30863:30860], addr_7715_7);

wire[31:0] addr_7716_7;

Selector_2 s7716_7(wires_1929_6[0], addr_1929_6, addr_positional[30867:30864], addr_7716_7);

wire[31:0] addr_7717_7;

Selector_2 s7717_7(wires_1929_6[1], addr_1929_6, addr_positional[30871:30868], addr_7717_7);

wire[31:0] addr_7718_7;

Selector_2 s7718_7(wires_1929_6[2], addr_1929_6, addr_positional[30875:30872], addr_7718_7);

wire[31:0] addr_7719_7;

Selector_2 s7719_7(wires_1929_6[3], addr_1929_6, addr_positional[30879:30876], addr_7719_7);

wire[31:0] addr_7720_7;

Selector_2 s7720_7(wires_1930_6[0], addr_1930_6, addr_positional[30883:30880], addr_7720_7);

wire[31:0] addr_7721_7;

Selector_2 s7721_7(wires_1930_6[1], addr_1930_6, addr_positional[30887:30884], addr_7721_7);

wire[31:0] addr_7722_7;

Selector_2 s7722_7(wires_1930_6[2], addr_1930_6, addr_positional[30891:30888], addr_7722_7);

wire[31:0] addr_7723_7;

Selector_2 s7723_7(wires_1930_6[3], addr_1930_6, addr_positional[30895:30892], addr_7723_7);

wire[31:0] addr_7724_7;

Selector_2 s7724_7(wires_1931_6[0], addr_1931_6, addr_positional[30899:30896], addr_7724_7);

wire[31:0] addr_7725_7;

Selector_2 s7725_7(wires_1931_6[1], addr_1931_6, addr_positional[30903:30900], addr_7725_7);

wire[31:0] addr_7726_7;

Selector_2 s7726_7(wires_1931_6[2], addr_1931_6, addr_positional[30907:30904], addr_7726_7);

wire[31:0] addr_7727_7;

Selector_2 s7727_7(wires_1931_6[3], addr_1931_6, addr_positional[30911:30908], addr_7727_7);

wire[31:0] addr_7728_7;

Selector_2 s7728_7(wires_1932_6[0], addr_1932_6, addr_positional[30915:30912], addr_7728_7);

wire[31:0] addr_7729_7;

Selector_2 s7729_7(wires_1932_6[1], addr_1932_6, addr_positional[30919:30916], addr_7729_7);

wire[31:0] addr_7730_7;

Selector_2 s7730_7(wires_1932_6[2], addr_1932_6, addr_positional[30923:30920], addr_7730_7);

wire[31:0] addr_7731_7;

Selector_2 s7731_7(wires_1932_6[3], addr_1932_6, addr_positional[30927:30924], addr_7731_7);

wire[31:0] addr_7732_7;

Selector_2 s7732_7(wires_1933_6[0], addr_1933_6, addr_positional[30931:30928], addr_7732_7);

wire[31:0] addr_7733_7;

Selector_2 s7733_7(wires_1933_6[1], addr_1933_6, addr_positional[30935:30932], addr_7733_7);

wire[31:0] addr_7734_7;

Selector_2 s7734_7(wires_1933_6[2], addr_1933_6, addr_positional[30939:30936], addr_7734_7);

wire[31:0] addr_7735_7;

Selector_2 s7735_7(wires_1933_6[3], addr_1933_6, addr_positional[30943:30940], addr_7735_7);

wire[31:0] addr_7736_7;

Selector_2 s7736_7(wires_1934_6[0], addr_1934_6, addr_positional[30947:30944], addr_7736_7);

wire[31:0] addr_7737_7;

Selector_2 s7737_7(wires_1934_6[1], addr_1934_6, addr_positional[30951:30948], addr_7737_7);

wire[31:0] addr_7738_7;

Selector_2 s7738_7(wires_1934_6[2], addr_1934_6, addr_positional[30955:30952], addr_7738_7);

wire[31:0] addr_7739_7;

Selector_2 s7739_7(wires_1934_6[3], addr_1934_6, addr_positional[30959:30956], addr_7739_7);

wire[31:0] addr_7740_7;

Selector_2 s7740_7(wires_1935_6[0], addr_1935_6, addr_positional[30963:30960], addr_7740_7);

wire[31:0] addr_7741_7;

Selector_2 s7741_7(wires_1935_6[1], addr_1935_6, addr_positional[30967:30964], addr_7741_7);

wire[31:0] addr_7742_7;

Selector_2 s7742_7(wires_1935_6[2], addr_1935_6, addr_positional[30971:30968], addr_7742_7);

wire[31:0] addr_7743_7;

Selector_2 s7743_7(wires_1935_6[3], addr_1935_6, addr_positional[30975:30972], addr_7743_7);

wire[31:0] addr_7744_7;

Selector_2 s7744_7(wires_1936_6[0], addr_1936_6, addr_positional[30979:30976], addr_7744_7);

wire[31:0] addr_7745_7;

Selector_2 s7745_7(wires_1936_6[1], addr_1936_6, addr_positional[30983:30980], addr_7745_7);

wire[31:0] addr_7746_7;

Selector_2 s7746_7(wires_1936_6[2], addr_1936_6, addr_positional[30987:30984], addr_7746_7);

wire[31:0] addr_7747_7;

Selector_2 s7747_7(wires_1936_6[3], addr_1936_6, addr_positional[30991:30988], addr_7747_7);

wire[31:0] addr_7748_7;

Selector_2 s7748_7(wires_1937_6[0], addr_1937_6, addr_positional[30995:30992], addr_7748_7);

wire[31:0] addr_7749_7;

Selector_2 s7749_7(wires_1937_6[1], addr_1937_6, addr_positional[30999:30996], addr_7749_7);

wire[31:0] addr_7750_7;

Selector_2 s7750_7(wires_1937_6[2], addr_1937_6, addr_positional[31003:31000], addr_7750_7);

wire[31:0] addr_7751_7;

Selector_2 s7751_7(wires_1937_6[3], addr_1937_6, addr_positional[31007:31004], addr_7751_7);

wire[31:0] addr_7752_7;

Selector_2 s7752_7(wires_1938_6[0], addr_1938_6, addr_positional[31011:31008], addr_7752_7);

wire[31:0] addr_7753_7;

Selector_2 s7753_7(wires_1938_6[1], addr_1938_6, addr_positional[31015:31012], addr_7753_7);

wire[31:0] addr_7754_7;

Selector_2 s7754_7(wires_1938_6[2], addr_1938_6, addr_positional[31019:31016], addr_7754_7);

wire[31:0] addr_7755_7;

Selector_2 s7755_7(wires_1938_6[3], addr_1938_6, addr_positional[31023:31020], addr_7755_7);

wire[31:0] addr_7756_7;

Selector_2 s7756_7(wires_1939_6[0], addr_1939_6, addr_positional[31027:31024], addr_7756_7);

wire[31:0] addr_7757_7;

Selector_2 s7757_7(wires_1939_6[1], addr_1939_6, addr_positional[31031:31028], addr_7757_7);

wire[31:0] addr_7758_7;

Selector_2 s7758_7(wires_1939_6[2], addr_1939_6, addr_positional[31035:31032], addr_7758_7);

wire[31:0] addr_7759_7;

Selector_2 s7759_7(wires_1939_6[3], addr_1939_6, addr_positional[31039:31036], addr_7759_7);

wire[31:0] addr_7760_7;

Selector_2 s7760_7(wires_1940_6[0], addr_1940_6, addr_positional[31043:31040], addr_7760_7);

wire[31:0] addr_7761_7;

Selector_2 s7761_7(wires_1940_6[1], addr_1940_6, addr_positional[31047:31044], addr_7761_7);

wire[31:0] addr_7762_7;

Selector_2 s7762_7(wires_1940_6[2], addr_1940_6, addr_positional[31051:31048], addr_7762_7);

wire[31:0] addr_7763_7;

Selector_2 s7763_7(wires_1940_6[3], addr_1940_6, addr_positional[31055:31052], addr_7763_7);

wire[31:0] addr_7764_7;

Selector_2 s7764_7(wires_1941_6[0], addr_1941_6, addr_positional[31059:31056], addr_7764_7);

wire[31:0] addr_7765_7;

Selector_2 s7765_7(wires_1941_6[1], addr_1941_6, addr_positional[31063:31060], addr_7765_7);

wire[31:0] addr_7766_7;

Selector_2 s7766_7(wires_1941_6[2], addr_1941_6, addr_positional[31067:31064], addr_7766_7);

wire[31:0] addr_7767_7;

Selector_2 s7767_7(wires_1941_6[3], addr_1941_6, addr_positional[31071:31068], addr_7767_7);

wire[31:0] addr_7768_7;

Selector_2 s7768_7(wires_1942_6[0], addr_1942_6, addr_positional[31075:31072], addr_7768_7);

wire[31:0] addr_7769_7;

Selector_2 s7769_7(wires_1942_6[1], addr_1942_6, addr_positional[31079:31076], addr_7769_7);

wire[31:0] addr_7770_7;

Selector_2 s7770_7(wires_1942_6[2], addr_1942_6, addr_positional[31083:31080], addr_7770_7);

wire[31:0] addr_7771_7;

Selector_2 s7771_7(wires_1942_6[3], addr_1942_6, addr_positional[31087:31084], addr_7771_7);

wire[31:0] addr_7772_7;

Selector_2 s7772_7(wires_1943_6[0], addr_1943_6, addr_positional[31091:31088], addr_7772_7);

wire[31:0] addr_7773_7;

Selector_2 s7773_7(wires_1943_6[1], addr_1943_6, addr_positional[31095:31092], addr_7773_7);

wire[31:0] addr_7774_7;

Selector_2 s7774_7(wires_1943_6[2], addr_1943_6, addr_positional[31099:31096], addr_7774_7);

wire[31:0] addr_7775_7;

Selector_2 s7775_7(wires_1943_6[3], addr_1943_6, addr_positional[31103:31100], addr_7775_7);

wire[31:0] addr_7776_7;

Selector_2 s7776_7(wires_1944_6[0], addr_1944_6, addr_positional[31107:31104], addr_7776_7);

wire[31:0] addr_7777_7;

Selector_2 s7777_7(wires_1944_6[1], addr_1944_6, addr_positional[31111:31108], addr_7777_7);

wire[31:0] addr_7778_7;

Selector_2 s7778_7(wires_1944_6[2], addr_1944_6, addr_positional[31115:31112], addr_7778_7);

wire[31:0] addr_7779_7;

Selector_2 s7779_7(wires_1944_6[3], addr_1944_6, addr_positional[31119:31116], addr_7779_7);

wire[31:0] addr_7780_7;

Selector_2 s7780_7(wires_1945_6[0], addr_1945_6, addr_positional[31123:31120], addr_7780_7);

wire[31:0] addr_7781_7;

Selector_2 s7781_7(wires_1945_6[1], addr_1945_6, addr_positional[31127:31124], addr_7781_7);

wire[31:0] addr_7782_7;

Selector_2 s7782_7(wires_1945_6[2], addr_1945_6, addr_positional[31131:31128], addr_7782_7);

wire[31:0] addr_7783_7;

Selector_2 s7783_7(wires_1945_6[3], addr_1945_6, addr_positional[31135:31132], addr_7783_7);

wire[31:0] addr_7784_7;

Selector_2 s7784_7(wires_1946_6[0], addr_1946_6, addr_positional[31139:31136], addr_7784_7);

wire[31:0] addr_7785_7;

Selector_2 s7785_7(wires_1946_6[1], addr_1946_6, addr_positional[31143:31140], addr_7785_7);

wire[31:0] addr_7786_7;

Selector_2 s7786_7(wires_1946_6[2], addr_1946_6, addr_positional[31147:31144], addr_7786_7);

wire[31:0] addr_7787_7;

Selector_2 s7787_7(wires_1946_6[3], addr_1946_6, addr_positional[31151:31148], addr_7787_7);

wire[31:0] addr_7788_7;

Selector_2 s7788_7(wires_1947_6[0], addr_1947_6, addr_positional[31155:31152], addr_7788_7);

wire[31:0] addr_7789_7;

Selector_2 s7789_7(wires_1947_6[1], addr_1947_6, addr_positional[31159:31156], addr_7789_7);

wire[31:0] addr_7790_7;

Selector_2 s7790_7(wires_1947_6[2], addr_1947_6, addr_positional[31163:31160], addr_7790_7);

wire[31:0] addr_7791_7;

Selector_2 s7791_7(wires_1947_6[3], addr_1947_6, addr_positional[31167:31164], addr_7791_7);

wire[31:0] addr_7792_7;

Selector_2 s7792_7(wires_1948_6[0], addr_1948_6, addr_positional[31171:31168], addr_7792_7);

wire[31:0] addr_7793_7;

Selector_2 s7793_7(wires_1948_6[1], addr_1948_6, addr_positional[31175:31172], addr_7793_7);

wire[31:0] addr_7794_7;

Selector_2 s7794_7(wires_1948_6[2], addr_1948_6, addr_positional[31179:31176], addr_7794_7);

wire[31:0] addr_7795_7;

Selector_2 s7795_7(wires_1948_6[3], addr_1948_6, addr_positional[31183:31180], addr_7795_7);

wire[31:0] addr_7796_7;

Selector_2 s7796_7(wires_1949_6[0], addr_1949_6, addr_positional[31187:31184], addr_7796_7);

wire[31:0] addr_7797_7;

Selector_2 s7797_7(wires_1949_6[1], addr_1949_6, addr_positional[31191:31188], addr_7797_7);

wire[31:0] addr_7798_7;

Selector_2 s7798_7(wires_1949_6[2], addr_1949_6, addr_positional[31195:31192], addr_7798_7);

wire[31:0] addr_7799_7;

Selector_2 s7799_7(wires_1949_6[3], addr_1949_6, addr_positional[31199:31196], addr_7799_7);

wire[31:0] addr_7800_7;

Selector_2 s7800_7(wires_1950_6[0], addr_1950_6, addr_positional[31203:31200], addr_7800_7);

wire[31:0] addr_7801_7;

Selector_2 s7801_7(wires_1950_6[1], addr_1950_6, addr_positional[31207:31204], addr_7801_7);

wire[31:0] addr_7802_7;

Selector_2 s7802_7(wires_1950_6[2], addr_1950_6, addr_positional[31211:31208], addr_7802_7);

wire[31:0] addr_7803_7;

Selector_2 s7803_7(wires_1950_6[3], addr_1950_6, addr_positional[31215:31212], addr_7803_7);

wire[31:0] addr_7804_7;

Selector_2 s7804_7(wires_1951_6[0], addr_1951_6, addr_positional[31219:31216], addr_7804_7);

wire[31:0] addr_7805_7;

Selector_2 s7805_7(wires_1951_6[1], addr_1951_6, addr_positional[31223:31220], addr_7805_7);

wire[31:0] addr_7806_7;

Selector_2 s7806_7(wires_1951_6[2], addr_1951_6, addr_positional[31227:31224], addr_7806_7);

wire[31:0] addr_7807_7;

Selector_2 s7807_7(wires_1951_6[3], addr_1951_6, addr_positional[31231:31228], addr_7807_7);

wire[31:0] addr_7808_7;

Selector_2 s7808_7(wires_1952_6[0], addr_1952_6, addr_positional[31235:31232], addr_7808_7);

wire[31:0] addr_7809_7;

Selector_2 s7809_7(wires_1952_6[1], addr_1952_6, addr_positional[31239:31236], addr_7809_7);

wire[31:0] addr_7810_7;

Selector_2 s7810_7(wires_1952_6[2], addr_1952_6, addr_positional[31243:31240], addr_7810_7);

wire[31:0] addr_7811_7;

Selector_2 s7811_7(wires_1952_6[3], addr_1952_6, addr_positional[31247:31244], addr_7811_7);

wire[31:0] addr_7812_7;

Selector_2 s7812_7(wires_1953_6[0], addr_1953_6, addr_positional[31251:31248], addr_7812_7);

wire[31:0] addr_7813_7;

Selector_2 s7813_7(wires_1953_6[1], addr_1953_6, addr_positional[31255:31252], addr_7813_7);

wire[31:0] addr_7814_7;

Selector_2 s7814_7(wires_1953_6[2], addr_1953_6, addr_positional[31259:31256], addr_7814_7);

wire[31:0] addr_7815_7;

Selector_2 s7815_7(wires_1953_6[3], addr_1953_6, addr_positional[31263:31260], addr_7815_7);

wire[31:0] addr_7816_7;

Selector_2 s7816_7(wires_1954_6[0], addr_1954_6, addr_positional[31267:31264], addr_7816_7);

wire[31:0] addr_7817_7;

Selector_2 s7817_7(wires_1954_6[1], addr_1954_6, addr_positional[31271:31268], addr_7817_7);

wire[31:0] addr_7818_7;

Selector_2 s7818_7(wires_1954_6[2], addr_1954_6, addr_positional[31275:31272], addr_7818_7);

wire[31:0] addr_7819_7;

Selector_2 s7819_7(wires_1954_6[3], addr_1954_6, addr_positional[31279:31276], addr_7819_7);

wire[31:0] addr_7820_7;

Selector_2 s7820_7(wires_1955_6[0], addr_1955_6, addr_positional[31283:31280], addr_7820_7);

wire[31:0] addr_7821_7;

Selector_2 s7821_7(wires_1955_6[1], addr_1955_6, addr_positional[31287:31284], addr_7821_7);

wire[31:0] addr_7822_7;

Selector_2 s7822_7(wires_1955_6[2], addr_1955_6, addr_positional[31291:31288], addr_7822_7);

wire[31:0] addr_7823_7;

Selector_2 s7823_7(wires_1955_6[3], addr_1955_6, addr_positional[31295:31292], addr_7823_7);

wire[31:0] addr_7824_7;

Selector_2 s7824_7(wires_1956_6[0], addr_1956_6, addr_positional[31299:31296], addr_7824_7);

wire[31:0] addr_7825_7;

Selector_2 s7825_7(wires_1956_6[1], addr_1956_6, addr_positional[31303:31300], addr_7825_7);

wire[31:0] addr_7826_7;

Selector_2 s7826_7(wires_1956_6[2], addr_1956_6, addr_positional[31307:31304], addr_7826_7);

wire[31:0] addr_7827_7;

Selector_2 s7827_7(wires_1956_6[3], addr_1956_6, addr_positional[31311:31308], addr_7827_7);

wire[31:0] addr_7828_7;

Selector_2 s7828_7(wires_1957_6[0], addr_1957_6, addr_positional[31315:31312], addr_7828_7);

wire[31:0] addr_7829_7;

Selector_2 s7829_7(wires_1957_6[1], addr_1957_6, addr_positional[31319:31316], addr_7829_7);

wire[31:0] addr_7830_7;

Selector_2 s7830_7(wires_1957_6[2], addr_1957_6, addr_positional[31323:31320], addr_7830_7);

wire[31:0] addr_7831_7;

Selector_2 s7831_7(wires_1957_6[3], addr_1957_6, addr_positional[31327:31324], addr_7831_7);

wire[31:0] addr_7832_7;

Selector_2 s7832_7(wires_1958_6[0], addr_1958_6, addr_positional[31331:31328], addr_7832_7);

wire[31:0] addr_7833_7;

Selector_2 s7833_7(wires_1958_6[1], addr_1958_6, addr_positional[31335:31332], addr_7833_7);

wire[31:0] addr_7834_7;

Selector_2 s7834_7(wires_1958_6[2], addr_1958_6, addr_positional[31339:31336], addr_7834_7);

wire[31:0] addr_7835_7;

Selector_2 s7835_7(wires_1958_6[3], addr_1958_6, addr_positional[31343:31340], addr_7835_7);

wire[31:0] addr_7836_7;

Selector_2 s7836_7(wires_1959_6[0], addr_1959_6, addr_positional[31347:31344], addr_7836_7);

wire[31:0] addr_7837_7;

Selector_2 s7837_7(wires_1959_6[1], addr_1959_6, addr_positional[31351:31348], addr_7837_7);

wire[31:0] addr_7838_7;

Selector_2 s7838_7(wires_1959_6[2], addr_1959_6, addr_positional[31355:31352], addr_7838_7);

wire[31:0] addr_7839_7;

Selector_2 s7839_7(wires_1959_6[3], addr_1959_6, addr_positional[31359:31356], addr_7839_7);

wire[31:0] addr_7840_7;

Selector_2 s7840_7(wires_1960_6[0], addr_1960_6, addr_positional[31363:31360], addr_7840_7);

wire[31:0] addr_7841_7;

Selector_2 s7841_7(wires_1960_6[1], addr_1960_6, addr_positional[31367:31364], addr_7841_7);

wire[31:0] addr_7842_7;

Selector_2 s7842_7(wires_1960_6[2], addr_1960_6, addr_positional[31371:31368], addr_7842_7);

wire[31:0] addr_7843_7;

Selector_2 s7843_7(wires_1960_6[3], addr_1960_6, addr_positional[31375:31372], addr_7843_7);

wire[31:0] addr_7844_7;

Selector_2 s7844_7(wires_1961_6[0], addr_1961_6, addr_positional[31379:31376], addr_7844_7);

wire[31:0] addr_7845_7;

Selector_2 s7845_7(wires_1961_6[1], addr_1961_6, addr_positional[31383:31380], addr_7845_7);

wire[31:0] addr_7846_7;

Selector_2 s7846_7(wires_1961_6[2], addr_1961_6, addr_positional[31387:31384], addr_7846_7);

wire[31:0] addr_7847_7;

Selector_2 s7847_7(wires_1961_6[3], addr_1961_6, addr_positional[31391:31388], addr_7847_7);

wire[31:0] addr_7848_7;

Selector_2 s7848_7(wires_1962_6[0], addr_1962_6, addr_positional[31395:31392], addr_7848_7);

wire[31:0] addr_7849_7;

Selector_2 s7849_7(wires_1962_6[1], addr_1962_6, addr_positional[31399:31396], addr_7849_7);

wire[31:0] addr_7850_7;

Selector_2 s7850_7(wires_1962_6[2], addr_1962_6, addr_positional[31403:31400], addr_7850_7);

wire[31:0] addr_7851_7;

Selector_2 s7851_7(wires_1962_6[3], addr_1962_6, addr_positional[31407:31404], addr_7851_7);

wire[31:0] addr_7852_7;

Selector_2 s7852_7(wires_1963_6[0], addr_1963_6, addr_positional[31411:31408], addr_7852_7);

wire[31:0] addr_7853_7;

Selector_2 s7853_7(wires_1963_6[1], addr_1963_6, addr_positional[31415:31412], addr_7853_7);

wire[31:0] addr_7854_7;

Selector_2 s7854_7(wires_1963_6[2], addr_1963_6, addr_positional[31419:31416], addr_7854_7);

wire[31:0] addr_7855_7;

Selector_2 s7855_7(wires_1963_6[3], addr_1963_6, addr_positional[31423:31420], addr_7855_7);

wire[31:0] addr_7856_7;

Selector_2 s7856_7(wires_1964_6[0], addr_1964_6, addr_positional[31427:31424], addr_7856_7);

wire[31:0] addr_7857_7;

Selector_2 s7857_7(wires_1964_6[1], addr_1964_6, addr_positional[31431:31428], addr_7857_7);

wire[31:0] addr_7858_7;

Selector_2 s7858_7(wires_1964_6[2], addr_1964_6, addr_positional[31435:31432], addr_7858_7);

wire[31:0] addr_7859_7;

Selector_2 s7859_7(wires_1964_6[3], addr_1964_6, addr_positional[31439:31436], addr_7859_7);

wire[31:0] addr_7860_7;

Selector_2 s7860_7(wires_1965_6[0], addr_1965_6, addr_positional[31443:31440], addr_7860_7);

wire[31:0] addr_7861_7;

Selector_2 s7861_7(wires_1965_6[1], addr_1965_6, addr_positional[31447:31444], addr_7861_7);

wire[31:0] addr_7862_7;

Selector_2 s7862_7(wires_1965_6[2], addr_1965_6, addr_positional[31451:31448], addr_7862_7);

wire[31:0] addr_7863_7;

Selector_2 s7863_7(wires_1965_6[3], addr_1965_6, addr_positional[31455:31452], addr_7863_7);

wire[31:0] addr_7864_7;

Selector_2 s7864_7(wires_1966_6[0], addr_1966_6, addr_positional[31459:31456], addr_7864_7);

wire[31:0] addr_7865_7;

Selector_2 s7865_7(wires_1966_6[1], addr_1966_6, addr_positional[31463:31460], addr_7865_7);

wire[31:0] addr_7866_7;

Selector_2 s7866_7(wires_1966_6[2], addr_1966_6, addr_positional[31467:31464], addr_7866_7);

wire[31:0] addr_7867_7;

Selector_2 s7867_7(wires_1966_6[3], addr_1966_6, addr_positional[31471:31468], addr_7867_7);

wire[31:0] addr_7868_7;

Selector_2 s7868_7(wires_1967_6[0], addr_1967_6, addr_positional[31475:31472], addr_7868_7);

wire[31:0] addr_7869_7;

Selector_2 s7869_7(wires_1967_6[1], addr_1967_6, addr_positional[31479:31476], addr_7869_7);

wire[31:0] addr_7870_7;

Selector_2 s7870_7(wires_1967_6[2], addr_1967_6, addr_positional[31483:31480], addr_7870_7);

wire[31:0] addr_7871_7;

Selector_2 s7871_7(wires_1967_6[3], addr_1967_6, addr_positional[31487:31484], addr_7871_7);

wire[31:0] addr_7872_7;

Selector_2 s7872_7(wires_1968_6[0], addr_1968_6, addr_positional[31491:31488], addr_7872_7);

wire[31:0] addr_7873_7;

Selector_2 s7873_7(wires_1968_6[1], addr_1968_6, addr_positional[31495:31492], addr_7873_7);

wire[31:0] addr_7874_7;

Selector_2 s7874_7(wires_1968_6[2], addr_1968_6, addr_positional[31499:31496], addr_7874_7);

wire[31:0] addr_7875_7;

Selector_2 s7875_7(wires_1968_6[3], addr_1968_6, addr_positional[31503:31500], addr_7875_7);

wire[31:0] addr_7876_7;

Selector_2 s7876_7(wires_1969_6[0], addr_1969_6, addr_positional[31507:31504], addr_7876_7);

wire[31:0] addr_7877_7;

Selector_2 s7877_7(wires_1969_6[1], addr_1969_6, addr_positional[31511:31508], addr_7877_7);

wire[31:0] addr_7878_7;

Selector_2 s7878_7(wires_1969_6[2], addr_1969_6, addr_positional[31515:31512], addr_7878_7);

wire[31:0] addr_7879_7;

Selector_2 s7879_7(wires_1969_6[3], addr_1969_6, addr_positional[31519:31516], addr_7879_7);

wire[31:0] addr_7880_7;

Selector_2 s7880_7(wires_1970_6[0], addr_1970_6, addr_positional[31523:31520], addr_7880_7);

wire[31:0] addr_7881_7;

Selector_2 s7881_7(wires_1970_6[1], addr_1970_6, addr_positional[31527:31524], addr_7881_7);

wire[31:0] addr_7882_7;

Selector_2 s7882_7(wires_1970_6[2], addr_1970_6, addr_positional[31531:31528], addr_7882_7);

wire[31:0] addr_7883_7;

Selector_2 s7883_7(wires_1970_6[3], addr_1970_6, addr_positional[31535:31532], addr_7883_7);

wire[31:0] addr_7884_7;

Selector_2 s7884_7(wires_1971_6[0], addr_1971_6, addr_positional[31539:31536], addr_7884_7);

wire[31:0] addr_7885_7;

Selector_2 s7885_7(wires_1971_6[1], addr_1971_6, addr_positional[31543:31540], addr_7885_7);

wire[31:0] addr_7886_7;

Selector_2 s7886_7(wires_1971_6[2], addr_1971_6, addr_positional[31547:31544], addr_7886_7);

wire[31:0] addr_7887_7;

Selector_2 s7887_7(wires_1971_6[3], addr_1971_6, addr_positional[31551:31548], addr_7887_7);

wire[31:0] addr_7888_7;

Selector_2 s7888_7(wires_1972_6[0], addr_1972_6, addr_positional[31555:31552], addr_7888_7);

wire[31:0] addr_7889_7;

Selector_2 s7889_7(wires_1972_6[1], addr_1972_6, addr_positional[31559:31556], addr_7889_7);

wire[31:0] addr_7890_7;

Selector_2 s7890_7(wires_1972_6[2], addr_1972_6, addr_positional[31563:31560], addr_7890_7);

wire[31:0] addr_7891_7;

Selector_2 s7891_7(wires_1972_6[3], addr_1972_6, addr_positional[31567:31564], addr_7891_7);

wire[31:0] addr_7892_7;

Selector_2 s7892_7(wires_1973_6[0], addr_1973_6, addr_positional[31571:31568], addr_7892_7);

wire[31:0] addr_7893_7;

Selector_2 s7893_7(wires_1973_6[1], addr_1973_6, addr_positional[31575:31572], addr_7893_7);

wire[31:0] addr_7894_7;

Selector_2 s7894_7(wires_1973_6[2], addr_1973_6, addr_positional[31579:31576], addr_7894_7);

wire[31:0] addr_7895_7;

Selector_2 s7895_7(wires_1973_6[3], addr_1973_6, addr_positional[31583:31580], addr_7895_7);

wire[31:0] addr_7896_7;

Selector_2 s7896_7(wires_1974_6[0], addr_1974_6, addr_positional[31587:31584], addr_7896_7);

wire[31:0] addr_7897_7;

Selector_2 s7897_7(wires_1974_6[1], addr_1974_6, addr_positional[31591:31588], addr_7897_7);

wire[31:0] addr_7898_7;

Selector_2 s7898_7(wires_1974_6[2], addr_1974_6, addr_positional[31595:31592], addr_7898_7);

wire[31:0] addr_7899_7;

Selector_2 s7899_7(wires_1974_6[3], addr_1974_6, addr_positional[31599:31596], addr_7899_7);

wire[31:0] addr_7900_7;

Selector_2 s7900_7(wires_1975_6[0], addr_1975_6, addr_positional[31603:31600], addr_7900_7);

wire[31:0] addr_7901_7;

Selector_2 s7901_7(wires_1975_6[1], addr_1975_6, addr_positional[31607:31604], addr_7901_7);

wire[31:0] addr_7902_7;

Selector_2 s7902_7(wires_1975_6[2], addr_1975_6, addr_positional[31611:31608], addr_7902_7);

wire[31:0] addr_7903_7;

Selector_2 s7903_7(wires_1975_6[3], addr_1975_6, addr_positional[31615:31612], addr_7903_7);

wire[31:0] addr_7904_7;

Selector_2 s7904_7(wires_1976_6[0], addr_1976_6, addr_positional[31619:31616], addr_7904_7);

wire[31:0] addr_7905_7;

Selector_2 s7905_7(wires_1976_6[1], addr_1976_6, addr_positional[31623:31620], addr_7905_7);

wire[31:0] addr_7906_7;

Selector_2 s7906_7(wires_1976_6[2], addr_1976_6, addr_positional[31627:31624], addr_7906_7);

wire[31:0] addr_7907_7;

Selector_2 s7907_7(wires_1976_6[3], addr_1976_6, addr_positional[31631:31628], addr_7907_7);

wire[31:0] addr_7908_7;

Selector_2 s7908_7(wires_1977_6[0], addr_1977_6, addr_positional[31635:31632], addr_7908_7);

wire[31:0] addr_7909_7;

Selector_2 s7909_7(wires_1977_6[1], addr_1977_6, addr_positional[31639:31636], addr_7909_7);

wire[31:0] addr_7910_7;

Selector_2 s7910_7(wires_1977_6[2], addr_1977_6, addr_positional[31643:31640], addr_7910_7);

wire[31:0] addr_7911_7;

Selector_2 s7911_7(wires_1977_6[3], addr_1977_6, addr_positional[31647:31644], addr_7911_7);

wire[31:0] addr_7912_7;

Selector_2 s7912_7(wires_1978_6[0], addr_1978_6, addr_positional[31651:31648], addr_7912_7);

wire[31:0] addr_7913_7;

Selector_2 s7913_7(wires_1978_6[1], addr_1978_6, addr_positional[31655:31652], addr_7913_7);

wire[31:0] addr_7914_7;

Selector_2 s7914_7(wires_1978_6[2], addr_1978_6, addr_positional[31659:31656], addr_7914_7);

wire[31:0] addr_7915_7;

Selector_2 s7915_7(wires_1978_6[3], addr_1978_6, addr_positional[31663:31660], addr_7915_7);

wire[31:0] addr_7916_7;

Selector_2 s7916_7(wires_1979_6[0], addr_1979_6, addr_positional[31667:31664], addr_7916_7);

wire[31:0] addr_7917_7;

Selector_2 s7917_7(wires_1979_6[1], addr_1979_6, addr_positional[31671:31668], addr_7917_7);

wire[31:0] addr_7918_7;

Selector_2 s7918_7(wires_1979_6[2], addr_1979_6, addr_positional[31675:31672], addr_7918_7);

wire[31:0] addr_7919_7;

Selector_2 s7919_7(wires_1979_6[3], addr_1979_6, addr_positional[31679:31676], addr_7919_7);

wire[31:0] addr_7920_7;

Selector_2 s7920_7(wires_1980_6[0], addr_1980_6, addr_positional[31683:31680], addr_7920_7);

wire[31:0] addr_7921_7;

Selector_2 s7921_7(wires_1980_6[1], addr_1980_6, addr_positional[31687:31684], addr_7921_7);

wire[31:0] addr_7922_7;

Selector_2 s7922_7(wires_1980_6[2], addr_1980_6, addr_positional[31691:31688], addr_7922_7);

wire[31:0] addr_7923_7;

Selector_2 s7923_7(wires_1980_6[3], addr_1980_6, addr_positional[31695:31692], addr_7923_7);

wire[31:0] addr_7924_7;

Selector_2 s7924_7(wires_1981_6[0], addr_1981_6, addr_positional[31699:31696], addr_7924_7);

wire[31:0] addr_7925_7;

Selector_2 s7925_7(wires_1981_6[1], addr_1981_6, addr_positional[31703:31700], addr_7925_7);

wire[31:0] addr_7926_7;

Selector_2 s7926_7(wires_1981_6[2], addr_1981_6, addr_positional[31707:31704], addr_7926_7);

wire[31:0] addr_7927_7;

Selector_2 s7927_7(wires_1981_6[3], addr_1981_6, addr_positional[31711:31708], addr_7927_7);

wire[31:0] addr_7928_7;

Selector_2 s7928_7(wires_1982_6[0], addr_1982_6, addr_positional[31715:31712], addr_7928_7);

wire[31:0] addr_7929_7;

Selector_2 s7929_7(wires_1982_6[1], addr_1982_6, addr_positional[31719:31716], addr_7929_7);

wire[31:0] addr_7930_7;

Selector_2 s7930_7(wires_1982_6[2], addr_1982_6, addr_positional[31723:31720], addr_7930_7);

wire[31:0] addr_7931_7;

Selector_2 s7931_7(wires_1982_6[3], addr_1982_6, addr_positional[31727:31724], addr_7931_7);

wire[31:0] addr_7932_7;

Selector_2 s7932_7(wires_1983_6[0], addr_1983_6, addr_positional[31731:31728], addr_7932_7);

wire[31:0] addr_7933_7;

Selector_2 s7933_7(wires_1983_6[1], addr_1983_6, addr_positional[31735:31732], addr_7933_7);

wire[31:0] addr_7934_7;

Selector_2 s7934_7(wires_1983_6[2], addr_1983_6, addr_positional[31739:31736], addr_7934_7);

wire[31:0] addr_7935_7;

Selector_2 s7935_7(wires_1983_6[3], addr_1983_6, addr_positional[31743:31740], addr_7935_7);

wire[31:0] addr_7936_7;

Selector_2 s7936_7(wires_1984_6[0], addr_1984_6, addr_positional[31747:31744], addr_7936_7);

wire[31:0] addr_7937_7;

Selector_2 s7937_7(wires_1984_6[1], addr_1984_6, addr_positional[31751:31748], addr_7937_7);

wire[31:0] addr_7938_7;

Selector_2 s7938_7(wires_1984_6[2], addr_1984_6, addr_positional[31755:31752], addr_7938_7);

wire[31:0] addr_7939_7;

Selector_2 s7939_7(wires_1984_6[3], addr_1984_6, addr_positional[31759:31756], addr_7939_7);

wire[31:0] addr_7940_7;

Selector_2 s7940_7(wires_1985_6[0], addr_1985_6, addr_positional[31763:31760], addr_7940_7);

wire[31:0] addr_7941_7;

Selector_2 s7941_7(wires_1985_6[1], addr_1985_6, addr_positional[31767:31764], addr_7941_7);

wire[31:0] addr_7942_7;

Selector_2 s7942_7(wires_1985_6[2], addr_1985_6, addr_positional[31771:31768], addr_7942_7);

wire[31:0] addr_7943_7;

Selector_2 s7943_7(wires_1985_6[3], addr_1985_6, addr_positional[31775:31772], addr_7943_7);

wire[31:0] addr_7944_7;

Selector_2 s7944_7(wires_1986_6[0], addr_1986_6, addr_positional[31779:31776], addr_7944_7);

wire[31:0] addr_7945_7;

Selector_2 s7945_7(wires_1986_6[1], addr_1986_6, addr_positional[31783:31780], addr_7945_7);

wire[31:0] addr_7946_7;

Selector_2 s7946_7(wires_1986_6[2], addr_1986_6, addr_positional[31787:31784], addr_7946_7);

wire[31:0] addr_7947_7;

Selector_2 s7947_7(wires_1986_6[3], addr_1986_6, addr_positional[31791:31788], addr_7947_7);

wire[31:0] addr_7948_7;

Selector_2 s7948_7(wires_1987_6[0], addr_1987_6, addr_positional[31795:31792], addr_7948_7);

wire[31:0] addr_7949_7;

Selector_2 s7949_7(wires_1987_6[1], addr_1987_6, addr_positional[31799:31796], addr_7949_7);

wire[31:0] addr_7950_7;

Selector_2 s7950_7(wires_1987_6[2], addr_1987_6, addr_positional[31803:31800], addr_7950_7);

wire[31:0] addr_7951_7;

Selector_2 s7951_7(wires_1987_6[3], addr_1987_6, addr_positional[31807:31804], addr_7951_7);

wire[31:0] addr_7952_7;

Selector_2 s7952_7(wires_1988_6[0], addr_1988_6, addr_positional[31811:31808], addr_7952_7);

wire[31:0] addr_7953_7;

Selector_2 s7953_7(wires_1988_6[1], addr_1988_6, addr_positional[31815:31812], addr_7953_7);

wire[31:0] addr_7954_7;

Selector_2 s7954_7(wires_1988_6[2], addr_1988_6, addr_positional[31819:31816], addr_7954_7);

wire[31:0] addr_7955_7;

Selector_2 s7955_7(wires_1988_6[3], addr_1988_6, addr_positional[31823:31820], addr_7955_7);

wire[31:0] addr_7956_7;

Selector_2 s7956_7(wires_1989_6[0], addr_1989_6, addr_positional[31827:31824], addr_7956_7);

wire[31:0] addr_7957_7;

Selector_2 s7957_7(wires_1989_6[1], addr_1989_6, addr_positional[31831:31828], addr_7957_7);

wire[31:0] addr_7958_7;

Selector_2 s7958_7(wires_1989_6[2], addr_1989_6, addr_positional[31835:31832], addr_7958_7);

wire[31:0] addr_7959_7;

Selector_2 s7959_7(wires_1989_6[3], addr_1989_6, addr_positional[31839:31836], addr_7959_7);

wire[31:0] addr_7960_7;

Selector_2 s7960_7(wires_1990_6[0], addr_1990_6, addr_positional[31843:31840], addr_7960_7);

wire[31:0] addr_7961_7;

Selector_2 s7961_7(wires_1990_6[1], addr_1990_6, addr_positional[31847:31844], addr_7961_7);

wire[31:0] addr_7962_7;

Selector_2 s7962_7(wires_1990_6[2], addr_1990_6, addr_positional[31851:31848], addr_7962_7);

wire[31:0] addr_7963_7;

Selector_2 s7963_7(wires_1990_6[3], addr_1990_6, addr_positional[31855:31852], addr_7963_7);

wire[31:0] addr_7964_7;

Selector_2 s7964_7(wires_1991_6[0], addr_1991_6, addr_positional[31859:31856], addr_7964_7);

wire[31:0] addr_7965_7;

Selector_2 s7965_7(wires_1991_6[1], addr_1991_6, addr_positional[31863:31860], addr_7965_7);

wire[31:0] addr_7966_7;

Selector_2 s7966_7(wires_1991_6[2], addr_1991_6, addr_positional[31867:31864], addr_7966_7);

wire[31:0] addr_7967_7;

Selector_2 s7967_7(wires_1991_6[3], addr_1991_6, addr_positional[31871:31868], addr_7967_7);

wire[31:0] addr_7968_7;

Selector_2 s7968_7(wires_1992_6[0], addr_1992_6, addr_positional[31875:31872], addr_7968_7);

wire[31:0] addr_7969_7;

Selector_2 s7969_7(wires_1992_6[1], addr_1992_6, addr_positional[31879:31876], addr_7969_7);

wire[31:0] addr_7970_7;

Selector_2 s7970_7(wires_1992_6[2], addr_1992_6, addr_positional[31883:31880], addr_7970_7);

wire[31:0] addr_7971_7;

Selector_2 s7971_7(wires_1992_6[3], addr_1992_6, addr_positional[31887:31884], addr_7971_7);

wire[31:0] addr_7972_7;

Selector_2 s7972_7(wires_1993_6[0], addr_1993_6, addr_positional[31891:31888], addr_7972_7);

wire[31:0] addr_7973_7;

Selector_2 s7973_7(wires_1993_6[1], addr_1993_6, addr_positional[31895:31892], addr_7973_7);

wire[31:0] addr_7974_7;

Selector_2 s7974_7(wires_1993_6[2], addr_1993_6, addr_positional[31899:31896], addr_7974_7);

wire[31:0] addr_7975_7;

Selector_2 s7975_7(wires_1993_6[3], addr_1993_6, addr_positional[31903:31900], addr_7975_7);

wire[31:0] addr_7976_7;

Selector_2 s7976_7(wires_1994_6[0], addr_1994_6, addr_positional[31907:31904], addr_7976_7);

wire[31:0] addr_7977_7;

Selector_2 s7977_7(wires_1994_6[1], addr_1994_6, addr_positional[31911:31908], addr_7977_7);

wire[31:0] addr_7978_7;

Selector_2 s7978_7(wires_1994_6[2], addr_1994_6, addr_positional[31915:31912], addr_7978_7);

wire[31:0] addr_7979_7;

Selector_2 s7979_7(wires_1994_6[3], addr_1994_6, addr_positional[31919:31916], addr_7979_7);

wire[31:0] addr_7980_7;

Selector_2 s7980_7(wires_1995_6[0], addr_1995_6, addr_positional[31923:31920], addr_7980_7);

wire[31:0] addr_7981_7;

Selector_2 s7981_7(wires_1995_6[1], addr_1995_6, addr_positional[31927:31924], addr_7981_7);

wire[31:0] addr_7982_7;

Selector_2 s7982_7(wires_1995_6[2], addr_1995_6, addr_positional[31931:31928], addr_7982_7);

wire[31:0] addr_7983_7;

Selector_2 s7983_7(wires_1995_6[3], addr_1995_6, addr_positional[31935:31932], addr_7983_7);

wire[31:0] addr_7984_7;

Selector_2 s7984_7(wires_1996_6[0], addr_1996_6, addr_positional[31939:31936], addr_7984_7);

wire[31:0] addr_7985_7;

Selector_2 s7985_7(wires_1996_6[1], addr_1996_6, addr_positional[31943:31940], addr_7985_7);

wire[31:0] addr_7986_7;

Selector_2 s7986_7(wires_1996_6[2], addr_1996_6, addr_positional[31947:31944], addr_7986_7);

wire[31:0] addr_7987_7;

Selector_2 s7987_7(wires_1996_6[3], addr_1996_6, addr_positional[31951:31948], addr_7987_7);

wire[31:0] addr_7988_7;

Selector_2 s7988_7(wires_1997_6[0], addr_1997_6, addr_positional[31955:31952], addr_7988_7);

wire[31:0] addr_7989_7;

Selector_2 s7989_7(wires_1997_6[1], addr_1997_6, addr_positional[31959:31956], addr_7989_7);

wire[31:0] addr_7990_7;

Selector_2 s7990_7(wires_1997_6[2], addr_1997_6, addr_positional[31963:31960], addr_7990_7);

wire[31:0] addr_7991_7;

Selector_2 s7991_7(wires_1997_6[3], addr_1997_6, addr_positional[31967:31964], addr_7991_7);

wire[31:0] addr_7992_7;

Selector_2 s7992_7(wires_1998_6[0], addr_1998_6, addr_positional[31971:31968], addr_7992_7);

wire[31:0] addr_7993_7;

Selector_2 s7993_7(wires_1998_6[1], addr_1998_6, addr_positional[31975:31972], addr_7993_7);

wire[31:0] addr_7994_7;

Selector_2 s7994_7(wires_1998_6[2], addr_1998_6, addr_positional[31979:31976], addr_7994_7);

wire[31:0] addr_7995_7;

Selector_2 s7995_7(wires_1998_6[3], addr_1998_6, addr_positional[31983:31980], addr_7995_7);

wire[31:0] addr_7996_7;

Selector_2 s7996_7(wires_1999_6[0], addr_1999_6, addr_positional[31987:31984], addr_7996_7);

wire[31:0] addr_7997_7;

Selector_2 s7997_7(wires_1999_6[1], addr_1999_6, addr_positional[31991:31988], addr_7997_7);

wire[31:0] addr_7998_7;

Selector_2 s7998_7(wires_1999_6[2], addr_1999_6, addr_positional[31995:31992], addr_7998_7);

wire[31:0] addr_7999_7;

Selector_2 s7999_7(wires_1999_6[3], addr_1999_6, addr_positional[31999:31996], addr_7999_7);

wire[31:0] addr_8000_7;

Selector_2 s8000_7(wires_2000_6[0], addr_2000_6, addr_positional[32003:32000], addr_8000_7);

wire[31:0] addr_8001_7;

Selector_2 s8001_7(wires_2000_6[1], addr_2000_6, addr_positional[32007:32004], addr_8001_7);

wire[31:0] addr_8002_7;

Selector_2 s8002_7(wires_2000_6[2], addr_2000_6, addr_positional[32011:32008], addr_8002_7);

wire[31:0] addr_8003_7;

Selector_2 s8003_7(wires_2000_6[3], addr_2000_6, addr_positional[32015:32012], addr_8003_7);

wire[31:0] addr_8004_7;

Selector_2 s8004_7(wires_2001_6[0], addr_2001_6, addr_positional[32019:32016], addr_8004_7);

wire[31:0] addr_8005_7;

Selector_2 s8005_7(wires_2001_6[1], addr_2001_6, addr_positional[32023:32020], addr_8005_7);

wire[31:0] addr_8006_7;

Selector_2 s8006_7(wires_2001_6[2], addr_2001_6, addr_positional[32027:32024], addr_8006_7);

wire[31:0] addr_8007_7;

Selector_2 s8007_7(wires_2001_6[3], addr_2001_6, addr_positional[32031:32028], addr_8007_7);

wire[31:0] addr_8008_7;

Selector_2 s8008_7(wires_2002_6[0], addr_2002_6, addr_positional[32035:32032], addr_8008_7);

wire[31:0] addr_8009_7;

Selector_2 s8009_7(wires_2002_6[1], addr_2002_6, addr_positional[32039:32036], addr_8009_7);

wire[31:0] addr_8010_7;

Selector_2 s8010_7(wires_2002_6[2], addr_2002_6, addr_positional[32043:32040], addr_8010_7);

wire[31:0] addr_8011_7;

Selector_2 s8011_7(wires_2002_6[3], addr_2002_6, addr_positional[32047:32044], addr_8011_7);

wire[31:0] addr_8012_7;

Selector_2 s8012_7(wires_2003_6[0], addr_2003_6, addr_positional[32051:32048], addr_8012_7);

wire[31:0] addr_8013_7;

Selector_2 s8013_7(wires_2003_6[1], addr_2003_6, addr_positional[32055:32052], addr_8013_7);

wire[31:0] addr_8014_7;

Selector_2 s8014_7(wires_2003_6[2], addr_2003_6, addr_positional[32059:32056], addr_8014_7);

wire[31:0] addr_8015_7;

Selector_2 s8015_7(wires_2003_6[3], addr_2003_6, addr_positional[32063:32060], addr_8015_7);

wire[31:0] addr_8016_7;

Selector_2 s8016_7(wires_2004_6[0], addr_2004_6, addr_positional[32067:32064], addr_8016_7);

wire[31:0] addr_8017_7;

Selector_2 s8017_7(wires_2004_6[1], addr_2004_6, addr_positional[32071:32068], addr_8017_7);

wire[31:0] addr_8018_7;

Selector_2 s8018_7(wires_2004_6[2], addr_2004_6, addr_positional[32075:32072], addr_8018_7);

wire[31:0] addr_8019_7;

Selector_2 s8019_7(wires_2004_6[3], addr_2004_6, addr_positional[32079:32076], addr_8019_7);

wire[31:0] addr_8020_7;

Selector_2 s8020_7(wires_2005_6[0], addr_2005_6, addr_positional[32083:32080], addr_8020_7);

wire[31:0] addr_8021_7;

Selector_2 s8021_7(wires_2005_6[1], addr_2005_6, addr_positional[32087:32084], addr_8021_7);

wire[31:0] addr_8022_7;

Selector_2 s8022_7(wires_2005_6[2], addr_2005_6, addr_positional[32091:32088], addr_8022_7);

wire[31:0] addr_8023_7;

Selector_2 s8023_7(wires_2005_6[3], addr_2005_6, addr_positional[32095:32092], addr_8023_7);

wire[31:0] addr_8024_7;

Selector_2 s8024_7(wires_2006_6[0], addr_2006_6, addr_positional[32099:32096], addr_8024_7);

wire[31:0] addr_8025_7;

Selector_2 s8025_7(wires_2006_6[1], addr_2006_6, addr_positional[32103:32100], addr_8025_7);

wire[31:0] addr_8026_7;

Selector_2 s8026_7(wires_2006_6[2], addr_2006_6, addr_positional[32107:32104], addr_8026_7);

wire[31:0] addr_8027_7;

Selector_2 s8027_7(wires_2006_6[3], addr_2006_6, addr_positional[32111:32108], addr_8027_7);

wire[31:0] addr_8028_7;

Selector_2 s8028_7(wires_2007_6[0], addr_2007_6, addr_positional[32115:32112], addr_8028_7);

wire[31:0] addr_8029_7;

Selector_2 s8029_7(wires_2007_6[1], addr_2007_6, addr_positional[32119:32116], addr_8029_7);

wire[31:0] addr_8030_7;

Selector_2 s8030_7(wires_2007_6[2], addr_2007_6, addr_positional[32123:32120], addr_8030_7);

wire[31:0] addr_8031_7;

Selector_2 s8031_7(wires_2007_6[3], addr_2007_6, addr_positional[32127:32124], addr_8031_7);

wire[31:0] addr_8032_7;

Selector_2 s8032_7(wires_2008_6[0], addr_2008_6, addr_positional[32131:32128], addr_8032_7);

wire[31:0] addr_8033_7;

Selector_2 s8033_7(wires_2008_6[1], addr_2008_6, addr_positional[32135:32132], addr_8033_7);

wire[31:0] addr_8034_7;

Selector_2 s8034_7(wires_2008_6[2], addr_2008_6, addr_positional[32139:32136], addr_8034_7);

wire[31:0] addr_8035_7;

Selector_2 s8035_7(wires_2008_6[3], addr_2008_6, addr_positional[32143:32140], addr_8035_7);

wire[31:0] addr_8036_7;

Selector_2 s8036_7(wires_2009_6[0], addr_2009_6, addr_positional[32147:32144], addr_8036_7);

wire[31:0] addr_8037_7;

Selector_2 s8037_7(wires_2009_6[1], addr_2009_6, addr_positional[32151:32148], addr_8037_7);

wire[31:0] addr_8038_7;

Selector_2 s8038_7(wires_2009_6[2], addr_2009_6, addr_positional[32155:32152], addr_8038_7);

wire[31:0] addr_8039_7;

Selector_2 s8039_7(wires_2009_6[3], addr_2009_6, addr_positional[32159:32156], addr_8039_7);

wire[31:0] addr_8040_7;

Selector_2 s8040_7(wires_2010_6[0], addr_2010_6, addr_positional[32163:32160], addr_8040_7);

wire[31:0] addr_8041_7;

Selector_2 s8041_7(wires_2010_6[1], addr_2010_6, addr_positional[32167:32164], addr_8041_7);

wire[31:0] addr_8042_7;

Selector_2 s8042_7(wires_2010_6[2], addr_2010_6, addr_positional[32171:32168], addr_8042_7);

wire[31:0] addr_8043_7;

Selector_2 s8043_7(wires_2010_6[3], addr_2010_6, addr_positional[32175:32172], addr_8043_7);

wire[31:0] addr_8044_7;

Selector_2 s8044_7(wires_2011_6[0], addr_2011_6, addr_positional[32179:32176], addr_8044_7);

wire[31:0] addr_8045_7;

Selector_2 s8045_7(wires_2011_6[1], addr_2011_6, addr_positional[32183:32180], addr_8045_7);

wire[31:0] addr_8046_7;

Selector_2 s8046_7(wires_2011_6[2], addr_2011_6, addr_positional[32187:32184], addr_8046_7);

wire[31:0] addr_8047_7;

Selector_2 s8047_7(wires_2011_6[3], addr_2011_6, addr_positional[32191:32188], addr_8047_7);

wire[31:0] addr_8048_7;

Selector_2 s8048_7(wires_2012_6[0], addr_2012_6, addr_positional[32195:32192], addr_8048_7);

wire[31:0] addr_8049_7;

Selector_2 s8049_7(wires_2012_6[1], addr_2012_6, addr_positional[32199:32196], addr_8049_7);

wire[31:0] addr_8050_7;

Selector_2 s8050_7(wires_2012_6[2], addr_2012_6, addr_positional[32203:32200], addr_8050_7);

wire[31:0] addr_8051_7;

Selector_2 s8051_7(wires_2012_6[3], addr_2012_6, addr_positional[32207:32204], addr_8051_7);

wire[31:0] addr_8052_7;

Selector_2 s8052_7(wires_2013_6[0], addr_2013_6, addr_positional[32211:32208], addr_8052_7);

wire[31:0] addr_8053_7;

Selector_2 s8053_7(wires_2013_6[1], addr_2013_6, addr_positional[32215:32212], addr_8053_7);

wire[31:0] addr_8054_7;

Selector_2 s8054_7(wires_2013_6[2], addr_2013_6, addr_positional[32219:32216], addr_8054_7);

wire[31:0] addr_8055_7;

Selector_2 s8055_7(wires_2013_6[3], addr_2013_6, addr_positional[32223:32220], addr_8055_7);

wire[31:0] addr_8056_7;

Selector_2 s8056_7(wires_2014_6[0], addr_2014_6, addr_positional[32227:32224], addr_8056_7);

wire[31:0] addr_8057_7;

Selector_2 s8057_7(wires_2014_6[1], addr_2014_6, addr_positional[32231:32228], addr_8057_7);

wire[31:0] addr_8058_7;

Selector_2 s8058_7(wires_2014_6[2], addr_2014_6, addr_positional[32235:32232], addr_8058_7);

wire[31:0] addr_8059_7;

Selector_2 s8059_7(wires_2014_6[3], addr_2014_6, addr_positional[32239:32236], addr_8059_7);

wire[31:0] addr_8060_7;

Selector_2 s8060_7(wires_2015_6[0], addr_2015_6, addr_positional[32243:32240], addr_8060_7);

wire[31:0] addr_8061_7;

Selector_2 s8061_7(wires_2015_6[1], addr_2015_6, addr_positional[32247:32244], addr_8061_7);

wire[31:0] addr_8062_7;

Selector_2 s8062_7(wires_2015_6[2], addr_2015_6, addr_positional[32251:32248], addr_8062_7);

wire[31:0] addr_8063_7;

Selector_2 s8063_7(wires_2015_6[3], addr_2015_6, addr_positional[32255:32252], addr_8063_7);

wire[31:0] addr_8064_7;

Selector_2 s8064_7(wires_2016_6[0], addr_2016_6, addr_positional[32259:32256], addr_8064_7);

wire[31:0] addr_8065_7;

Selector_2 s8065_7(wires_2016_6[1], addr_2016_6, addr_positional[32263:32260], addr_8065_7);

wire[31:0] addr_8066_7;

Selector_2 s8066_7(wires_2016_6[2], addr_2016_6, addr_positional[32267:32264], addr_8066_7);

wire[31:0] addr_8067_7;

Selector_2 s8067_7(wires_2016_6[3], addr_2016_6, addr_positional[32271:32268], addr_8067_7);

wire[31:0] addr_8068_7;

Selector_2 s8068_7(wires_2017_6[0], addr_2017_6, addr_positional[32275:32272], addr_8068_7);

wire[31:0] addr_8069_7;

Selector_2 s8069_7(wires_2017_6[1], addr_2017_6, addr_positional[32279:32276], addr_8069_7);

wire[31:0] addr_8070_7;

Selector_2 s8070_7(wires_2017_6[2], addr_2017_6, addr_positional[32283:32280], addr_8070_7);

wire[31:0] addr_8071_7;

Selector_2 s8071_7(wires_2017_6[3], addr_2017_6, addr_positional[32287:32284], addr_8071_7);

wire[31:0] addr_8072_7;

Selector_2 s8072_7(wires_2018_6[0], addr_2018_6, addr_positional[32291:32288], addr_8072_7);

wire[31:0] addr_8073_7;

Selector_2 s8073_7(wires_2018_6[1], addr_2018_6, addr_positional[32295:32292], addr_8073_7);

wire[31:0] addr_8074_7;

Selector_2 s8074_7(wires_2018_6[2], addr_2018_6, addr_positional[32299:32296], addr_8074_7);

wire[31:0] addr_8075_7;

Selector_2 s8075_7(wires_2018_6[3], addr_2018_6, addr_positional[32303:32300], addr_8075_7);

wire[31:0] addr_8076_7;

Selector_2 s8076_7(wires_2019_6[0], addr_2019_6, addr_positional[32307:32304], addr_8076_7);

wire[31:0] addr_8077_7;

Selector_2 s8077_7(wires_2019_6[1], addr_2019_6, addr_positional[32311:32308], addr_8077_7);

wire[31:0] addr_8078_7;

Selector_2 s8078_7(wires_2019_6[2], addr_2019_6, addr_positional[32315:32312], addr_8078_7);

wire[31:0] addr_8079_7;

Selector_2 s8079_7(wires_2019_6[3], addr_2019_6, addr_positional[32319:32316], addr_8079_7);

wire[31:0] addr_8080_7;

Selector_2 s8080_7(wires_2020_6[0], addr_2020_6, addr_positional[32323:32320], addr_8080_7);

wire[31:0] addr_8081_7;

Selector_2 s8081_7(wires_2020_6[1], addr_2020_6, addr_positional[32327:32324], addr_8081_7);

wire[31:0] addr_8082_7;

Selector_2 s8082_7(wires_2020_6[2], addr_2020_6, addr_positional[32331:32328], addr_8082_7);

wire[31:0] addr_8083_7;

Selector_2 s8083_7(wires_2020_6[3], addr_2020_6, addr_positional[32335:32332], addr_8083_7);

wire[31:0] addr_8084_7;

Selector_2 s8084_7(wires_2021_6[0], addr_2021_6, addr_positional[32339:32336], addr_8084_7);

wire[31:0] addr_8085_7;

Selector_2 s8085_7(wires_2021_6[1], addr_2021_6, addr_positional[32343:32340], addr_8085_7);

wire[31:0] addr_8086_7;

Selector_2 s8086_7(wires_2021_6[2], addr_2021_6, addr_positional[32347:32344], addr_8086_7);

wire[31:0] addr_8087_7;

Selector_2 s8087_7(wires_2021_6[3], addr_2021_6, addr_positional[32351:32348], addr_8087_7);

wire[31:0] addr_8088_7;

Selector_2 s8088_7(wires_2022_6[0], addr_2022_6, addr_positional[32355:32352], addr_8088_7);

wire[31:0] addr_8089_7;

Selector_2 s8089_7(wires_2022_6[1], addr_2022_6, addr_positional[32359:32356], addr_8089_7);

wire[31:0] addr_8090_7;

Selector_2 s8090_7(wires_2022_6[2], addr_2022_6, addr_positional[32363:32360], addr_8090_7);

wire[31:0] addr_8091_7;

Selector_2 s8091_7(wires_2022_6[3], addr_2022_6, addr_positional[32367:32364], addr_8091_7);

wire[31:0] addr_8092_7;

Selector_2 s8092_7(wires_2023_6[0], addr_2023_6, addr_positional[32371:32368], addr_8092_7);

wire[31:0] addr_8093_7;

Selector_2 s8093_7(wires_2023_6[1], addr_2023_6, addr_positional[32375:32372], addr_8093_7);

wire[31:0] addr_8094_7;

Selector_2 s8094_7(wires_2023_6[2], addr_2023_6, addr_positional[32379:32376], addr_8094_7);

wire[31:0] addr_8095_7;

Selector_2 s8095_7(wires_2023_6[3], addr_2023_6, addr_positional[32383:32380], addr_8095_7);

wire[31:0] addr_8096_7;

Selector_2 s8096_7(wires_2024_6[0], addr_2024_6, addr_positional[32387:32384], addr_8096_7);

wire[31:0] addr_8097_7;

Selector_2 s8097_7(wires_2024_6[1], addr_2024_6, addr_positional[32391:32388], addr_8097_7);

wire[31:0] addr_8098_7;

Selector_2 s8098_7(wires_2024_6[2], addr_2024_6, addr_positional[32395:32392], addr_8098_7);

wire[31:0] addr_8099_7;

Selector_2 s8099_7(wires_2024_6[3], addr_2024_6, addr_positional[32399:32396], addr_8099_7);

wire[31:0] addr_8100_7;

Selector_2 s8100_7(wires_2025_6[0], addr_2025_6, addr_positional[32403:32400], addr_8100_7);

wire[31:0] addr_8101_7;

Selector_2 s8101_7(wires_2025_6[1], addr_2025_6, addr_positional[32407:32404], addr_8101_7);

wire[31:0] addr_8102_7;

Selector_2 s8102_7(wires_2025_6[2], addr_2025_6, addr_positional[32411:32408], addr_8102_7);

wire[31:0] addr_8103_7;

Selector_2 s8103_7(wires_2025_6[3], addr_2025_6, addr_positional[32415:32412], addr_8103_7);

wire[31:0] addr_8104_7;

Selector_2 s8104_7(wires_2026_6[0], addr_2026_6, addr_positional[32419:32416], addr_8104_7);

wire[31:0] addr_8105_7;

Selector_2 s8105_7(wires_2026_6[1], addr_2026_6, addr_positional[32423:32420], addr_8105_7);

wire[31:0] addr_8106_7;

Selector_2 s8106_7(wires_2026_6[2], addr_2026_6, addr_positional[32427:32424], addr_8106_7);

wire[31:0] addr_8107_7;

Selector_2 s8107_7(wires_2026_6[3], addr_2026_6, addr_positional[32431:32428], addr_8107_7);

wire[31:0] addr_8108_7;

Selector_2 s8108_7(wires_2027_6[0], addr_2027_6, addr_positional[32435:32432], addr_8108_7);

wire[31:0] addr_8109_7;

Selector_2 s8109_7(wires_2027_6[1], addr_2027_6, addr_positional[32439:32436], addr_8109_7);

wire[31:0] addr_8110_7;

Selector_2 s8110_7(wires_2027_6[2], addr_2027_6, addr_positional[32443:32440], addr_8110_7);

wire[31:0] addr_8111_7;

Selector_2 s8111_7(wires_2027_6[3], addr_2027_6, addr_positional[32447:32444], addr_8111_7);

wire[31:0] addr_8112_7;

Selector_2 s8112_7(wires_2028_6[0], addr_2028_6, addr_positional[32451:32448], addr_8112_7);

wire[31:0] addr_8113_7;

Selector_2 s8113_7(wires_2028_6[1], addr_2028_6, addr_positional[32455:32452], addr_8113_7);

wire[31:0] addr_8114_7;

Selector_2 s8114_7(wires_2028_6[2], addr_2028_6, addr_positional[32459:32456], addr_8114_7);

wire[31:0] addr_8115_7;

Selector_2 s8115_7(wires_2028_6[3], addr_2028_6, addr_positional[32463:32460], addr_8115_7);

wire[31:0] addr_8116_7;

Selector_2 s8116_7(wires_2029_6[0], addr_2029_6, addr_positional[32467:32464], addr_8116_7);

wire[31:0] addr_8117_7;

Selector_2 s8117_7(wires_2029_6[1], addr_2029_6, addr_positional[32471:32468], addr_8117_7);

wire[31:0] addr_8118_7;

Selector_2 s8118_7(wires_2029_6[2], addr_2029_6, addr_positional[32475:32472], addr_8118_7);

wire[31:0] addr_8119_7;

Selector_2 s8119_7(wires_2029_6[3], addr_2029_6, addr_positional[32479:32476], addr_8119_7);

wire[31:0] addr_8120_7;

Selector_2 s8120_7(wires_2030_6[0], addr_2030_6, addr_positional[32483:32480], addr_8120_7);

wire[31:0] addr_8121_7;

Selector_2 s8121_7(wires_2030_6[1], addr_2030_6, addr_positional[32487:32484], addr_8121_7);

wire[31:0] addr_8122_7;

Selector_2 s8122_7(wires_2030_6[2], addr_2030_6, addr_positional[32491:32488], addr_8122_7);

wire[31:0] addr_8123_7;

Selector_2 s8123_7(wires_2030_6[3], addr_2030_6, addr_positional[32495:32492], addr_8123_7);

wire[31:0] addr_8124_7;

Selector_2 s8124_7(wires_2031_6[0], addr_2031_6, addr_positional[32499:32496], addr_8124_7);

wire[31:0] addr_8125_7;

Selector_2 s8125_7(wires_2031_6[1], addr_2031_6, addr_positional[32503:32500], addr_8125_7);

wire[31:0] addr_8126_7;

Selector_2 s8126_7(wires_2031_6[2], addr_2031_6, addr_positional[32507:32504], addr_8126_7);

wire[31:0] addr_8127_7;

Selector_2 s8127_7(wires_2031_6[3], addr_2031_6, addr_positional[32511:32508], addr_8127_7);

wire[31:0] addr_8128_7;

Selector_2 s8128_7(wires_2032_6[0], addr_2032_6, addr_positional[32515:32512], addr_8128_7);

wire[31:0] addr_8129_7;

Selector_2 s8129_7(wires_2032_6[1], addr_2032_6, addr_positional[32519:32516], addr_8129_7);

wire[31:0] addr_8130_7;

Selector_2 s8130_7(wires_2032_6[2], addr_2032_6, addr_positional[32523:32520], addr_8130_7);

wire[31:0] addr_8131_7;

Selector_2 s8131_7(wires_2032_6[3], addr_2032_6, addr_positional[32527:32524], addr_8131_7);

wire[31:0] addr_8132_7;

Selector_2 s8132_7(wires_2033_6[0], addr_2033_6, addr_positional[32531:32528], addr_8132_7);

wire[31:0] addr_8133_7;

Selector_2 s8133_7(wires_2033_6[1], addr_2033_6, addr_positional[32535:32532], addr_8133_7);

wire[31:0] addr_8134_7;

Selector_2 s8134_7(wires_2033_6[2], addr_2033_6, addr_positional[32539:32536], addr_8134_7);

wire[31:0] addr_8135_7;

Selector_2 s8135_7(wires_2033_6[3], addr_2033_6, addr_positional[32543:32540], addr_8135_7);

wire[31:0] addr_8136_7;

Selector_2 s8136_7(wires_2034_6[0], addr_2034_6, addr_positional[32547:32544], addr_8136_7);

wire[31:0] addr_8137_7;

Selector_2 s8137_7(wires_2034_6[1], addr_2034_6, addr_positional[32551:32548], addr_8137_7);

wire[31:0] addr_8138_7;

Selector_2 s8138_7(wires_2034_6[2], addr_2034_6, addr_positional[32555:32552], addr_8138_7);

wire[31:0] addr_8139_7;

Selector_2 s8139_7(wires_2034_6[3], addr_2034_6, addr_positional[32559:32556], addr_8139_7);

wire[31:0] addr_8140_7;

Selector_2 s8140_7(wires_2035_6[0], addr_2035_6, addr_positional[32563:32560], addr_8140_7);

wire[31:0] addr_8141_7;

Selector_2 s8141_7(wires_2035_6[1], addr_2035_6, addr_positional[32567:32564], addr_8141_7);

wire[31:0] addr_8142_7;

Selector_2 s8142_7(wires_2035_6[2], addr_2035_6, addr_positional[32571:32568], addr_8142_7);

wire[31:0] addr_8143_7;

Selector_2 s8143_7(wires_2035_6[3], addr_2035_6, addr_positional[32575:32572], addr_8143_7);

wire[31:0] addr_8144_7;

Selector_2 s8144_7(wires_2036_6[0], addr_2036_6, addr_positional[32579:32576], addr_8144_7);

wire[31:0] addr_8145_7;

Selector_2 s8145_7(wires_2036_6[1], addr_2036_6, addr_positional[32583:32580], addr_8145_7);

wire[31:0] addr_8146_7;

Selector_2 s8146_7(wires_2036_6[2], addr_2036_6, addr_positional[32587:32584], addr_8146_7);

wire[31:0] addr_8147_7;

Selector_2 s8147_7(wires_2036_6[3], addr_2036_6, addr_positional[32591:32588], addr_8147_7);

wire[31:0] addr_8148_7;

Selector_2 s8148_7(wires_2037_6[0], addr_2037_6, addr_positional[32595:32592], addr_8148_7);

wire[31:0] addr_8149_7;

Selector_2 s8149_7(wires_2037_6[1], addr_2037_6, addr_positional[32599:32596], addr_8149_7);

wire[31:0] addr_8150_7;

Selector_2 s8150_7(wires_2037_6[2], addr_2037_6, addr_positional[32603:32600], addr_8150_7);

wire[31:0] addr_8151_7;

Selector_2 s8151_7(wires_2037_6[3], addr_2037_6, addr_positional[32607:32604], addr_8151_7);

wire[31:0] addr_8152_7;

Selector_2 s8152_7(wires_2038_6[0], addr_2038_6, addr_positional[32611:32608], addr_8152_7);

wire[31:0] addr_8153_7;

Selector_2 s8153_7(wires_2038_6[1], addr_2038_6, addr_positional[32615:32612], addr_8153_7);

wire[31:0] addr_8154_7;

Selector_2 s8154_7(wires_2038_6[2], addr_2038_6, addr_positional[32619:32616], addr_8154_7);

wire[31:0] addr_8155_7;

Selector_2 s8155_7(wires_2038_6[3], addr_2038_6, addr_positional[32623:32620], addr_8155_7);

wire[31:0] addr_8156_7;

Selector_2 s8156_7(wires_2039_6[0], addr_2039_6, addr_positional[32627:32624], addr_8156_7);

wire[31:0] addr_8157_7;

Selector_2 s8157_7(wires_2039_6[1], addr_2039_6, addr_positional[32631:32628], addr_8157_7);

wire[31:0] addr_8158_7;

Selector_2 s8158_7(wires_2039_6[2], addr_2039_6, addr_positional[32635:32632], addr_8158_7);

wire[31:0] addr_8159_7;

Selector_2 s8159_7(wires_2039_6[3], addr_2039_6, addr_positional[32639:32636], addr_8159_7);

wire[31:0] addr_8160_7;

Selector_2 s8160_7(wires_2040_6[0], addr_2040_6, addr_positional[32643:32640], addr_8160_7);

wire[31:0] addr_8161_7;

Selector_2 s8161_7(wires_2040_6[1], addr_2040_6, addr_positional[32647:32644], addr_8161_7);

wire[31:0] addr_8162_7;

Selector_2 s8162_7(wires_2040_6[2], addr_2040_6, addr_positional[32651:32648], addr_8162_7);

wire[31:0] addr_8163_7;

Selector_2 s8163_7(wires_2040_6[3], addr_2040_6, addr_positional[32655:32652], addr_8163_7);

wire[31:0] addr_8164_7;

Selector_2 s8164_7(wires_2041_6[0], addr_2041_6, addr_positional[32659:32656], addr_8164_7);

wire[31:0] addr_8165_7;

Selector_2 s8165_7(wires_2041_6[1], addr_2041_6, addr_positional[32663:32660], addr_8165_7);

wire[31:0] addr_8166_7;

Selector_2 s8166_7(wires_2041_6[2], addr_2041_6, addr_positional[32667:32664], addr_8166_7);

wire[31:0] addr_8167_7;

Selector_2 s8167_7(wires_2041_6[3], addr_2041_6, addr_positional[32671:32668], addr_8167_7);

wire[31:0] addr_8168_7;

Selector_2 s8168_7(wires_2042_6[0], addr_2042_6, addr_positional[32675:32672], addr_8168_7);

wire[31:0] addr_8169_7;

Selector_2 s8169_7(wires_2042_6[1], addr_2042_6, addr_positional[32679:32676], addr_8169_7);

wire[31:0] addr_8170_7;

Selector_2 s8170_7(wires_2042_6[2], addr_2042_6, addr_positional[32683:32680], addr_8170_7);

wire[31:0] addr_8171_7;

Selector_2 s8171_7(wires_2042_6[3], addr_2042_6, addr_positional[32687:32684], addr_8171_7);

wire[31:0] addr_8172_7;

Selector_2 s8172_7(wires_2043_6[0], addr_2043_6, addr_positional[32691:32688], addr_8172_7);

wire[31:0] addr_8173_7;

Selector_2 s8173_7(wires_2043_6[1], addr_2043_6, addr_positional[32695:32692], addr_8173_7);

wire[31:0] addr_8174_7;

Selector_2 s8174_7(wires_2043_6[2], addr_2043_6, addr_positional[32699:32696], addr_8174_7);

wire[31:0] addr_8175_7;

Selector_2 s8175_7(wires_2043_6[3], addr_2043_6, addr_positional[32703:32700], addr_8175_7);

wire[31:0] addr_8176_7;

Selector_2 s8176_7(wires_2044_6[0], addr_2044_6, addr_positional[32707:32704], addr_8176_7);

wire[31:0] addr_8177_7;

Selector_2 s8177_7(wires_2044_6[1], addr_2044_6, addr_positional[32711:32708], addr_8177_7);

wire[31:0] addr_8178_7;

Selector_2 s8178_7(wires_2044_6[2], addr_2044_6, addr_positional[32715:32712], addr_8178_7);

wire[31:0] addr_8179_7;

Selector_2 s8179_7(wires_2044_6[3], addr_2044_6, addr_positional[32719:32716], addr_8179_7);

wire[31:0] addr_8180_7;

Selector_2 s8180_7(wires_2045_6[0], addr_2045_6, addr_positional[32723:32720], addr_8180_7);

wire[31:0] addr_8181_7;

Selector_2 s8181_7(wires_2045_6[1], addr_2045_6, addr_positional[32727:32724], addr_8181_7);

wire[31:0] addr_8182_7;

Selector_2 s8182_7(wires_2045_6[2], addr_2045_6, addr_positional[32731:32728], addr_8182_7);

wire[31:0] addr_8183_7;

Selector_2 s8183_7(wires_2045_6[3], addr_2045_6, addr_positional[32735:32732], addr_8183_7);

wire[31:0] addr_8184_7;

Selector_2 s8184_7(wires_2046_6[0], addr_2046_6, addr_positional[32739:32736], addr_8184_7);

wire[31:0] addr_8185_7;

Selector_2 s8185_7(wires_2046_6[1], addr_2046_6, addr_positional[32743:32740], addr_8185_7);

wire[31:0] addr_8186_7;

Selector_2 s8186_7(wires_2046_6[2], addr_2046_6, addr_positional[32747:32744], addr_8186_7);

wire[31:0] addr_8187_7;

Selector_2 s8187_7(wires_2046_6[3], addr_2046_6, addr_positional[32751:32748], addr_8187_7);

wire[31:0] addr_8188_7;

Selector_2 s8188_7(wires_2047_6[0], addr_2047_6, addr_positional[32755:32752], addr_8188_7);

wire[31:0] addr_8189_7;

Selector_2 s8189_7(wires_2047_6[1], addr_2047_6, addr_positional[32759:32756], addr_8189_7);

wire[31:0] addr_8190_7;

Selector_2 s8190_7(wires_2047_6[2], addr_2047_6, addr_positional[32763:32760], addr_8190_7);

wire[31:0] addr_8191_7;

Selector_2 s8191_7(wires_2047_6[3], addr_2047_6, addr_positional[32767:32764], addr_8191_7);

wire[31:0] addr_8192_7;

Selector_2 s8192_7(wires_2048_6[0], addr_2048_6, addr_positional[32771:32768], addr_8192_7);

wire[31:0] addr_8193_7;

Selector_2 s8193_7(wires_2048_6[1], addr_2048_6, addr_positional[32775:32772], addr_8193_7);

wire[31:0] addr_8194_7;

Selector_2 s8194_7(wires_2048_6[2], addr_2048_6, addr_positional[32779:32776], addr_8194_7);

wire[31:0] addr_8195_7;

Selector_2 s8195_7(wires_2048_6[3], addr_2048_6, addr_positional[32783:32780], addr_8195_7);

wire[31:0] addr_8196_7;

Selector_2 s8196_7(wires_2049_6[0], addr_2049_6, addr_positional[32787:32784], addr_8196_7);

wire[31:0] addr_8197_7;

Selector_2 s8197_7(wires_2049_6[1], addr_2049_6, addr_positional[32791:32788], addr_8197_7);

wire[31:0] addr_8198_7;

Selector_2 s8198_7(wires_2049_6[2], addr_2049_6, addr_positional[32795:32792], addr_8198_7);

wire[31:0] addr_8199_7;

Selector_2 s8199_7(wires_2049_6[3], addr_2049_6, addr_positional[32799:32796], addr_8199_7);

wire[31:0] addr_8200_7;

Selector_2 s8200_7(wires_2050_6[0], addr_2050_6, addr_positional[32803:32800], addr_8200_7);

wire[31:0] addr_8201_7;

Selector_2 s8201_7(wires_2050_6[1], addr_2050_6, addr_positional[32807:32804], addr_8201_7);

wire[31:0] addr_8202_7;

Selector_2 s8202_7(wires_2050_6[2], addr_2050_6, addr_positional[32811:32808], addr_8202_7);

wire[31:0] addr_8203_7;

Selector_2 s8203_7(wires_2050_6[3], addr_2050_6, addr_positional[32815:32812], addr_8203_7);

wire[31:0] addr_8204_7;

Selector_2 s8204_7(wires_2051_6[0], addr_2051_6, addr_positional[32819:32816], addr_8204_7);

wire[31:0] addr_8205_7;

Selector_2 s8205_7(wires_2051_6[1], addr_2051_6, addr_positional[32823:32820], addr_8205_7);

wire[31:0] addr_8206_7;

Selector_2 s8206_7(wires_2051_6[2], addr_2051_6, addr_positional[32827:32824], addr_8206_7);

wire[31:0] addr_8207_7;

Selector_2 s8207_7(wires_2051_6[3], addr_2051_6, addr_positional[32831:32828], addr_8207_7);

wire[31:0] addr_8208_7;

Selector_2 s8208_7(wires_2052_6[0], addr_2052_6, addr_positional[32835:32832], addr_8208_7);

wire[31:0] addr_8209_7;

Selector_2 s8209_7(wires_2052_6[1], addr_2052_6, addr_positional[32839:32836], addr_8209_7);

wire[31:0] addr_8210_7;

Selector_2 s8210_7(wires_2052_6[2], addr_2052_6, addr_positional[32843:32840], addr_8210_7);

wire[31:0] addr_8211_7;

Selector_2 s8211_7(wires_2052_6[3], addr_2052_6, addr_positional[32847:32844], addr_8211_7);

wire[31:0] addr_8212_7;

Selector_2 s8212_7(wires_2053_6[0], addr_2053_6, addr_positional[32851:32848], addr_8212_7);

wire[31:0] addr_8213_7;

Selector_2 s8213_7(wires_2053_6[1], addr_2053_6, addr_positional[32855:32852], addr_8213_7);

wire[31:0] addr_8214_7;

Selector_2 s8214_7(wires_2053_6[2], addr_2053_6, addr_positional[32859:32856], addr_8214_7);

wire[31:0] addr_8215_7;

Selector_2 s8215_7(wires_2053_6[3], addr_2053_6, addr_positional[32863:32860], addr_8215_7);

wire[31:0] addr_8216_7;

Selector_2 s8216_7(wires_2054_6[0], addr_2054_6, addr_positional[32867:32864], addr_8216_7);

wire[31:0] addr_8217_7;

Selector_2 s8217_7(wires_2054_6[1], addr_2054_6, addr_positional[32871:32868], addr_8217_7);

wire[31:0] addr_8218_7;

Selector_2 s8218_7(wires_2054_6[2], addr_2054_6, addr_positional[32875:32872], addr_8218_7);

wire[31:0] addr_8219_7;

Selector_2 s8219_7(wires_2054_6[3], addr_2054_6, addr_positional[32879:32876], addr_8219_7);

wire[31:0] addr_8220_7;

Selector_2 s8220_7(wires_2055_6[0], addr_2055_6, addr_positional[32883:32880], addr_8220_7);

wire[31:0] addr_8221_7;

Selector_2 s8221_7(wires_2055_6[1], addr_2055_6, addr_positional[32887:32884], addr_8221_7);

wire[31:0] addr_8222_7;

Selector_2 s8222_7(wires_2055_6[2], addr_2055_6, addr_positional[32891:32888], addr_8222_7);

wire[31:0] addr_8223_7;

Selector_2 s8223_7(wires_2055_6[3], addr_2055_6, addr_positional[32895:32892], addr_8223_7);

wire[31:0] addr_8224_7;

Selector_2 s8224_7(wires_2056_6[0], addr_2056_6, addr_positional[32899:32896], addr_8224_7);

wire[31:0] addr_8225_7;

Selector_2 s8225_7(wires_2056_6[1], addr_2056_6, addr_positional[32903:32900], addr_8225_7);

wire[31:0] addr_8226_7;

Selector_2 s8226_7(wires_2056_6[2], addr_2056_6, addr_positional[32907:32904], addr_8226_7);

wire[31:0] addr_8227_7;

Selector_2 s8227_7(wires_2056_6[3], addr_2056_6, addr_positional[32911:32908], addr_8227_7);

wire[31:0] addr_8228_7;

Selector_2 s8228_7(wires_2057_6[0], addr_2057_6, addr_positional[32915:32912], addr_8228_7);

wire[31:0] addr_8229_7;

Selector_2 s8229_7(wires_2057_6[1], addr_2057_6, addr_positional[32919:32916], addr_8229_7);

wire[31:0] addr_8230_7;

Selector_2 s8230_7(wires_2057_6[2], addr_2057_6, addr_positional[32923:32920], addr_8230_7);

wire[31:0] addr_8231_7;

Selector_2 s8231_7(wires_2057_6[3], addr_2057_6, addr_positional[32927:32924], addr_8231_7);

wire[31:0] addr_8232_7;

Selector_2 s8232_7(wires_2058_6[0], addr_2058_6, addr_positional[32931:32928], addr_8232_7);

wire[31:0] addr_8233_7;

Selector_2 s8233_7(wires_2058_6[1], addr_2058_6, addr_positional[32935:32932], addr_8233_7);

wire[31:0] addr_8234_7;

Selector_2 s8234_7(wires_2058_6[2], addr_2058_6, addr_positional[32939:32936], addr_8234_7);

wire[31:0] addr_8235_7;

Selector_2 s8235_7(wires_2058_6[3], addr_2058_6, addr_positional[32943:32940], addr_8235_7);

wire[31:0] addr_8236_7;

Selector_2 s8236_7(wires_2059_6[0], addr_2059_6, addr_positional[32947:32944], addr_8236_7);

wire[31:0] addr_8237_7;

Selector_2 s8237_7(wires_2059_6[1], addr_2059_6, addr_positional[32951:32948], addr_8237_7);

wire[31:0] addr_8238_7;

Selector_2 s8238_7(wires_2059_6[2], addr_2059_6, addr_positional[32955:32952], addr_8238_7);

wire[31:0] addr_8239_7;

Selector_2 s8239_7(wires_2059_6[3], addr_2059_6, addr_positional[32959:32956], addr_8239_7);

wire[31:0] addr_8240_7;

Selector_2 s8240_7(wires_2060_6[0], addr_2060_6, addr_positional[32963:32960], addr_8240_7);

wire[31:0] addr_8241_7;

Selector_2 s8241_7(wires_2060_6[1], addr_2060_6, addr_positional[32967:32964], addr_8241_7);

wire[31:0] addr_8242_7;

Selector_2 s8242_7(wires_2060_6[2], addr_2060_6, addr_positional[32971:32968], addr_8242_7);

wire[31:0] addr_8243_7;

Selector_2 s8243_7(wires_2060_6[3], addr_2060_6, addr_positional[32975:32972], addr_8243_7);

wire[31:0] addr_8244_7;

Selector_2 s8244_7(wires_2061_6[0], addr_2061_6, addr_positional[32979:32976], addr_8244_7);

wire[31:0] addr_8245_7;

Selector_2 s8245_7(wires_2061_6[1], addr_2061_6, addr_positional[32983:32980], addr_8245_7);

wire[31:0] addr_8246_7;

Selector_2 s8246_7(wires_2061_6[2], addr_2061_6, addr_positional[32987:32984], addr_8246_7);

wire[31:0] addr_8247_7;

Selector_2 s8247_7(wires_2061_6[3], addr_2061_6, addr_positional[32991:32988], addr_8247_7);

wire[31:0] addr_8248_7;

Selector_2 s8248_7(wires_2062_6[0], addr_2062_6, addr_positional[32995:32992], addr_8248_7);

wire[31:0] addr_8249_7;

Selector_2 s8249_7(wires_2062_6[1], addr_2062_6, addr_positional[32999:32996], addr_8249_7);

wire[31:0] addr_8250_7;

Selector_2 s8250_7(wires_2062_6[2], addr_2062_6, addr_positional[33003:33000], addr_8250_7);

wire[31:0] addr_8251_7;

Selector_2 s8251_7(wires_2062_6[3], addr_2062_6, addr_positional[33007:33004], addr_8251_7);

wire[31:0] addr_8252_7;

Selector_2 s8252_7(wires_2063_6[0], addr_2063_6, addr_positional[33011:33008], addr_8252_7);

wire[31:0] addr_8253_7;

Selector_2 s8253_7(wires_2063_6[1], addr_2063_6, addr_positional[33015:33012], addr_8253_7);

wire[31:0] addr_8254_7;

Selector_2 s8254_7(wires_2063_6[2], addr_2063_6, addr_positional[33019:33016], addr_8254_7);

wire[31:0] addr_8255_7;

Selector_2 s8255_7(wires_2063_6[3], addr_2063_6, addr_positional[33023:33020], addr_8255_7);

wire[31:0] addr_8256_7;

Selector_2 s8256_7(wires_2064_6[0], addr_2064_6, addr_positional[33027:33024], addr_8256_7);

wire[31:0] addr_8257_7;

Selector_2 s8257_7(wires_2064_6[1], addr_2064_6, addr_positional[33031:33028], addr_8257_7);

wire[31:0] addr_8258_7;

Selector_2 s8258_7(wires_2064_6[2], addr_2064_6, addr_positional[33035:33032], addr_8258_7);

wire[31:0] addr_8259_7;

Selector_2 s8259_7(wires_2064_6[3], addr_2064_6, addr_positional[33039:33036], addr_8259_7);

wire[31:0] addr_8260_7;

Selector_2 s8260_7(wires_2065_6[0], addr_2065_6, addr_positional[33043:33040], addr_8260_7);

wire[31:0] addr_8261_7;

Selector_2 s8261_7(wires_2065_6[1], addr_2065_6, addr_positional[33047:33044], addr_8261_7);

wire[31:0] addr_8262_7;

Selector_2 s8262_7(wires_2065_6[2], addr_2065_6, addr_positional[33051:33048], addr_8262_7);

wire[31:0] addr_8263_7;

Selector_2 s8263_7(wires_2065_6[3], addr_2065_6, addr_positional[33055:33052], addr_8263_7);

wire[31:0] addr_8264_7;

Selector_2 s8264_7(wires_2066_6[0], addr_2066_6, addr_positional[33059:33056], addr_8264_7);

wire[31:0] addr_8265_7;

Selector_2 s8265_7(wires_2066_6[1], addr_2066_6, addr_positional[33063:33060], addr_8265_7);

wire[31:0] addr_8266_7;

Selector_2 s8266_7(wires_2066_6[2], addr_2066_6, addr_positional[33067:33064], addr_8266_7);

wire[31:0] addr_8267_7;

Selector_2 s8267_7(wires_2066_6[3], addr_2066_6, addr_positional[33071:33068], addr_8267_7);

wire[31:0] addr_8268_7;

Selector_2 s8268_7(wires_2067_6[0], addr_2067_6, addr_positional[33075:33072], addr_8268_7);

wire[31:0] addr_8269_7;

Selector_2 s8269_7(wires_2067_6[1], addr_2067_6, addr_positional[33079:33076], addr_8269_7);

wire[31:0] addr_8270_7;

Selector_2 s8270_7(wires_2067_6[2], addr_2067_6, addr_positional[33083:33080], addr_8270_7);

wire[31:0] addr_8271_7;

Selector_2 s8271_7(wires_2067_6[3], addr_2067_6, addr_positional[33087:33084], addr_8271_7);

wire[31:0] addr_8272_7;

Selector_2 s8272_7(wires_2068_6[0], addr_2068_6, addr_positional[33091:33088], addr_8272_7);

wire[31:0] addr_8273_7;

Selector_2 s8273_7(wires_2068_6[1], addr_2068_6, addr_positional[33095:33092], addr_8273_7);

wire[31:0] addr_8274_7;

Selector_2 s8274_7(wires_2068_6[2], addr_2068_6, addr_positional[33099:33096], addr_8274_7);

wire[31:0] addr_8275_7;

Selector_2 s8275_7(wires_2068_6[3], addr_2068_6, addr_positional[33103:33100], addr_8275_7);

wire[31:0] addr_8276_7;

Selector_2 s8276_7(wires_2069_6[0], addr_2069_6, addr_positional[33107:33104], addr_8276_7);

wire[31:0] addr_8277_7;

Selector_2 s8277_7(wires_2069_6[1], addr_2069_6, addr_positional[33111:33108], addr_8277_7);

wire[31:0] addr_8278_7;

Selector_2 s8278_7(wires_2069_6[2], addr_2069_6, addr_positional[33115:33112], addr_8278_7);

wire[31:0] addr_8279_7;

Selector_2 s8279_7(wires_2069_6[3], addr_2069_6, addr_positional[33119:33116], addr_8279_7);

wire[31:0] addr_8280_7;

Selector_2 s8280_7(wires_2070_6[0], addr_2070_6, addr_positional[33123:33120], addr_8280_7);

wire[31:0] addr_8281_7;

Selector_2 s8281_7(wires_2070_6[1], addr_2070_6, addr_positional[33127:33124], addr_8281_7);

wire[31:0] addr_8282_7;

Selector_2 s8282_7(wires_2070_6[2], addr_2070_6, addr_positional[33131:33128], addr_8282_7);

wire[31:0] addr_8283_7;

Selector_2 s8283_7(wires_2070_6[3], addr_2070_6, addr_positional[33135:33132], addr_8283_7);

wire[31:0] addr_8284_7;

Selector_2 s8284_7(wires_2071_6[0], addr_2071_6, addr_positional[33139:33136], addr_8284_7);

wire[31:0] addr_8285_7;

Selector_2 s8285_7(wires_2071_6[1], addr_2071_6, addr_positional[33143:33140], addr_8285_7);

wire[31:0] addr_8286_7;

Selector_2 s8286_7(wires_2071_6[2], addr_2071_6, addr_positional[33147:33144], addr_8286_7);

wire[31:0] addr_8287_7;

Selector_2 s8287_7(wires_2071_6[3], addr_2071_6, addr_positional[33151:33148], addr_8287_7);

wire[31:0] addr_8288_7;

Selector_2 s8288_7(wires_2072_6[0], addr_2072_6, addr_positional[33155:33152], addr_8288_7);

wire[31:0] addr_8289_7;

Selector_2 s8289_7(wires_2072_6[1], addr_2072_6, addr_positional[33159:33156], addr_8289_7);

wire[31:0] addr_8290_7;

Selector_2 s8290_7(wires_2072_6[2], addr_2072_6, addr_positional[33163:33160], addr_8290_7);

wire[31:0] addr_8291_7;

Selector_2 s8291_7(wires_2072_6[3], addr_2072_6, addr_positional[33167:33164], addr_8291_7);

wire[31:0] addr_8292_7;

Selector_2 s8292_7(wires_2073_6[0], addr_2073_6, addr_positional[33171:33168], addr_8292_7);

wire[31:0] addr_8293_7;

Selector_2 s8293_7(wires_2073_6[1], addr_2073_6, addr_positional[33175:33172], addr_8293_7);

wire[31:0] addr_8294_7;

Selector_2 s8294_7(wires_2073_6[2], addr_2073_6, addr_positional[33179:33176], addr_8294_7);

wire[31:0] addr_8295_7;

Selector_2 s8295_7(wires_2073_6[3], addr_2073_6, addr_positional[33183:33180], addr_8295_7);

wire[31:0] addr_8296_7;

Selector_2 s8296_7(wires_2074_6[0], addr_2074_6, addr_positional[33187:33184], addr_8296_7);

wire[31:0] addr_8297_7;

Selector_2 s8297_7(wires_2074_6[1], addr_2074_6, addr_positional[33191:33188], addr_8297_7);

wire[31:0] addr_8298_7;

Selector_2 s8298_7(wires_2074_6[2], addr_2074_6, addr_positional[33195:33192], addr_8298_7);

wire[31:0] addr_8299_7;

Selector_2 s8299_7(wires_2074_6[3], addr_2074_6, addr_positional[33199:33196], addr_8299_7);

wire[31:0] addr_8300_7;

Selector_2 s8300_7(wires_2075_6[0], addr_2075_6, addr_positional[33203:33200], addr_8300_7);

wire[31:0] addr_8301_7;

Selector_2 s8301_7(wires_2075_6[1], addr_2075_6, addr_positional[33207:33204], addr_8301_7);

wire[31:0] addr_8302_7;

Selector_2 s8302_7(wires_2075_6[2], addr_2075_6, addr_positional[33211:33208], addr_8302_7);

wire[31:0] addr_8303_7;

Selector_2 s8303_7(wires_2075_6[3], addr_2075_6, addr_positional[33215:33212], addr_8303_7);

wire[31:0] addr_8304_7;

Selector_2 s8304_7(wires_2076_6[0], addr_2076_6, addr_positional[33219:33216], addr_8304_7);

wire[31:0] addr_8305_7;

Selector_2 s8305_7(wires_2076_6[1], addr_2076_6, addr_positional[33223:33220], addr_8305_7);

wire[31:0] addr_8306_7;

Selector_2 s8306_7(wires_2076_6[2], addr_2076_6, addr_positional[33227:33224], addr_8306_7);

wire[31:0] addr_8307_7;

Selector_2 s8307_7(wires_2076_6[3], addr_2076_6, addr_positional[33231:33228], addr_8307_7);

wire[31:0] addr_8308_7;

Selector_2 s8308_7(wires_2077_6[0], addr_2077_6, addr_positional[33235:33232], addr_8308_7);

wire[31:0] addr_8309_7;

Selector_2 s8309_7(wires_2077_6[1], addr_2077_6, addr_positional[33239:33236], addr_8309_7);

wire[31:0] addr_8310_7;

Selector_2 s8310_7(wires_2077_6[2], addr_2077_6, addr_positional[33243:33240], addr_8310_7);

wire[31:0] addr_8311_7;

Selector_2 s8311_7(wires_2077_6[3], addr_2077_6, addr_positional[33247:33244], addr_8311_7);

wire[31:0] addr_8312_7;

Selector_2 s8312_7(wires_2078_6[0], addr_2078_6, addr_positional[33251:33248], addr_8312_7);

wire[31:0] addr_8313_7;

Selector_2 s8313_7(wires_2078_6[1], addr_2078_6, addr_positional[33255:33252], addr_8313_7);

wire[31:0] addr_8314_7;

Selector_2 s8314_7(wires_2078_6[2], addr_2078_6, addr_positional[33259:33256], addr_8314_7);

wire[31:0] addr_8315_7;

Selector_2 s8315_7(wires_2078_6[3], addr_2078_6, addr_positional[33263:33260], addr_8315_7);

wire[31:0] addr_8316_7;

Selector_2 s8316_7(wires_2079_6[0], addr_2079_6, addr_positional[33267:33264], addr_8316_7);

wire[31:0] addr_8317_7;

Selector_2 s8317_7(wires_2079_6[1], addr_2079_6, addr_positional[33271:33268], addr_8317_7);

wire[31:0] addr_8318_7;

Selector_2 s8318_7(wires_2079_6[2], addr_2079_6, addr_positional[33275:33272], addr_8318_7);

wire[31:0] addr_8319_7;

Selector_2 s8319_7(wires_2079_6[3], addr_2079_6, addr_positional[33279:33276], addr_8319_7);

wire[31:0] addr_8320_7;

Selector_2 s8320_7(wires_2080_6[0], addr_2080_6, addr_positional[33283:33280], addr_8320_7);

wire[31:0] addr_8321_7;

Selector_2 s8321_7(wires_2080_6[1], addr_2080_6, addr_positional[33287:33284], addr_8321_7);

wire[31:0] addr_8322_7;

Selector_2 s8322_7(wires_2080_6[2], addr_2080_6, addr_positional[33291:33288], addr_8322_7);

wire[31:0] addr_8323_7;

Selector_2 s8323_7(wires_2080_6[3], addr_2080_6, addr_positional[33295:33292], addr_8323_7);

wire[31:0] addr_8324_7;

Selector_2 s8324_7(wires_2081_6[0], addr_2081_6, addr_positional[33299:33296], addr_8324_7);

wire[31:0] addr_8325_7;

Selector_2 s8325_7(wires_2081_6[1], addr_2081_6, addr_positional[33303:33300], addr_8325_7);

wire[31:0] addr_8326_7;

Selector_2 s8326_7(wires_2081_6[2], addr_2081_6, addr_positional[33307:33304], addr_8326_7);

wire[31:0] addr_8327_7;

Selector_2 s8327_7(wires_2081_6[3], addr_2081_6, addr_positional[33311:33308], addr_8327_7);

wire[31:0] addr_8328_7;

Selector_2 s8328_7(wires_2082_6[0], addr_2082_6, addr_positional[33315:33312], addr_8328_7);

wire[31:0] addr_8329_7;

Selector_2 s8329_7(wires_2082_6[1], addr_2082_6, addr_positional[33319:33316], addr_8329_7);

wire[31:0] addr_8330_7;

Selector_2 s8330_7(wires_2082_6[2], addr_2082_6, addr_positional[33323:33320], addr_8330_7);

wire[31:0] addr_8331_7;

Selector_2 s8331_7(wires_2082_6[3], addr_2082_6, addr_positional[33327:33324], addr_8331_7);

wire[31:0] addr_8332_7;

Selector_2 s8332_7(wires_2083_6[0], addr_2083_6, addr_positional[33331:33328], addr_8332_7);

wire[31:0] addr_8333_7;

Selector_2 s8333_7(wires_2083_6[1], addr_2083_6, addr_positional[33335:33332], addr_8333_7);

wire[31:0] addr_8334_7;

Selector_2 s8334_7(wires_2083_6[2], addr_2083_6, addr_positional[33339:33336], addr_8334_7);

wire[31:0] addr_8335_7;

Selector_2 s8335_7(wires_2083_6[3], addr_2083_6, addr_positional[33343:33340], addr_8335_7);

wire[31:0] addr_8336_7;

Selector_2 s8336_7(wires_2084_6[0], addr_2084_6, addr_positional[33347:33344], addr_8336_7);

wire[31:0] addr_8337_7;

Selector_2 s8337_7(wires_2084_6[1], addr_2084_6, addr_positional[33351:33348], addr_8337_7);

wire[31:0] addr_8338_7;

Selector_2 s8338_7(wires_2084_6[2], addr_2084_6, addr_positional[33355:33352], addr_8338_7);

wire[31:0] addr_8339_7;

Selector_2 s8339_7(wires_2084_6[3], addr_2084_6, addr_positional[33359:33356], addr_8339_7);

wire[31:0] addr_8340_7;

Selector_2 s8340_7(wires_2085_6[0], addr_2085_6, addr_positional[33363:33360], addr_8340_7);

wire[31:0] addr_8341_7;

Selector_2 s8341_7(wires_2085_6[1], addr_2085_6, addr_positional[33367:33364], addr_8341_7);

wire[31:0] addr_8342_7;

Selector_2 s8342_7(wires_2085_6[2], addr_2085_6, addr_positional[33371:33368], addr_8342_7);

wire[31:0] addr_8343_7;

Selector_2 s8343_7(wires_2085_6[3], addr_2085_6, addr_positional[33375:33372], addr_8343_7);

wire[31:0] addr_8344_7;

Selector_2 s8344_7(wires_2086_6[0], addr_2086_6, addr_positional[33379:33376], addr_8344_7);

wire[31:0] addr_8345_7;

Selector_2 s8345_7(wires_2086_6[1], addr_2086_6, addr_positional[33383:33380], addr_8345_7);

wire[31:0] addr_8346_7;

Selector_2 s8346_7(wires_2086_6[2], addr_2086_6, addr_positional[33387:33384], addr_8346_7);

wire[31:0] addr_8347_7;

Selector_2 s8347_7(wires_2086_6[3], addr_2086_6, addr_positional[33391:33388], addr_8347_7);

wire[31:0] addr_8348_7;

Selector_2 s8348_7(wires_2087_6[0], addr_2087_6, addr_positional[33395:33392], addr_8348_7);

wire[31:0] addr_8349_7;

Selector_2 s8349_7(wires_2087_6[1], addr_2087_6, addr_positional[33399:33396], addr_8349_7);

wire[31:0] addr_8350_7;

Selector_2 s8350_7(wires_2087_6[2], addr_2087_6, addr_positional[33403:33400], addr_8350_7);

wire[31:0] addr_8351_7;

Selector_2 s8351_7(wires_2087_6[3], addr_2087_6, addr_positional[33407:33404], addr_8351_7);

wire[31:0] addr_8352_7;

Selector_2 s8352_7(wires_2088_6[0], addr_2088_6, addr_positional[33411:33408], addr_8352_7);

wire[31:0] addr_8353_7;

Selector_2 s8353_7(wires_2088_6[1], addr_2088_6, addr_positional[33415:33412], addr_8353_7);

wire[31:0] addr_8354_7;

Selector_2 s8354_7(wires_2088_6[2], addr_2088_6, addr_positional[33419:33416], addr_8354_7);

wire[31:0] addr_8355_7;

Selector_2 s8355_7(wires_2088_6[3], addr_2088_6, addr_positional[33423:33420], addr_8355_7);

wire[31:0] addr_8356_7;

Selector_2 s8356_7(wires_2089_6[0], addr_2089_6, addr_positional[33427:33424], addr_8356_7);

wire[31:0] addr_8357_7;

Selector_2 s8357_7(wires_2089_6[1], addr_2089_6, addr_positional[33431:33428], addr_8357_7);

wire[31:0] addr_8358_7;

Selector_2 s8358_7(wires_2089_6[2], addr_2089_6, addr_positional[33435:33432], addr_8358_7);

wire[31:0] addr_8359_7;

Selector_2 s8359_7(wires_2089_6[3], addr_2089_6, addr_positional[33439:33436], addr_8359_7);

wire[31:0] addr_8360_7;

Selector_2 s8360_7(wires_2090_6[0], addr_2090_6, addr_positional[33443:33440], addr_8360_7);

wire[31:0] addr_8361_7;

Selector_2 s8361_7(wires_2090_6[1], addr_2090_6, addr_positional[33447:33444], addr_8361_7);

wire[31:0] addr_8362_7;

Selector_2 s8362_7(wires_2090_6[2], addr_2090_6, addr_positional[33451:33448], addr_8362_7);

wire[31:0] addr_8363_7;

Selector_2 s8363_7(wires_2090_6[3], addr_2090_6, addr_positional[33455:33452], addr_8363_7);

wire[31:0] addr_8364_7;

Selector_2 s8364_7(wires_2091_6[0], addr_2091_6, addr_positional[33459:33456], addr_8364_7);

wire[31:0] addr_8365_7;

Selector_2 s8365_7(wires_2091_6[1], addr_2091_6, addr_positional[33463:33460], addr_8365_7);

wire[31:0] addr_8366_7;

Selector_2 s8366_7(wires_2091_6[2], addr_2091_6, addr_positional[33467:33464], addr_8366_7);

wire[31:0] addr_8367_7;

Selector_2 s8367_7(wires_2091_6[3], addr_2091_6, addr_positional[33471:33468], addr_8367_7);

wire[31:0] addr_8368_7;

Selector_2 s8368_7(wires_2092_6[0], addr_2092_6, addr_positional[33475:33472], addr_8368_7);

wire[31:0] addr_8369_7;

Selector_2 s8369_7(wires_2092_6[1], addr_2092_6, addr_positional[33479:33476], addr_8369_7);

wire[31:0] addr_8370_7;

Selector_2 s8370_7(wires_2092_6[2], addr_2092_6, addr_positional[33483:33480], addr_8370_7);

wire[31:0] addr_8371_7;

Selector_2 s8371_7(wires_2092_6[3], addr_2092_6, addr_positional[33487:33484], addr_8371_7);

wire[31:0] addr_8372_7;

Selector_2 s8372_7(wires_2093_6[0], addr_2093_6, addr_positional[33491:33488], addr_8372_7);

wire[31:0] addr_8373_7;

Selector_2 s8373_7(wires_2093_6[1], addr_2093_6, addr_positional[33495:33492], addr_8373_7);

wire[31:0] addr_8374_7;

Selector_2 s8374_7(wires_2093_6[2], addr_2093_6, addr_positional[33499:33496], addr_8374_7);

wire[31:0] addr_8375_7;

Selector_2 s8375_7(wires_2093_6[3], addr_2093_6, addr_positional[33503:33500], addr_8375_7);

wire[31:0] addr_8376_7;

Selector_2 s8376_7(wires_2094_6[0], addr_2094_6, addr_positional[33507:33504], addr_8376_7);

wire[31:0] addr_8377_7;

Selector_2 s8377_7(wires_2094_6[1], addr_2094_6, addr_positional[33511:33508], addr_8377_7);

wire[31:0] addr_8378_7;

Selector_2 s8378_7(wires_2094_6[2], addr_2094_6, addr_positional[33515:33512], addr_8378_7);

wire[31:0] addr_8379_7;

Selector_2 s8379_7(wires_2094_6[3], addr_2094_6, addr_positional[33519:33516], addr_8379_7);

wire[31:0] addr_8380_7;

Selector_2 s8380_7(wires_2095_6[0], addr_2095_6, addr_positional[33523:33520], addr_8380_7);

wire[31:0] addr_8381_7;

Selector_2 s8381_7(wires_2095_6[1], addr_2095_6, addr_positional[33527:33524], addr_8381_7);

wire[31:0] addr_8382_7;

Selector_2 s8382_7(wires_2095_6[2], addr_2095_6, addr_positional[33531:33528], addr_8382_7);

wire[31:0] addr_8383_7;

Selector_2 s8383_7(wires_2095_6[3], addr_2095_6, addr_positional[33535:33532], addr_8383_7);

wire[31:0] addr_8384_7;

Selector_2 s8384_7(wires_2096_6[0], addr_2096_6, addr_positional[33539:33536], addr_8384_7);

wire[31:0] addr_8385_7;

Selector_2 s8385_7(wires_2096_6[1], addr_2096_6, addr_positional[33543:33540], addr_8385_7);

wire[31:0] addr_8386_7;

Selector_2 s8386_7(wires_2096_6[2], addr_2096_6, addr_positional[33547:33544], addr_8386_7);

wire[31:0] addr_8387_7;

Selector_2 s8387_7(wires_2096_6[3], addr_2096_6, addr_positional[33551:33548], addr_8387_7);

wire[31:0] addr_8388_7;

Selector_2 s8388_7(wires_2097_6[0], addr_2097_6, addr_positional[33555:33552], addr_8388_7);

wire[31:0] addr_8389_7;

Selector_2 s8389_7(wires_2097_6[1], addr_2097_6, addr_positional[33559:33556], addr_8389_7);

wire[31:0] addr_8390_7;

Selector_2 s8390_7(wires_2097_6[2], addr_2097_6, addr_positional[33563:33560], addr_8390_7);

wire[31:0] addr_8391_7;

Selector_2 s8391_7(wires_2097_6[3], addr_2097_6, addr_positional[33567:33564], addr_8391_7);

wire[31:0] addr_8392_7;

Selector_2 s8392_7(wires_2098_6[0], addr_2098_6, addr_positional[33571:33568], addr_8392_7);

wire[31:0] addr_8393_7;

Selector_2 s8393_7(wires_2098_6[1], addr_2098_6, addr_positional[33575:33572], addr_8393_7);

wire[31:0] addr_8394_7;

Selector_2 s8394_7(wires_2098_6[2], addr_2098_6, addr_positional[33579:33576], addr_8394_7);

wire[31:0] addr_8395_7;

Selector_2 s8395_7(wires_2098_6[3], addr_2098_6, addr_positional[33583:33580], addr_8395_7);

wire[31:0] addr_8396_7;

Selector_2 s8396_7(wires_2099_6[0], addr_2099_6, addr_positional[33587:33584], addr_8396_7);

wire[31:0] addr_8397_7;

Selector_2 s8397_7(wires_2099_6[1], addr_2099_6, addr_positional[33591:33588], addr_8397_7);

wire[31:0] addr_8398_7;

Selector_2 s8398_7(wires_2099_6[2], addr_2099_6, addr_positional[33595:33592], addr_8398_7);

wire[31:0] addr_8399_7;

Selector_2 s8399_7(wires_2099_6[3], addr_2099_6, addr_positional[33599:33596], addr_8399_7);

wire[31:0] addr_8400_7;

Selector_2 s8400_7(wires_2100_6[0], addr_2100_6, addr_positional[33603:33600], addr_8400_7);

wire[31:0] addr_8401_7;

Selector_2 s8401_7(wires_2100_6[1], addr_2100_6, addr_positional[33607:33604], addr_8401_7);

wire[31:0] addr_8402_7;

Selector_2 s8402_7(wires_2100_6[2], addr_2100_6, addr_positional[33611:33608], addr_8402_7);

wire[31:0] addr_8403_7;

Selector_2 s8403_7(wires_2100_6[3], addr_2100_6, addr_positional[33615:33612], addr_8403_7);

wire[31:0] addr_8404_7;

Selector_2 s8404_7(wires_2101_6[0], addr_2101_6, addr_positional[33619:33616], addr_8404_7);

wire[31:0] addr_8405_7;

Selector_2 s8405_7(wires_2101_6[1], addr_2101_6, addr_positional[33623:33620], addr_8405_7);

wire[31:0] addr_8406_7;

Selector_2 s8406_7(wires_2101_6[2], addr_2101_6, addr_positional[33627:33624], addr_8406_7);

wire[31:0] addr_8407_7;

Selector_2 s8407_7(wires_2101_6[3], addr_2101_6, addr_positional[33631:33628], addr_8407_7);

wire[31:0] addr_8408_7;

Selector_2 s8408_7(wires_2102_6[0], addr_2102_6, addr_positional[33635:33632], addr_8408_7);

wire[31:0] addr_8409_7;

Selector_2 s8409_7(wires_2102_6[1], addr_2102_6, addr_positional[33639:33636], addr_8409_7);

wire[31:0] addr_8410_7;

Selector_2 s8410_7(wires_2102_6[2], addr_2102_6, addr_positional[33643:33640], addr_8410_7);

wire[31:0] addr_8411_7;

Selector_2 s8411_7(wires_2102_6[3], addr_2102_6, addr_positional[33647:33644], addr_8411_7);

wire[31:0] addr_8412_7;

Selector_2 s8412_7(wires_2103_6[0], addr_2103_6, addr_positional[33651:33648], addr_8412_7);

wire[31:0] addr_8413_7;

Selector_2 s8413_7(wires_2103_6[1], addr_2103_6, addr_positional[33655:33652], addr_8413_7);

wire[31:0] addr_8414_7;

Selector_2 s8414_7(wires_2103_6[2], addr_2103_6, addr_positional[33659:33656], addr_8414_7);

wire[31:0] addr_8415_7;

Selector_2 s8415_7(wires_2103_6[3], addr_2103_6, addr_positional[33663:33660], addr_8415_7);

wire[31:0] addr_8416_7;

Selector_2 s8416_7(wires_2104_6[0], addr_2104_6, addr_positional[33667:33664], addr_8416_7);

wire[31:0] addr_8417_7;

Selector_2 s8417_7(wires_2104_6[1], addr_2104_6, addr_positional[33671:33668], addr_8417_7);

wire[31:0] addr_8418_7;

Selector_2 s8418_7(wires_2104_6[2], addr_2104_6, addr_positional[33675:33672], addr_8418_7);

wire[31:0] addr_8419_7;

Selector_2 s8419_7(wires_2104_6[3], addr_2104_6, addr_positional[33679:33676], addr_8419_7);

wire[31:0] addr_8420_7;

Selector_2 s8420_7(wires_2105_6[0], addr_2105_6, addr_positional[33683:33680], addr_8420_7);

wire[31:0] addr_8421_7;

Selector_2 s8421_7(wires_2105_6[1], addr_2105_6, addr_positional[33687:33684], addr_8421_7);

wire[31:0] addr_8422_7;

Selector_2 s8422_7(wires_2105_6[2], addr_2105_6, addr_positional[33691:33688], addr_8422_7);

wire[31:0] addr_8423_7;

Selector_2 s8423_7(wires_2105_6[3], addr_2105_6, addr_positional[33695:33692], addr_8423_7);

wire[31:0] addr_8424_7;

Selector_2 s8424_7(wires_2106_6[0], addr_2106_6, addr_positional[33699:33696], addr_8424_7);

wire[31:0] addr_8425_7;

Selector_2 s8425_7(wires_2106_6[1], addr_2106_6, addr_positional[33703:33700], addr_8425_7);

wire[31:0] addr_8426_7;

Selector_2 s8426_7(wires_2106_6[2], addr_2106_6, addr_positional[33707:33704], addr_8426_7);

wire[31:0] addr_8427_7;

Selector_2 s8427_7(wires_2106_6[3], addr_2106_6, addr_positional[33711:33708], addr_8427_7);

wire[31:0] addr_8428_7;

Selector_2 s8428_7(wires_2107_6[0], addr_2107_6, addr_positional[33715:33712], addr_8428_7);

wire[31:0] addr_8429_7;

Selector_2 s8429_7(wires_2107_6[1], addr_2107_6, addr_positional[33719:33716], addr_8429_7);

wire[31:0] addr_8430_7;

Selector_2 s8430_7(wires_2107_6[2], addr_2107_6, addr_positional[33723:33720], addr_8430_7);

wire[31:0] addr_8431_7;

Selector_2 s8431_7(wires_2107_6[3], addr_2107_6, addr_positional[33727:33724], addr_8431_7);

wire[31:0] addr_8432_7;

Selector_2 s8432_7(wires_2108_6[0], addr_2108_6, addr_positional[33731:33728], addr_8432_7);

wire[31:0] addr_8433_7;

Selector_2 s8433_7(wires_2108_6[1], addr_2108_6, addr_positional[33735:33732], addr_8433_7);

wire[31:0] addr_8434_7;

Selector_2 s8434_7(wires_2108_6[2], addr_2108_6, addr_positional[33739:33736], addr_8434_7);

wire[31:0] addr_8435_7;

Selector_2 s8435_7(wires_2108_6[3], addr_2108_6, addr_positional[33743:33740], addr_8435_7);

wire[31:0] addr_8436_7;

Selector_2 s8436_7(wires_2109_6[0], addr_2109_6, addr_positional[33747:33744], addr_8436_7);

wire[31:0] addr_8437_7;

Selector_2 s8437_7(wires_2109_6[1], addr_2109_6, addr_positional[33751:33748], addr_8437_7);

wire[31:0] addr_8438_7;

Selector_2 s8438_7(wires_2109_6[2], addr_2109_6, addr_positional[33755:33752], addr_8438_7);

wire[31:0] addr_8439_7;

Selector_2 s8439_7(wires_2109_6[3], addr_2109_6, addr_positional[33759:33756], addr_8439_7);

wire[31:0] addr_8440_7;

Selector_2 s8440_7(wires_2110_6[0], addr_2110_6, addr_positional[33763:33760], addr_8440_7);

wire[31:0] addr_8441_7;

Selector_2 s8441_7(wires_2110_6[1], addr_2110_6, addr_positional[33767:33764], addr_8441_7);

wire[31:0] addr_8442_7;

Selector_2 s8442_7(wires_2110_6[2], addr_2110_6, addr_positional[33771:33768], addr_8442_7);

wire[31:0] addr_8443_7;

Selector_2 s8443_7(wires_2110_6[3], addr_2110_6, addr_positional[33775:33772], addr_8443_7);

wire[31:0] addr_8444_7;

Selector_2 s8444_7(wires_2111_6[0], addr_2111_6, addr_positional[33779:33776], addr_8444_7);

wire[31:0] addr_8445_7;

Selector_2 s8445_7(wires_2111_6[1], addr_2111_6, addr_positional[33783:33780], addr_8445_7);

wire[31:0] addr_8446_7;

Selector_2 s8446_7(wires_2111_6[2], addr_2111_6, addr_positional[33787:33784], addr_8446_7);

wire[31:0] addr_8447_7;

Selector_2 s8447_7(wires_2111_6[3], addr_2111_6, addr_positional[33791:33788], addr_8447_7);

wire[31:0] addr_8448_7;

Selector_2 s8448_7(wires_2112_6[0], addr_2112_6, addr_positional[33795:33792], addr_8448_7);

wire[31:0] addr_8449_7;

Selector_2 s8449_7(wires_2112_6[1], addr_2112_6, addr_positional[33799:33796], addr_8449_7);

wire[31:0] addr_8450_7;

Selector_2 s8450_7(wires_2112_6[2], addr_2112_6, addr_positional[33803:33800], addr_8450_7);

wire[31:0] addr_8451_7;

Selector_2 s8451_7(wires_2112_6[3], addr_2112_6, addr_positional[33807:33804], addr_8451_7);

wire[31:0] addr_8452_7;

Selector_2 s8452_7(wires_2113_6[0], addr_2113_6, addr_positional[33811:33808], addr_8452_7);

wire[31:0] addr_8453_7;

Selector_2 s8453_7(wires_2113_6[1], addr_2113_6, addr_positional[33815:33812], addr_8453_7);

wire[31:0] addr_8454_7;

Selector_2 s8454_7(wires_2113_6[2], addr_2113_6, addr_positional[33819:33816], addr_8454_7);

wire[31:0] addr_8455_7;

Selector_2 s8455_7(wires_2113_6[3], addr_2113_6, addr_positional[33823:33820], addr_8455_7);

wire[31:0] addr_8456_7;

Selector_2 s8456_7(wires_2114_6[0], addr_2114_6, addr_positional[33827:33824], addr_8456_7);

wire[31:0] addr_8457_7;

Selector_2 s8457_7(wires_2114_6[1], addr_2114_6, addr_positional[33831:33828], addr_8457_7);

wire[31:0] addr_8458_7;

Selector_2 s8458_7(wires_2114_6[2], addr_2114_6, addr_positional[33835:33832], addr_8458_7);

wire[31:0] addr_8459_7;

Selector_2 s8459_7(wires_2114_6[3], addr_2114_6, addr_positional[33839:33836], addr_8459_7);

wire[31:0] addr_8460_7;

Selector_2 s8460_7(wires_2115_6[0], addr_2115_6, addr_positional[33843:33840], addr_8460_7);

wire[31:0] addr_8461_7;

Selector_2 s8461_7(wires_2115_6[1], addr_2115_6, addr_positional[33847:33844], addr_8461_7);

wire[31:0] addr_8462_7;

Selector_2 s8462_7(wires_2115_6[2], addr_2115_6, addr_positional[33851:33848], addr_8462_7);

wire[31:0] addr_8463_7;

Selector_2 s8463_7(wires_2115_6[3], addr_2115_6, addr_positional[33855:33852], addr_8463_7);

wire[31:0] addr_8464_7;

Selector_2 s8464_7(wires_2116_6[0], addr_2116_6, addr_positional[33859:33856], addr_8464_7);

wire[31:0] addr_8465_7;

Selector_2 s8465_7(wires_2116_6[1], addr_2116_6, addr_positional[33863:33860], addr_8465_7);

wire[31:0] addr_8466_7;

Selector_2 s8466_7(wires_2116_6[2], addr_2116_6, addr_positional[33867:33864], addr_8466_7);

wire[31:0] addr_8467_7;

Selector_2 s8467_7(wires_2116_6[3], addr_2116_6, addr_positional[33871:33868], addr_8467_7);

wire[31:0] addr_8468_7;

Selector_2 s8468_7(wires_2117_6[0], addr_2117_6, addr_positional[33875:33872], addr_8468_7);

wire[31:0] addr_8469_7;

Selector_2 s8469_7(wires_2117_6[1], addr_2117_6, addr_positional[33879:33876], addr_8469_7);

wire[31:0] addr_8470_7;

Selector_2 s8470_7(wires_2117_6[2], addr_2117_6, addr_positional[33883:33880], addr_8470_7);

wire[31:0] addr_8471_7;

Selector_2 s8471_7(wires_2117_6[3], addr_2117_6, addr_positional[33887:33884], addr_8471_7);

wire[31:0] addr_8472_7;

Selector_2 s8472_7(wires_2118_6[0], addr_2118_6, addr_positional[33891:33888], addr_8472_7);

wire[31:0] addr_8473_7;

Selector_2 s8473_7(wires_2118_6[1], addr_2118_6, addr_positional[33895:33892], addr_8473_7);

wire[31:0] addr_8474_7;

Selector_2 s8474_7(wires_2118_6[2], addr_2118_6, addr_positional[33899:33896], addr_8474_7);

wire[31:0] addr_8475_7;

Selector_2 s8475_7(wires_2118_6[3], addr_2118_6, addr_positional[33903:33900], addr_8475_7);

wire[31:0] addr_8476_7;

Selector_2 s8476_7(wires_2119_6[0], addr_2119_6, addr_positional[33907:33904], addr_8476_7);

wire[31:0] addr_8477_7;

Selector_2 s8477_7(wires_2119_6[1], addr_2119_6, addr_positional[33911:33908], addr_8477_7);

wire[31:0] addr_8478_7;

Selector_2 s8478_7(wires_2119_6[2], addr_2119_6, addr_positional[33915:33912], addr_8478_7);

wire[31:0] addr_8479_7;

Selector_2 s8479_7(wires_2119_6[3], addr_2119_6, addr_positional[33919:33916], addr_8479_7);

wire[31:0] addr_8480_7;

Selector_2 s8480_7(wires_2120_6[0], addr_2120_6, addr_positional[33923:33920], addr_8480_7);

wire[31:0] addr_8481_7;

Selector_2 s8481_7(wires_2120_6[1], addr_2120_6, addr_positional[33927:33924], addr_8481_7);

wire[31:0] addr_8482_7;

Selector_2 s8482_7(wires_2120_6[2], addr_2120_6, addr_positional[33931:33928], addr_8482_7);

wire[31:0] addr_8483_7;

Selector_2 s8483_7(wires_2120_6[3], addr_2120_6, addr_positional[33935:33932], addr_8483_7);

wire[31:0] addr_8484_7;

Selector_2 s8484_7(wires_2121_6[0], addr_2121_6, addr_positional[33939:33936], addr_8484_7);

wire[31:0] addr_8485_7;

Selector_2 s8485_7(wires_2121_6[1], addr_2121_6, addr_positional[33943:33940], addr_8485_7);

wire[31:0] addr_8486_7;

Selector_2 s8486_7(wires_2121_6[2], addr_2121_6, addr_positional[33947:33944], addr_8486_7);

wire[31:0] addr_8487_7;

Selector_2 s8487_7(wires_2121_6[3], addr_2121_6, addr_positional[33951:33948], addr_8487_7);

wire[31:0] addr_8488_7;

Selector_2 s8488_7(wires_2122_6[0], addr_2122_6, addr_positional[33955:33952], addr_8488_7);

wire[31:0] addr_8489_7;

Selector_2 s8489_7(wires_2122_6[1], addr_2122_6, addr_positional[33959:33956], addr_8489_7);

wire[31:0] addr_8490_7;

Selector_2 s8490_7(wires_2122_6[2], addr_2122_6, addr_positional[33963:33960], addr_8490_7);

wire[31:0] addr_8491_7;

Selector_2 s8491_7(wires_2122_6[3], addr_2122_6, addr_positional[33967:33964], addr_8491_7);

wire[31:0] addr_8492_7;

Selector_2 s8492_7(wires_2123_6[0], addr_2123_6, addr_positional[33971:33968], addr_8492_7);

wire[31:0] addr_8493_7;

Selector_2 s8493_7(wires_2123_6[1], addr_2123_6, addr_positional[33975:33972], addr_8493_7);

wire[31:0] addr_8494_7;

Selector_2 s8494_7(wires_2123_6[2], addr_2123_6, addr_positional[33979:33976], addr_8494_7);

wire[31:0] addr_8495_7;

Selector_2 s8495_7(wires_2123_6[3], addr_2123_6, addr_positional[33983:33980], addr_8495_7);

wire[31:0] addr_8496_7;

Selector_2 s8496_7(wires_2124_6[0], addr_2124_6, addr_positional[33987:33984], addr_8496_7);

wire[31:0] addr_8497_7;

Selector_2 s8497_7(wires_2124_6[1], addr_2124_6, addr_positional[33991:33988], addr_8497_7);

wire[31:0] addr_8498_7;

Selector_2 s8498_7(wires_2124_6[2], addr_2124_6, addr_positional[33995:33992], addr_8498_7);

wire[31:0] addr_8499_7;

Selector_2 s8499_7(wires_2124_6[3], addr_2124_6, addr_positional[33999:33996], addr_8499_7);

wire[31:0] addr_8500_7;

Selector_2 s8500_7(wires_2125_6[0], addr_2125_6, addr_positional[34003:34000], addr_8500_7);

wire[31:0] addr_8501_7;

Selector_2 s8501_7(wires_2125_6[1], addr_2125_6, addr_positional[34007:34004], addr_8501_7);

wire[31:0] addr_8502_7;

Selector_2 s8502_7(wires_2125_6[2], addr_2125_6, addr_positional[34011:34008], addr_8502_7);

wire[31:0] addr_8503_7;

Selector_2 s8503_7(wires_2125_6[3], addr_2125_6, addr_positional[34015:34012], addr_8503_7);

wire[31:0] addr_8504_7;

Selector_2 s8504_7(wires_2126_6[0], addr_2126_6, addr_positional[34019:34016], addr_8504_7);

wire[31:0] addr_8505_7;

Selector_2 s8505_7(wires_2126_6[1], addr_2126_6, addr_positional[34023:34020], addr_8505_7);

wire[31:0] addr_8506_7;

Selector_2 s8506_7(wires_2126_6[2], addr_2126_6, addr_positional[34027:34024], addr_8506_7);

wire[31:0] addr_8507_7;

Selector_2 s8507_7(wires_2126_6[3], addr_2126_6, addr_positional[34031:34028], addr_8507_7);

wire[31:0] addr_8508_7;

Selector_2 s8508_7(wires_2127_6[0], addr_2127_6, addr_positional[34035:34032], addr_8508_7);

wire[31:0] addr_8509_7;

Selector_2 s8509_7(wires_2127_6[1], addr_2127_6, addr_positional[34039:34036], addr_8509_7);

wire[31:0] addr_8510_7;

Selector_2 s8510_7(wires_2127_6[2], addr_2127_6, addr_positional[34043:34040], addr_8510_7);

wire[31:0] addr_8511_7;

Selector_2 s8511_7(wires_2127_6[3], addr_2127_6, addr_positional[34047:34044], addr_8511_7);

wire[31:0] addr_8512_7;

Selector_2 s8512_7(wires_2128_6[0], addr_2128_6, addr_positional[34051:34048], addr_8512_7);

wire[31:0] addr_8513_7;

Selector_2 s8513_7(wires_2128_6[1], addr_2128_6, addr_positional[34055:34052], addr_8513_7);

wire[31:0] addr_8514_7;

Selector_2 s8514_7(wires_2128_6[2], addr_2128_6, addr_positional[34059:34056], addr_8514_7);

wire[31:0] addr_8515_7;

Selector_2 s8515_7(wires_2128_6[3], addr_2128_6, addr_positional[34063:34060], addr_8515_7);

wire[31:0] addr_8516_7;

Selector_2 s8516_7(wires_2129_6[0], addr_2129_6, addr_positional[34067:34064], addr_8516_7);

wire[31:0] addr_8517_7;

Selector_2 s8517_7(wires_2129_6[1], addr_2129_6, addr_positional[34071:34068], addr_8517_7);

wire[31:0] addr_8518_7;

Selector_2 s8518_7(wires_2129_6[2], addr_2129_6, addr_positional[34075:34072], addr_8518_7);

wire[31:0] addr_8519_7;

Selector_2 s8519_7(wires_2129_6[3], addr_2129_6, addr_positional[34079:34076], addr_8519_7);

wire[31:0] addr_8520_7;

Selector_2 s8520_7(wires_2130_6[0], addr_2130_6, addr_positional[34083:34080], addr_8520_7);

wire[31:0] addr_8521_7;

Selector_2 s8521_7(wires_2130_6[1], addr_2130_6, addr_positional[34087:34084], addr_8521_7);

wire[31:0] addr_8522_7;

Selector_2 s8522_7(wires_2130_6[2], addr_2130_6, addr_positional[34091:34088], addr_8522_7);

wire[31:0] addr_8523_7;

Selector_2 s8523_7(wires_2130_6[3], addr_2130_6, addr_positional[34095:34092], addr_8523_7);

wire[31:0] addr_8524_7;

Selector_2 s8524_7(wires_2131_6[0], addr_2131_6, addr_positional[34099:34096], addr_8524_7);

wire[31:0] addr_8525_7;

Selector_2 s8525_7(wires_2131_6[1], addr_2131_6, addr_positional[34103:34100], addr_8525_7);

wire[31:0] addr_8526_7;

Selector_2 s8526_7(wires_2131_6[2], addr_2131_6, addr_positional[34107:34104], addr_8526_7);

wire[31:0] addr_8527_7;

Selector_2 s8527_7(wires_2131_6[3], addr_2131_6, addr_positional[34111:34108], addr_8527_7);

wire[31:0] addr_8528_7;

Selector_2 s8528_7(wires_2132_6[0], addr_2132_6, addr_positional[34115:34112], addr_8528_7);

wire[31:0] addr_8529_7;

Selector_2 s8529_7(wires_2132_6[1], addr_2132_6, addr_positional[34119:34116], addr_8529_7);

wire[31:0] addr_8530_7;

Selector_2 s8530_7(wires_2132_6[2], addr_2132_6, addr_positional[34123:34120], addr_8530_7);

wire[31:0] addr_8531_7;

Selector_2 s8531_7(wires_2132_6[3], addr_2132_6, addr_positional[34127:34124], addr_8531_7);

wire[31:0] addr_8532_7;

Selector_2 s8532_7(wires_2133_6[0], addr_2133_6, addr_positional[34131:34128], addr_8532_7);

wire[31:0] addr_8533_7;

Selector_2 s8533_7(wires_2133_6[1], addr_2133_6, addr_positional[34135:34132], addr_8533_7);

wire[31:0] addr_8534_7;

Selector_2 s8534_7(wires_2133_6[2], addr_2133_6, addr_positional[34139:34136], addr_8534_7);

wire[31:0] addr_8535_7;

Selector_2 s8535_7(wires_2133_6[3], addr_2133_6, addr_positional[34143:34140], addr_8535_7);

wire[31:0] addr_8536_7;

Selector_2 s8536_7(wires_2134_6[0], addr_2134_6, addr_positional[34147:34144], addr_8536_7);

wire[31:0] addr_8537_7;

Selector_2 s8537_7(wires_2134_6[1], addr_2134_6, addr_positional[34151:34148], addr_8537_7);

wire[31:0] addr_8538_7;

Selector_2 s8538_7(wires_2134_6[2], addr_2134_6, addr_positional[34155:34152], addr_8538_7);

wire[31:0] addr_8539_7;

Selector_2 s8539_7(wires_2134_6[3], addr_2134_6, addr_positional[34159:34156], addr_8539_7);

wire[31:0] addr_8540_7;

Selector_2 s8540_7(wires_2135_6[0], addr_2135_6, addr_positional[34163:34160], addr_8540_7);

wire[31:0] addr_8541_7;

Selector_2 s8541_7(wires_2135_6[1], addr_2135_6, addr_positional[34167:34164], addr_8541_7);

wire[31:0] addr_8542_7;

Selector_2 s8542_7(wires_2135_6[2], addr_2135_6, addr_positional[34171:34168], addr_8542_7);

wire[31:0] addr_8543_7;

Selector_2 s8543_7(wires_2135_6[3], addr_2135_6, addr_positional[34175:34172], addr_8543_7);

wire[31:0] addr_8544_7;

Selector_2 s8544_7(wires_2136_6[0], addr_2136_6, addr_positional[34179:34176], addr_8544_7);

wire[31:0] addr_8545_7;

Selector_2 s8545_7(wires_2136_6[1], addr_2136_6, addr_positional[34183:34180], addr_8545_7);

wire[31:0] addr_8546_7;

Selector_2 s8546_7(wires_2136_6[2], addr_2136_6, addr_positional[34187:34184], addr_8546_7);

wire[31:0] addr_8547_7;

Selector_2 s8547_7(wires_2136_6[3], addr_2136_6, addr_positional[34191:34188], addr_8547_7);

wire[31:0] addr_8548_7;

Selector_2 s8548_7(wires_2137_6[0], addr_2137_6, addr_positional[34195:34192], addr_8548_7);

wire[31:0] addr_8549_7;

Selector_2 s8549_7(wires_2137_6[1], addr_2137_6, addr_positional[34199:34196], addr_8549_7);

wire[31:0] addr_8550_7;

Selector_2 s8550_7(wires_2137_6[2], addr_2137_6, addr_positional[34203:34200], addr_8550_7);

wire[31:0] addr_8551_7;

Selector_2 s8551_7(wires_2137_6[3], addr_2137_6, addr_positional[34207:34204], addr_8551_7);

wire[31:0] addr_8552_7;

Selector_2 s8552_7(wires_2138_6[0], addr_2138_6, addr_positional[34211:34208], addr_8552_7);

wire[31:0] addr_8553_7;

Selector_2 s8553_7(wires_2138_6[1], addr_2138_6, addr_positional[34215:34212], addr_8553_7);

wire[31:0] addr_8554_7;

Selector_2 s8554_7(wires_2138_6[2], addr_2138_6, addr_positional[34219:34216], addr_8554_7);

wire[31:0] addr_8555_7;

Selector_2 s8555_7(wires_2138_6[3], addr_2138_6, addr_positional[34223:34220], addr_8555_7);

wire[31:0] addr_8556_7;

Selector_2 s8556_7(wires_2139_6[0], addr_2139_6, addr_positional[34227:34224], addr_8556_7);

wire[31:0] addr_8557_7;

Selector_2 s8557_7(wires_2139_6[1], addr_2139_6, addr_positional[34231:34228], addr_8557_7);

wire[31:0] addr_8558_7;

Selector_2 s8558_7(wires_2139_6[2], addr_2139_6, addr_positional[34235:34232], addr_8558_7);

wire[31:0] addr_8559_7;

Selector_2 s8559_7(wires_2139_6[3], addr_2139_6, addr_positional[34239:34236], addr_8559_7);

wire[31:0] addr_8560_7;

Selector_2 s8560_7(wires_2140_6[0], addr_2140_6, addr_positional[34243:34240], addr_8560_7);

wire[31:0] addr_8561_7;

Selector_2 s8561_7(wires_2140_6[1], addr_2140_6, addr_positional[34247:34244], addr_8561_7);

wire[31:0] addr_8562_7;

Selector_2 s8562_7(wires_2140_6[2], addr_2140_6, addr_positional[34251:34248], addr_8562_7);

wire[31:0] addr_8563_7;

Selector_2 s8563_7(wires_2140_6[3], addr_2140_6, addr_positional[34255:34252], addr_8563_7);

wire[31:0] addr_8564_7;

Selector_2 s8564_7(wires_2141_6[0], addr_2141_6, addr_positional[34259:34256], addr_8564_7);

wire[31:0] addr_8565_7;

Selector_2 s8565_7(wires_2141_6[1], addr_2141_6, addr_positional[34263:34260], addr_8565_7);

wire[31:0] addr_8566_7;

Selector_2 s8566_7(wires_2141_6[2], addr_2141_6, addr_positional[34267:34264], addr_8566_7);

wire[31:0] addr_8567_7;

Selector_2 s8567_7(wires_2141_6[3], addr_2141_6, addr_positional[34271:34268], addr_8567_7);

wire[31:0] addr_8568_7;

Selector_2 s8568_7(wires_2142_6[0], addr_2142_6, addr_positional[34275:34272], addr_8568_7);

wire[31:0] addr_8569_7;

Selector_2 s8569_7(wires_2142_6[1], addr_2142_6, addr_positional[34279:34276], addr_8569_7);

wire[31:0] addr_8570_7;

Selector_2 s8570_7(wires_2142_6[2], addr_2142_6, addr_positional[34283:34280], addr_8570_7);

wire[31:0] addr_8571_7;

Selector_2 s8571_7(wires_2142_6[3], addr_2142_6, addr_positional[34287:34284], addr_8571_7);

wire[31:0] addr_8572_7;

Selector_2 s8572_7(wires_2143_6[0], addr_2143_6, addr_positional[34291:34288], addr_8572_7);

wire[31:0] addr_8573_7;

Selector_2 s8573_7(wires_2143_6[1], addr_2143_6, addr_positional[34295:34292], addr_8573_7);

wire[31:0] addr_8574_7;

Selector_2 s8574_7(wires_2143_6[2], addr_2143_6, addr_positional[34299:34296], addr_8574_7);

wire[31:0] addr_8575_7;

Selector_2 s8575_7(wires_2143_6[3], addr_2143_6, addr_positional[34303:34300], addr_8575_7);

wire[31:0] addr_8576_7;

Selector_2 s8576_7(wires_2144_6[0], addr_2144_6, addr_positional[34307:34304], addr_8576_7);

wire[31:0] addr_8577_7;

Selector_2 s8577_7(wires_2144_6[1], addr_2144_6, addr_positional[34311:34308], addr_8577_7);

wire[31:0] addr_8578_7;

Selector_2 s8578_7(wires_2144_6[2], addr_2144_6, addr_positional[34315:34312], addr_8578_7);

wire[31:0] addr_8579_7;

Selector_2 s8579_7(wires_2144_6[3], addr_2144_6, addr_positional[34319:34316], addr_8579_7);

wire[31:0] addr_8580_7;

Selector_2 s8580_7(wires_2145_6[0], addr_2145_6, addr_positional[34323:34320], addr_8580_7);

wire[31:0] addr_8581_7;

Selector_2 s8581_7(wires_2145_6[1], addr_2145_6, addr_positional[34327:34324], addr_8581_7);

wire[31:0] addr_8582_7;

Selector_2 s8582_7(wires_2145_6[2], addr_2145_6, addr_positional[34331:34328], addr_8582_7);

wire[31:0] addr_8583_7;

Selector_2 s8583_7(wires_2145_6[3], addr_2145_6, addr_positional[34335:34332], addr_8583_7);

wire[31:0] addr_8584_7;

Selector_2 s8584_7(wires_2146_6[0], addr_2146_6, addr_positional[34339:34336], addr_8584_7);

wire[31:0] addr_8585_7;

Selector_2 s8585_7(wires_2146_6[1], addr_2146_6, addr_positional[34343:34340], addr_8585_7);

wire[31:0] addr_8586_7;

Selector_2 s8586_7(wires_2146_6[2], addr_2146_6, addr_positional[34347:34344], addr_8586_7);

wire[31:0] addr_8587_7;

Selector_2 s8587_7(wires_2146_6[3], addr_2146_6, addr_positional[34351:34348], addr_8587_7);

wire[31:0] addr_8588_7;

Selector_2 s8588_7(wires_2147_6[0], addr_2147_6, addr_positional[34355:34352], addr_8588_7);

wire[31:0] addr_8589_7;

Selector_2 s8589_7(wires_2147_6[1], addr_2147_6, addr_positional[34359:34356], addr_8589_7);

wire[31:0] addr_8590_7;

Selector_2 s8590_7(wires_2147_6[2], addr_2147_6, addr_positional[34363:34360], addr_8590_7);

wire[31:0] addr_8591_7;

Selector_2 s8591_7(wires_2147_6[3], addr_2147_6, addr_positional[34367:34364], addr_8591_7);

wire[31:0] addr_8592_7;

Selector_2 s8592_7(wires_2148_6[0], addr_2148_6, addr_positional[34371:34368], addr_8592_7);

wire[31:0] addr_8593_7;

Selector_2 s8593_7(wires_2148_6[1], addr_2148_6, addr_positional[34375:34372], addr_8593_7);

wire[31:0] addr_8594_7;

Selector_2 s8594_7(wires_2148_6[2], addr_2148_6, addr_positional[34379:34376], addr_8594_7);

wire[31:0] addr_8595_7;

Selector_2 s8595_7(wires_2148_6[3], addr_2148_6, addr_positional[34383:34380], addr_8595_7);

wire[31:0] addr_8596_7;

Selector_2 s8596_7(wires_2149_6[0], addr_2149_6, addr_positional[34387:34384], addr_8596_7);

wire[31:0] addr_8597_7;

Selector_2 s8597_7(wires_2149_6[1], addr_2149_6, addr_positional[34391:34388], addr_8597_7);

wire[31:0] addr_8598_7;

Selector_2 s8598_7(wires_2149_6[2], addr_2149_6, addr_positional[34395:34392], addr_8598_7);

wire[31:0] addr_8599_7;

Selector_2 s8599_7(wires_2149_6[3], addr_2149_6, addr_positional[34399:34396], addr_8599_7);

wire[31:0] addr_8600_7;

Selector_2 s8600_7(wires_2150_6[0], addr_2150_6, addr_positional[34403:34400], addr_8600_7);

wire[31:0] addr_8601_7;

Selector_2 s8601_7(wires_2150_6[1], addr_2150_6, addr_positional[34407:34404], addr_8601_7);

wire[31:0] addr_8602_7;

Selector_2 s8602_7(wires_2150_6[2], addr_2150_6, addr_positional[34411:34408], addr_8602_7);

wire[31:0] addr_8603_7;

Selector_2 s8603_7(wires_2150_6[3], addr_2150_6, addr_positional[34415:34412], addr_8603_7);

wire[31:0] addr_8604_7;

Selector_2 s8604_7(wires_2151_6[0], addr_2151_6, addr_positional[34419:34416], addr_8604_7);

wire[31:0] addr_8605_7;

Selector_2 s8605_7(wires_2151_6[1], addr_2151_6, addr_positional[34423:34420], addr_8605_7);

wire[31:0] addr_8606_7;

Selector_2 s8606_7(wires_2151_6[2], addr_2151_6, addr_positional[34427:34424], addr_8606_7);

wire[31:0] addr_8607_7;

Selector_2 s8607_7(wires_2151_6[3], addr_2151_6, addr_positional[34431:34428], addr_8607_7);

wire[31:0] addr_8608_7;

Selector_2 s8608_7(wires_2152_6[0], addr_2152_6, addr_positional[34435:34432], addr_8608_7);

wire[31:0] addr_8609_7;

Selector_2 s8609_7(wires_2152_6[1], addr_2152_6, addr_positional[34439:34436], addr_8609_7);

wire[31:0] addr_8610_7;

Selector_2 s8610_7(wires_2152_6[2], addr_2152_6, addr_positional[34443:34440], addr_8610_7);

wire[31:0] addr_8611_7;

Selector_2 s8611_7(wires_2152_6[3], addr_2152_6, addr_positional[34447:34444], addr_8611_7);

wire[31:0] addr_8612_7;

Selector_2 s8612_7(wires_2153_6[0], addr_2153_6, addr_positional[34451:34448], addr_8612_7);

wire[31:0] addr_8613_7;

Selector_2 s8613_7(wires_2153_6[1], addr_2153_6, addr_positional[34455:34452], addr_8613_7);

wire[31:0] addr_8614_7;

Selector_2 s8614_7(wires_2153_6[2], addr_2153_6, addr_positional[34459:34456], addr_8614_7);

wire[31:0] addr_8615_7;

Selector_2 s8615_7(wires_2153_6[3], addr_2153_6, addr_positional[34463:34460], addr_8615_7);

wire[31:0] addr_8616_7;

Selector_2 s8616_7(wires_2154_6[0], addr_2154_6, addr_positional[34467:34464], addr_8616_7);

wire[31:0] addr_8617_7;

Selector_2 s8617_7(wires_2154_6[1], addr_2154_6, addr_positional[34471:34468], addr_8617_7);

wire[31:0] addr_8618_7;

Selector_2 s8618_7(wires_2154_6[2], addr_2154_6, addr_positional[34475:34472], addr_8618_7);

wire[31:0] addr_8619_7;

Selector_2 s8619_7(wires_2154_6[3], addr_2154_6, addr_positional[34479:34476], addr_8619_7);

wire[31:0] addr_8620_7;

Selector_2 s8620_7(wires_2155_6[0], addr_2155_6, addr_positional[34483:34480], addr_8620_7);

wire[31:0] addr_8621_7;

Selector_2 s8621_7(wires_2155_6[1], addr_2155_6, addr_positional[34487:34484], addr_8621_7);

wire[31:0] addr_8622_7;

Selector_2 s8622_7(wires_2155_6[2], addr_2155_6, addr_positional[34491:34488], addr_8622_7);

wire[31:0] addr_8623_7;

Selector_2 s8623_7(wires_2155_6[3], addr_2155_6, addr_positional[34495:34492], addr_8623_7);

wire[31:0] addr_8624_7;

Selector_2 s8624_7(wires_2156_6[0], addr_2156_6, addr_positional[34499:34496], addr_8624_7);

wire[31:0] addr_8625_7;

Selector_2 s8625_7(wires_2156_6[1], addr_2156_6, addr_positional[34503:34500], addr_8625_7);

wire[31:0] addr_8626_7;

Selector_2 s8626_7(wires_2156_6[2], addr_2156_6, addr_positional[34507:34504], addr_8626_7);

wire[31:0] addr_8627_7;

Selector_2 s8627_7(wires_2156_6[3], addr_2156_6, addr_positional[34511:34508], addr_8627_7);

wire[31:0] addr_8628_7;

Selector_2 s8628_7(wires_2157_6[0], addr_2157_6, addr_positional[34515:34512], addr_8628_7);

wire[31:0] addr_8629_7;

Selector_2 s8629_7(wires_2157_6[1], addr_2157_6, addr_positional[34519:34516], addr_8629_7);

wire[31:0] addr_8630_7;

Selector_2 s8630_7(wires_2157_6[2], addr_2157_6, addr_positional[34523:34520], addr_8630_7);

wire[31:0] addr_8631_7;

Selector_2 s8631_7(wires_2157_6[3], addr_2157_6, addr_positional[34527:34524], addr_8631_7);

wire[31:0] addr_8632_7;

Selector_2 s8632_7(wires_2158_6[0], addr_2158_6, addr_positional[34531:34528], addr_8632_7);

wire[31:0] addr_8633_7;

Selector_2 s8633_7(wires_2158_6[1], addr_2158_6, addr_positional[34535:34532], addr_8633_7);

wire[31:0] addr_8634_7;

Selector_2 s8634_7(wires_2158_6[2], addr_2158_6, addr_positional[34539:34536], addr_8634_7);

wire[31:0] addr_8635_7;

Selector_2 s8635_7(wires_2158_6[3], addr_2158_6, addr_positional[34543:34540], addr_8635_7);

wire[31:0] addr_8636_7;

Selector_2 s8636_7(wires_2159_6[0], addr_2159_6, addr_positional[34547:34544], addr_8636_7);

wire[31:0] addr_8637_7;

Selector_2 s8637_7(wires_2159_6[1], addr_2159_6, addr_positional[34551:34548], addr_8637_7);

wire[31:0] addr_8638_7;

Selector_2 s8638_7(wires_2159_6[2], addr_2159_6, addr_positional[34555:34552], addr_8638_7);

wire[31:0] addr_8639_7;

Selector_2 s8639_7(wires_2159_6[3], addr_2159_6, addr_positional[34559:34556], addr_8639_7);

wire[31:0] addr_8640_7;

Selector_2 s8640_7(wires_2160_6[0], addr_2160_6, addr_positional[34563:34560], addr_8640_7);

wire[31:0] addr_8641_7;

Selector_2 s8641_7(wires_2160_6[1], addr_2160_6, addr_positional[34567:34564], addr_8641_7);

wire[31:0] addr_8642_7;

Selector_2 s8642_7(wires_2160_6[2], addr_2160_6, addr_positional[34571:34568], addr_8642_7);

wire[31:0] addr_8643_7;

Selector_2 s8643_7(wires_2160_6[3], addr_2160_6, addr_positional[34575:34572], addr_8643_7);

wire[31:0] addr_8644_7;

Selector_2 s8644_7(wires_2161_6[0], addr_2161_6, addr_positional[34579:34576], addr_8644_7);

wire[31:0] addr_8645_7;

Selector_2 s8645_7(wires_2161_6[1], addr_2161_6, addr_positional[34583:34580], addr_8645_7);

wire[31:0] addr_8646_7;

Selector_2 s8646_7(wires_2161_6[2], addr_2161_6, addr_positional[34587:34584], addr_8646_7);

wire[31:0] addr_8647_7;

Selector_2 s8647_7(wires_2161_6[3], addr_2161_6, addr_positional[34591:34588], addr_8647_7);

wire[31:0] addr_8648_7;

Selector_2 s8648_7(wires_2162_6[0], addr_2162_6, addr_positional[34595:34592], addr_8648_7);

wire[31:0] addr_8649_7;

Selector_2 s8649_7(wires_2162_6[1], addr_2162_6, addr_positional[34599:34596], addr_8649_7);

wire[31:0] addr_8650_7;

Selector_2 s8650_7(wires_2162_6[2], addr_2162_6, addr_positional[34603:34600], addr_8650_7);

wire[31:0] addr_8651_7;

Selector_2 s8651_7(wires_2162_6[3], addr_2162_6, addr_positional[34607:34604], addr_8651_7);

wire[31:0] addr_8652_7;

Selector_2 s8652_7(wires_2163_6[0], addr_2163_6, addr_positional[34611:34608], addr_8652_7);

wire[31:0] addr_8653_7;

Selector_2 s8653_7(wires_2163_6[1], addr_2163_6, addr_positional[34615:34612], addr_8653_7);

wire[31:0] addr_8654_7;

Selector_2 s8654_7(wires_2163_6[2], addr_2163_6, addr_positional[34619:34616], addr_8654_7);

wire[31:0] addr_8655_7;

Selector_2 s8655_7(wires_2163_6[3], addr_2163_6, addr_positional[34623:34620], addr_8655_7);

wire[31:0] addr_8656_7;

Selector_2 s8656_7(wires_2164_6[0], addr_2164_6, addr_positional[34627:34624], addr_8656_7);

wire[31:0] addr_8657_7;

Selector_2 s8657_7(wires_2164_6[1], addr_2164_6, addr_positional[34631:34628], addr_8657_7);

wire[31:0] addr_8658_7;

Selector_2 s8658_7(wires_2164_6[2], addr_2164_6, addr_positional[34635:34632], addr_8658_7);

wire[31:0] addr_8659_7;

Selector_2 s8659_7(wires_2164_6[3], addr_2164_6, addr_positional[34639:34636], addr_8659_7);

wire[31:0] addr_8660_7;

Selector_2 s8660_7(wires_2165_6[0], addr_2165_6, addr_positional[34643:34640], addr_8660_7);

wire[31:0] addr_8661_7;

Selector_2 s8661_7(wires_2165_6[1], addr_2165_6, addr_positional[34647:34644], addr_8661_7);

wire[31:0] addr_8662_7;

Selector_2 s8662_7(wires_2165_6[2], addr_2165_6, addr_positional[34651:34648], addr_8662_7);

wire[31:0] addr_8663_7;

Selector_2 s8663_7(wires_2165_6[3], addr_2165_6, addr_positional[34655:34652], addr_8663_7);

wire[31:0] addr_8664_7;

Selector_2 s8664_7(wires_2166_6[0], addr_2166_6, addr_positional[34659:34656], addr_8664_7);

wire[31:0] addr_8665_7;

Selector_2 s8665_7(wires_2166_6[1], addr_2166_6, addr_positional[34663:34660], addr_8665_7);

wire[31:0] addr_8666_7;

Selector_2 s8666_7(wires_2166_6[2], addr_2166_6, addr_positional[34667:34664], addr_8666_7);

wire[31:0] addr_8667_7;

Selector_2 s8667_7(wires_2166_6[3], addr_2166_6, addr_positional[34671:34668], addr_8667_7);

wire[31:0] addr_8668_7;

Selector_2 s8668_7(wires_2167_6[0], addr_2167_6, addr_positional[34675:34672], addr_8668_7);

wire[31:0] addr_8669_7;

Selector_2 s8669_7(wires_2167_6[1], addr_2167_6, addr_positional[34679:34676], addr_8669_7);

wire[31:0] addr_8670_7;

Selector_2 s8670_7(wires_2167_6[2], addr_2167_6, addr_positional[34683:34680], addr_8670_7);

wire[31:0] addr_8671_7;

Selector_2 s8671_7(wires_2167_6[3], addr_2167_6, addr_positional[34687:34684], addr_8671_7);

wire[31:0] addr_8672_7;

Selector_2 s8672_7(wires_2168_6[0], addr_2168_6, addr_positional[34691:34688], addr_8672_7);

wire[31:0] addr_8673_7;

Selector_2 s8673_7(wires_2168_6[1], addr_2168_6, addr_positional[34695:34692], addr_8673_7);

wire[31:0] addr_8674_7;

Selector_2 s8674_7(wires_2168_6[2], addr_2168_6, addr_positional[34699:34696], addr_8674_7);

wire[31:0] addr_8675_7;

Selector_2 s8675_7(wires_2168_6[3], addr_2168_6, addr_positional[34703:34700], addr_8675_7);

wire[31:0] addr_8676_7;

Selector_2 s8676_7(wires_2169_6[0], addr_2169_6, addr_positional[34707:34704], addr_8676_7);

wire[31:0] addr_8677_7;

Selector_2 s8677_7(wires_2169_6[1], addr_2169_6, addr_positional[34711:34708], addr_8677_7);

wire[31:0] addr_8678_7;

Selector_2 s8678_7(wires_2169_6[2], addr_2169_6, addr_positional[34715:34712], addr_8678_7);

wire[31:0] addr_8679_7;

Selector_2 s8679_7(wires_2169_6[3], addr_2169_6, addr_positional[34719:34716], addr_8679_7);

wire[31:0] addr_8680_7;

Selector_2 s8680_7(wires_2170_6[0], addr_2170_6, addr_positional[34723:34720], addr_8680_7);

wire[31:0] addr_8681_7;

Selector_2 s8681_7(wires_2170_6[1], addr_2170_6, addr_positional[34727:34724], addr_8681_7);

wire[31:0] addr_8682_7;

Selector_2 s8682_7(wires_2170_6[2], addr_2170_6, addr_positional[34731:34728], addr_8682_7);

wire[31:0] addr_8683_7;

Selector_2 s8683_7(wires_2170_6[3], addr_2170_6, addr_positional[34735:34732], addr_8683_7);

wire[31:0] addr_8684_7;

Selector_2 s8684_7(wires_2171_6[0], addr_2171_6, addr_positional[34739:34736], addr_8684_7);

wire[31:0] addr_8685_7;

Selector_2 s8685_7(wires_2171_6[1], addr_2171_6, addr_positional[34743:34740], addr_8685_7);

wire[31:0] addr_8686_7;

Selector_2 s8686_7(wires_2171_6[2], addr_2171_6, addr_positional[34747:34744], addr_8686_7);

wire[31:0] addr_8687_7;

Selector_2 s8687_7(wires_2171_6[3], addr_2171_6, addr_positional[34751:34748], addr_8687_7);

wire[31:0] addr_8688_7;

Selector_2 s8688_7(wires_2172_6[0], addr_2172_6, addr_positional[34755:34752], addr_8688_7);

wire[31:0] addr_8689_7;

Selector_2 s8689_7(wires_2172_6[1], addr_2172_6, addr_positional[34759:34756], addr_8689_7);

wire[31:0] addr_8690_7;

Selector_2 s8690_7(wires_2172_6[2], addr_2172_6, addr_positional[34763:34760], addr_8690_7);

wire[31:0] addr_8691_7;

Selector_2 s8691_7(wires_2172_6[3], addr_2172_6, addr_positional[34767:34764], addr_8691_7);

wire[31:0] addr_8692_7;

Selector_2 s8692_7(wires_2173_6[0], addr_2173_6, addr_positional[34771:34768], addr_8692_7);

wire[31:0] addr_8693_7;

Selector_2 s8693_7(wires_2173_6[1], addr_2173_6, addr_positional[34775:34772], addr_8693_7);

wire[31:0] addr_8694_7;

Selector_2 s8694_7(wires_2173_6[2], addr_2173_6, addr_positional[34779:34776], addr_8694_7);

wire[31:0] addr_8695_7;

Selector_2 s8695_7(wires_2173_6[3], addr_2173_6, addr_positional[34783:34780], addr_8695_7);

wire[31:0] addr_8696_7;

Selector_2 s8696_7(wires_2174_6[0], addr_2174_6, addr_positional[34787:34784], addr_8696_7);

wire[31:0] addr_8697_7;

Selector_2 s8697_7(wires_2174_6[1], addr_2174_6, addr_positional[34791:34788], addr_8697_7);

wire[31:0] addr_8698_7;

Selector_2 s8698_7(wires_2174_6[2], addr_2174_6, addr_positional[34795:34792], addr_8698_7);

wire[31:0] addr_8699_7;

Selector_2 s8699_7(wires_2174_6[3], addr_2174_6, addr_positional[34799:34796], addr_8699_7);

wire[31:0] addr_8700_7;

Selector_2 s8700_7(wires_2175_6[0], addr_2175_6, addr_positional[34803:34800], addr_8700_7);

wire[31:0] addr_8701_7;

Selector_2 s8701_7(wires_2175_6[1], addr_2175_6, addr_positional[34807:34804], addr_8701_7);

wire[31:0] addr_8702_7;

Selector_2 s8702_7(wires_2175_6[2], addr_2175_6, addr_positional[34811:34808], addr_8702_7);

wire[31:0] addr_8703_7;

Selector_2 s8703_7(wires_2175_6[3], addr_2175_6, addr_positional[34815:34812], addr_8703_7);

wire[31:0] addr_8704_7;

Selector_2 s8704_7(wires_2176_6[0], addr_2176_6, addr_positional[34819:34816], addr_8704_7);

wire[31:0] addr_8705_7;

Selector_2 s8705_7(wires_2176_6[1], addr_2176_6, addr_positional[34823:34820], addr_8705_7);

wire[31:0] addr_8706_7;

Selector_2 s8706_7(wires_2176_6[2], addr_2176_6, addr_positional[34827:34824], addr_8706_7);

wire[31:0] addr_8707_7;

Selector_2 s8707_7(wires_2176_6[3], addr_2176_6, addr_positional[34831:34828], addr_8707_7);

wire[31:0] addr_8708_7;

Selector_2 s8708_7(wires_2177_6[0], addr_2177_6, addr_positional[34835:34832], addr_8708_7);

wire[31:0] addr_8709_7;

Selector_2 s8709_7(wires_2177_6[1], addr_2177_6, addr_positional[34839:34836], addr_8709_7);

wire[31:0] addr_8710_7;

Selector_2 s8710_7(wires_2177_6[2], addr_2177_6, addr_positional[34843:34840], addr_8710_7);

wire[31:0] addr_8711_7;

Selector_2 s8711_7(wires_2177_6[3], addr_2177_6, addr_positional[34847:34844], addr_8711_7);

wire[31:0] addr_8712_7;

Selector_2 s8712_7(wires_2178_6[0], addr_2178_6, addr_positional[34851:34848], addr_8712_7);

wire[31:0] addr_8713_7;

Selector_2 s8713_7(wires_2178_6[1], addr_2178_6, addr_positional[34855:34852], addr_8713_7);

wire[31:0] addr_8714_7;

Selector_2 s8714_7(wires_2178_6[2], addr_2178_6, addr_positional[34859:34856], addr_8714_7);

wire[31:0] addr_8715_7;

Selector_2 s8715_7(wires_2178_6[3], addr_2178_6, addr_positional[34863:34860], addr_8715_7);

wire[31:0] addr_8716_7;

Selector_2 s8716_7(wires_2179_6[0], addr_2179_6, addr_positional[34867:34864], addr_8716_7);

wire[31:0] addr_8717_7;

Selector_2 s8717_7(wires_2179_6[1], addr_2179_6, addr_positional[34871:34868], addr_8717_7);

wire[31:0] addr_8718_7;

Selector_2 s8718_7(wires_2179_6[2], addr_2179_6, addr_positional[34875:34872], addr_8718_7);

wire[31:0] addr_8719_7;

Selector_2 s8719_7(wires_2179_6[3], addr_2179_6, addr_positional[34879:34876], addr_8719_7);

wire[31:0] addr_8720_7;

Selector_2 s8720_7(wires_2180_6[0], addr_2180_6, addr_positional[34883:34880], addr_8720_7);

wire[31:0] addr_8721_7;

Selector_2 s8721_7(wires_2180_6[1], addr_2180_6, addr_positional[34887:34884], addr_8721_7);

wire[31:0] addr_8722_7;

Selector_2 s8722_7(wires_2180_6[2], addr_2180_6, addr_positional[34891:34888], addr_8722_7);

wire[31:0] addr_8723_7;

Selector_2 s8723_7(wires_2180_6[3], addr_2180_6, addr_positional[34895:34892], addr_8723_7);

wire[31:0] addr_8724_7;

Selector_2 s8724_7(wires_2181_6[0], addr_2181_6, addr_positional[34899:34896], addr_8724_7);

wire[31:0] addr_8725_7;

Selector_2 s8725_7(wires_2181_6[1], addr_2181_6, addr_positional[34903:34900], addr_8725_7);

wire[31:0] addr_8726_7;

Selector_2 s8726_7(wires_2181_6[2], addr_2181_6, addr_positional[34907:34904], addr_8726_7);

wire[31:0] addr_8727_7;

Selector_2 s8727_7(wires_2181_6[3], addr_2181_6, addr_positional[34911:34908], addr_8727_7);

wire[31:0] addr_8728_7;

Selector_2 s8728_7(wires_2182_6[0], addr_2182_6, addr_positional[34915:34912], addr_8728_7);

wire[31:0] addr_8729_7;

Selector_2 s8729_7(wires_2182_6[1], addr_2182_6, addr_positional[34919:34916], addr_8729_7);

wire[31:0] addr_8730_7;

Selector_2 s8730_7(wires_2182_6[2], addr_2182_6, addr_positional[34923:34920], addr_8730_7);

wire[31:0] addr_8731_7;

Selector_2 s8731_7(wires_2182_6[3], addr_2182_6, addr_positional[34927:34924], addr_8731_7);

wire[31:0] addr_8732_7;

Selector_2 s8732_7(wires_2183_6[0], addr_2183_6, addr_positional[34931:34928], addr_8732_7);

wire[31:0] addr_8733_7;

Selector_2 s8733_7(wires_2183_6[1], addr_2183_6, addr_positional[34935:34932], addr_8733_7);

wire[31:0] addr_8734_7;

Selector_2 s8734_7(wires_2183_6[2], addr_2183_6, addr_positional[34939:34936], addr_8734_7);

wire[31:0] addr_8735_7;

Selector_2 s8735_7(wires_2183_6[3], addr_2183_6, addr_positional[34943:34940], addr_8735_7);

wire[31:0] addr_8736_7;

Selector_2 s8736_7(wires_2184_6[0], addr_2184_6, addr_positional[34947:34944], addr_8736_7);

wire[31:0] addr_8737_7;

Selector_2 s8737_7(wires_2184_6[1], addr_2184_6, addr_positional[34951:34948], addr_8737_7);

wire[31:0] addr_8738_7;

Selector_2 s8738_7(wires_2184_6[2], addr_2184_6, addr_positional[34955:34952], addr_8738_7);

wire[31:0] addr_8739_7;

Selector_2 s8739_7(wires_2184_6[3], addr_2184_6, addr_positional[34959:34956], addr_8739_7);

wire[31:0] addr_8740_7;

Selector_2 s8740_7(wires_2185_6[0], addr_2185_6, addr_positional[34963:34960], addr_8740_7);

wire[31:0] addr_8741_7;

Selector_2 s8741_7(wires_2185_6[1], addr_2185_6, addr_positional[34967:34964], addr_8741_7);

wire[31:0] addr_8742_7;

Selector_2 s8742_7(wires_2185_6[2], addr_2185_6, addr_positional[34971:34968], addr_8742_7);

wire[31:0] addr_8743_7;

Selector_2 s8743_7(wires_2185_6[3], addr_2185_6, addr_positional[34975:34972], addr_8743_7);

wire[31:0] addr_8744_7;

Selector_2 s8744_7(wires_2186_6[0], addr_2186_6, addr_positional[34979:34976], addr_8744_7);

wire[31:0] addr_8745_7;

Selector_2 s8745_7(wires_2186_6[1], addr_2186_6, addr_positional[34983:34980], addr_8745_7);

wire[31:0] addr_8746_7;

Selector_2 s8746_7(wires_2186_6[2], addr_2186_6, addr_positional[34987:34984], addr_8746_7);

wire[31:0] addr_8747_7;

Selector_2 s8747_7(wires_2186_6[3], addr_2186_6, addr_positional[34991:34988], addr_8747_7);

wire[31:0] addr_8748_7;

Selector_2 s8748_7(wires_2187_6[0], addr_2187_6, addr_positional[34995:34992], addr_8748_7);

wire[31:0] addr_8749_7;

Selector_2 s8749_7(wires_2187_6[1], addr_2187_6, addr_positional[34999:34996], addr_8749_7);

wire[31:0] addr_8750_7;

Selector_2 s8750_7(wires_2187_6[2], addr_2187_6, addr_positional[35003:35000], addr_8750_7);

wire[31:0] addr_8751_7;

Selector_2 s8751_7(wires_2187_6[3], addr_2187_6, addr_positional[35007:35004], addr_8751_7);

wire[31:0] addr_8752_7;

Selector_2 s8752_7(wires_2188_6[0], addr_2188_6, addr_positional[35011:35008], addr_8752_7);

wire[31:0] addr_8753_7;

Selector_2 s8753_7(wires_2188_6[1], addr_2188_6, addr_positional[35015:35012], addr_8753_7);

wire[31:0] addr_8754_7;

Selector_2 s8754_7(wires_2188_6[2], addr_2188_6, addr_positional[35019:35016], addr_8754_7);

wire[31:0] addr_8755_7;

Selector_2 s8755_7(wires_2188_6[3], addr_2188_6, addr_positional[35023:35020], addr_8755_7);

wire[31:0] addr_8756_7;

Selector_2 s8756_7(wires_2189_6[0], addr_2189_6, addr_positional[35027:35024], addr_8756_7);

wire[31:0] addr_8757_7;

Selector_2 s8757_7(wires_2189_6[1], addr_2189_6, addr_positional[35031:35028], addr_8757_7);

wire[31:0] addr_8758_7;

Selector_2 s8758_7(wires_2189_6[2], addr_2189_6, addr_positional[35035:35032], addr_8758_7);

wire[31:0] addr_8759_7;

Selector_2 s8759_7(wires_2189_6[3], addr_2189_6, addr_positional[35039:35036], addr_8759_7);

wire[31:0] addr_8760_7;

Selector_2 s8760_7(wires_2190_6[0], addr_2190_6, addr_positional[35043:35040], addr_8760_7);

wire[31:0] addr_8761_7;

Selector_2 s8761_7(wires_2190_6[1], addr_2190_6, addr_positional[35047:35044], addr_8761_7);

wire[31:0] addr_8762_7;

Selector_2 s8762_7(wires_2190_6[2], addr_2190_6, addr_positional[35051:35048], addr_8762_7);

wire[31:0] addr_8763_7;

Selector_2 s8763_7(wires_2190_6[3], addr_2190_6, addr_positional[35055:35052], addr_8763_7);

wire[31:0] addr_8764_7;

Selector_2 s8764_7(wires_2191_6[0], addr_2191_6, addr_positional[35059:35056], addr_8764_7);

wire[31:0] addr_8765_7;

Selector_2 s8765_7(wires_2191_6[1], addr_2191_6, addr_positional[35063:35060], addr_8765_7);

wire[31:0] addr_8766_7;

Selector_2 s8766_7(wires_2191_6[2], addr_2191_6, addr_positional[35067:35064], addr_8766_7);

wire[31:0] addr_8767_7;

Selector_2 s8767_7(wires_2191_6[3], addr_2191_6, addr_positional[35071:35068], addr_8767_7);

wire[31:0] addr_8768_7;

Selector_2 s8768_7(wires_2192_6[0], addr_2192_6, addr_positional[35075:35072], addr_8768_7);

wire[31:0] addr_8769_7;

Selector_2 s8769_7(wires_2192_6[1], addr_2192_6, addr_positional[35079:35076], addr_8769_7);

wire[31:0] addr_8770_7;

Selector_2 s8770_7(wires_2192_6[2], addr_2192_6, addr_positional[35083:35080], addr_8770_7);

wire[31:0] addr_8771_7;

Selector_2 s8771_7(wires_2192_6[3], addr_2192_6, addr_positional[35087:35084], addr_8771_7);

wire[31:0] addr_8772_7;

Selector_2 s8772_7(wires_2193_6[0], addr_2193_6, addr_positional[35091:35088], addr_8772_7);

wire[31:0] addr_8773_7;

Selector_2 s8773_7(wires_2193_6[1], addr_2193_6, addr_positional[35095:35092], addr_8773_7);

wire[31:0] addr_8774_7;

Selector_2 s8774_7(wires_2193_6[2], addr_2193_6, addr_positional[35099:35096], addr_8774_7);

wire[31:0] addr_8775_7;

Selector_2 s8775_7(wires_2193_6[3], addr_2193_6, addr_positional[35103:35100], addr_8775_7);

wire[31:0] addr_8776_7;

Selector_2 s8776_7(wires_2194_6[0], addr_2194_6, addr_positional[35107:35104], addr_8776_7);

wire[31:0] addr_8777_7;

Selector_2 s8777_7(wires_2194_6[1], addr_2194_6, addr_positional[35111:35108], addr_8777_7);

wire[31:0] addr_8778_7;

Selector_2 s8778_7(wires_2194_6[2], addr_2194_6, addr_positional[35115:35112], addr_8778_7);

wire[31:0] addr_8779_7;

Selector_2 s8779_7(wires_2194_6[3], addr_2194_6, addr_positional[35119:35116], addr_8779_7);

wire[31:0] addr_8780_7;

Selector_2 s8780_7(wires_2195_6[0], addr_2195_6, addr_positional[35123:35120], addr_8780_7);

wire[31:0] addr_8781_7;

Selector_2 s8781_7(wires_2195_6[1], addr_2195_6, addr_positional[35127:35124], addr_8781_7);

wire[31:0] addr_8782_7;

Selector_2 s8782_7(wires_2195_6[2], addr_2195_6, addr_positional[35131:35128], addr_8782_7);

wire[31:0] addr_8783_7;

Selector_2 s8783_7(wires_2195_6[3], addr_2195_6, addr_positional[35135:35132], addr_8783_7);

wire[31:0] addr_8784_7;

Selector_2 s8784_7(wires_2196_6[0], addr_2196_6, addr_positional[35139:35136], addr_8784_7);

wire[31:0] addr_8785_7;

Selector_2 s8785_7(wires_2196_6[1], addr_2196_6, addr_positional[35143:35140], addr_8785_7);

wire[31:0] addr_8786_7;

Selector_2 s8786_7(wires_2196_6[2], addr_2196_6, addr_positional[35147:35144], addr_8786_7);

wire[31:0] addr_8787_7;

Selector_2 s8787_7(wires_2196_6[3], addr_2196_6, addr_positional[35151:35148], addr_8787_7);

wire[31:0] addr_8788_7;

Selector_2 s8788_7(wires_2197_6[0], addr_2197_6, addr_positional[35155:35152], addr_8788_7);

wire[31:0] addr_8789_7;

Selector_2 s8789_7(wires_2197_6[1], addr_2197_6, addr_positional[35159:35156], addr_8789_7);

wire[31:0] addr_8790_7;

Selector_2 s8790_7(wires_2197_6[2], addr_2197_6, addr_positional[35163:35160], addr_8790_7);

wire[31:0] addr_8791_7;

Selector_2 s8791_7(wires_2197_6[3], addr_2197_6, addr_positional[35167:35164], addr_8791_7);

wire[31:0] addr_8792_7;

Selector_2 s8792_7(wires_2198_6[0], addr_2198_6, addr_positional[35171:35168], addr_8792_7);

wire[31:0] addr_8793_7;

Selector_2 s8793_7(wires_2198_6[1], addr_2198_6, addr_positional[35175:35172], addr_8793_7);

wire[31:0] addr_8794_7;

Selector_2 s8794_7(wires_2198_6[2], addr_2198_6, addr_positional[35179:35176], addr_8794_7);

wire[31:0] addr_8795_7;

Selector_2 s8795_7(wires_2198_6[3], addr_2198_6, addr_positional[35183:35180], addr_8795_7);

wire[31:0] addr_8796_7;

Selector_2 s8796_7(wires_2199_6[0], addr_2199_6, addr_positional[35187:35184], addr_8796_7);

wire[31:0] addr_8797_7;

Selector_2 s8797_7(wires_2199_6[1], addr_2199_6, addr_positional[35191:35188], addr_8797_7);

wire[31:0] addr_8798_7;

Selector_2 s8798_7(wires_2199_6[2], addr_2199_6, addr_positional[35195:35192], addr_8798_7);

wire[31:0] addr_8799_7;

Selector_2 s8799_7(wires_2199_6[3], addr_2199_6, addr_positional[35199:35196], addr_8799_7);

wire[31:0] addr_8800_7;

Selector_2 s8800_7(wires_2200_6[0], addr_2200_6, addr_positional[35203:35200], addr_8800_7);

wire[31:0] addr_8801_7;

Selector_2 s8801_7(wires_2200_6[1], addr_2200_6, addr_positional[35207:35204], addr_8801_7);

wire[31:0] addr_8802_7;

Selector_2 s8802_7(wires_2200_6[2], addr_2200_6, addr_positional[35211:35208], addr_8802_7);

wire[31:0] addr_8803_7;

Selector_2 s8803_7(wires_2200_6[3], addr_2200_6, addr_positional[35215:35212], addr_8803_7);

wire[31:0] addr_8804_7;

Selector_2 s8804_7(wires_2201_6[0], addr_2201_6, addr_positional[35219:35216], addr_8804_7);

wire[31:0] addr_8805_7;

Selector_2 s8805_7(wires_2201_6[1], addr_2201_6, addr_positional[35223:35220], addr_8805_7);

wire[31:0] addr_8806_7;

Selector_2 s8806_7(wires_2201_6[2], addr_2201_6, addr_positional[35227:35224], addr_8806_7);

wire[31:0] addr_8807_7;

Selector_2 s8807_7(wires_2201_6[3], addr_2201_6, addr_positional[35231:35228], addr_8807_7);

wire[31:0] addr_8808_7;

Selector_2 s8808_7(wires_2202_6[0], addr_2202_6, addr_positional[35235:35232], addr_8808_7);

wire[31:0] addr_8809_7;

Selector_2 s8809_7(wires_2202_6[1], addr_2202_6, addr_positional[35239:35236], addr_8809_7);

wire[31:0] addr_8810_7;

Selector_2 s8810_7(wires_2202_6[2], addr_2202_6, addr_positional[35243:35240], addr_8810_7);

wire[31:0] addr_8811_7;

Selector_2 s8811_7(wires_2202_6[3], addr_2202_6, addr_positional[35247:35244], addr_8811_7);

wire[31:0] addr_8812_7;

Selector_2 s8812_7(wires_2203_6[0], addr_2203_6, addr_positional[35251:35248], addr_8812_7);

wire[31:0] addr_8813_7;

Selector_2 s8813_7(wires_2203_6[1], addr_2203_6, addr_positional[35255:35252], addr_8813_7);

wire[31:0] addr_8814_7;

Selector_2 s8814_7(wires_2203_6[2], addr_2203_6, addr_positional[35259:35256], addr_8814_7);

wire[31:0] addr_8815_7;

Selector_2 s8815_7(wires_2203_6[3], addr_2203_6, addr_positional[35263:35260], addr_8815_7);

wire[31:0] addr_8816_7;

Selector_2 s8816_7(wires_2204_6[0], addr_2204_6, addr_positional[35267:35264], addr_8816_7);

wire[31:0] addr_8817_7;

Selector_2 s8817_7(wires_2204_6[1], addr_2204_6, addr_positional[35271:35268], addr_8817_7);

wire[31:0] addr_8818_7;

Selector_2 s8818_7(wires_2204_6[2], addr_2204_6, addr_positional[35275:35272], addr_8818_7);

wire[31:0] addr_8819_7;

Selector_2 s8819_7(wires_2204_6[3], addr_2204_6, addr_positional[35279:35276], addr_8819_7);

wire[31:0] addr_8820_7;

Selector_2 s8820_7(wires_2205_6[0], addr_2205_6, addr_positional[35283:35280], addr_8820_7);

wire[31:0] addr_8821_7;

Selector_2 s8821_7(wires_2205_6[1], addr_2205_6, addr_positional[35287:35284], addr_8821_7);

wire[31:0] addr_8822_7;

Selector_2 s8822_7(wires_2205_6[2], addr_2205_6, addr_positional[35291:35288], addr_8822_7);

wire[31:0] addr_8823_7;

Selector_2 s8823_7(wires_2205_6[3], addr_2205_6, addr_positional[35295:35292], addr_8823_7);

wire[31:0] addr_8824_7;

Selector_2 s8824_7(wires_2206_6[0], addr_2206_6, addr_positional[35299:35296], addr_8824_7);

wire[31:0] addr_8825_7;

Selector_2 s8825_7(wires_2206_6[1], addr_2206_6, addr_positional[35303:35300], addr_8825_7);

wire[31:0] addr_8826_7;

Selector_2 s8826_7(wires_2206_6[2], addr_2206_6, addr_positional[35307:35304], addr_8826_7);

wire[31:0] addr_8827_7;

Selector_2 s8827_7(wires_2206_6[3], addr_2206_6, addr_positional[35311:35308], addr_8827_7);

wire[31:0] addr_8828_7;

Selector_2 s8828_7(wires_2207_6[0], addr_2207_6, addr_positional[35315:35312], addr_8828_7);

wire[31:0] addr_8829_7;

Selector_2 s8829_7(wires_2207_6[1], addr_2207_6, addr_positional[35319:35316], addr_8829_7);

wire[31:0] addr_8830_7;

Selector_2 s8830_7(wires_2207_6[2], addr_2207_6, addr_positional[35323:35320], addr_8830_7);

wire[31:0] addr_8831_7;

Selector_2 s8831_7(wires_2207_6[3], addr_2207_6, addr_positional[35327:35324], addr_8831_7);

wire[31:0] addr_8832_7;

Selector_2 s8832_7(wires_2208_6[0], addr_2208_6, addr_positional[35331:35328], addr_8832_7);

wire[31:0] addr_8833_7;

Selector_2 s8833_7(wires_2208_6[1], addr_2208_6, addr_positional[35335:35332], addr_8833_7);

wire[31:0] addr_8834_7;

Selector_2 s8834_7(wires_2208_6[2], addr_2208_6, addr_positional[35339:35336], addr_8834_7);

wire[31:0] addr_8835_7;

Selector_2 s8835_7(wires_2208_6[3], addr_2208_6, addr_positional[35343:35340], addr_8835_7);

wire[31:0] addr_8836_7;

Selector_2 s8836_7(wires_2209_6[0], addr_2209_6, addr_positional[35347:35344], addr_8836_7);

wire[31:0] addr_8837_7;

Selector_2 s8837_7(wires_2209_6[1], addr_2209_6, addr_positional[35351:35348], addr_8837_7);

wire[31:0] addr_8838_7;

Selector_2 s8838_7(wires_2209_6[2], addr_2209_6, addr_positional[35355:35352], addr_8838_7);

wire[31:0] addr_8839_7;

Selector_2 s8839_7(wires_2209_6[3], addr_2209_6, addr_positional[35359:35356], addr_8839_7);

wire[31:0] addr_8840_7;

Selector_2 s8840_7(wires_2210_6[0], addr_2210_6, addr_positional[35363:35360], addr_8840_7);

wire[31:0] addr_8841_7;

Selector_2 s8841_7(wires_2210_6[1], addr_2210_6, addr_positional[35367:35364], addr_8841_7);

wire[31:0] addr_8842_7;

Selector_2 s8842_7(wires_2210_6[2], addr_2210_6, addr_positional[35371:35368], addr_8842_7);

wire[31:0] addr_8843_7;

Selector_2 s8843_7(wires_2210_6[3], addr_2210_6, addr_positional[35375:35372], addr_8843_7);

wire[31:0] addr_8844_7;

Selector_2 s8844_7(wires_2211_6[0], addr_2211_6, addr_positional[35379:35376], addr_8844_7);

wire[31:0] addr_8845_7;

Selector_2 s8845_7(wires_2211_6[1], addr_2211_6, addr_positional[35383:35380], addr_8845_7);

wire[31:0] addr_8846_7;

Selector_2 s8846_7(wires_2211_6[2], addr_2211_6, addr_positional[35387:35384], addr_8846_7);

wire[31:0] addr_8847_7;

Selector_2 s8847_7(wires_2211_6[3], addr_2211_6, addr_positional[35391:35388], addr_8847_7);

wire[31:0] addr_8848_7;

Selector_2 s8848_7(wires_2212_6[0], addr_2212_6, addr_positional[35395:35392], addr_8848_7);

wire[31:0] addr_8849_7;

Selector_2 s8849_7(wires_2212_6[1], addr_2212_6, addr_positional[35399:35396], addr_8849_7);

wire[31:0] addr_8850_7;

Selector_2 s8850_7(wires_2212_6[2], addr_2212_6, addr_positional[35403:35400], addr_8850_7);

wire[31:0] addr_8851_7;

Selector_2 s8851_7(wires_2212_6[3], addr_2212_6, addr_positional[35407:35404], addr_8851_7);

wire[31:0] addr_8852_7;

Selector_2 s8852_7(wires_2213_6[0], addr_2213_6, addr_positional[35411:35408], addr_8852_7);

wire[31:0] addr_8853_7;

Selector_2 s8853_7(wires_2213_6[1], addr_2213_6, addr_positional[35415:35412], addr_8853_7);

wire[31:0] addr_8854_7;

Selector_2 s8854_7(wires_2213_6[2], addr_2213_6, addr_positional[35419:35416], addr_8854_7);

wire[31:0] addr_8855_7;

Selector_2 s8855_7(wires_2213_6[3], addr_2213_6, addr_positional[35423:35420], addr_8855_7);

wire[31:0] addr_8856_7;

Selector_2 s8856_7(wires_2214_6[0], addr_2214_6, addr_positional[35427:35424], addr_8856_7);

wire[31:0] addr_8857_7;

Selector_2 s8857_7(wires_2214_6[1], addr_2214_6, addr_positional[35431:35428], addr_8857_7);

wire[31:0] addr_8858_7;

Selector_2 s8858_7(wires_2214_6[2], addr_2214_6, addr_positional[35435:35432], addr_8858_7);

wire[31:0] addr_8859_7;

Selector_2 s8859_7(wires_2214_6[3], addr_2214_6, addr_positional[35439:35436], addr_8859_7);

wire[31:0] addr_8860_7;

Selector_2 s8860_7(wires_2215_6[0], addr_2215_6, addr_positional[35443:35440], addr_8860_7);

wire[31:0] addr_8861_7;

Selector_2 s8861_7(wires_2215_6[1], addr_2215_6, addr_positional[35447:35444], addr_8861_7);

wire[31:0] addr_8862_7;

Selector_2 s8862_7(wires_2215_6[2], addr_2215_6, addr_positional[35451:35448], addr_8862_7);

wire[31:0] addr_8863_7;

Selector_2 s8863_7(wires_2215_6[3], addr_2215_6, addr_positional[35455:35452], addr_8863_7);

wire[31:0] addr_8864_7;

Selector_2 s8864_7(wires_2216_6[0], addr_2216_6, addr_positional[35459:35456], addr_8864_7);

wire[31:0] addr_8865_7;

Selector_2 s8865_7(wires_2216_6[1], addr_2216_6, addr_positional[35463:35460], addr_8865_7);

wire[31:0] addr_8866_7;

Selector_2 s8866_7(wires_2216_6[2], addr_2216_6, addr_positional[35467:35464], addr_8866_7);

wire[31:0] addr_8867_7;

Selector_2 s8867_7(wires_2216_6[3], addr_2216_6, addr_positional[35471:35468], addr_8867_7);

wire[31:0] addr_8868_7;

Selector_2 s8868_7(wires_2217_6[0], addr_2217_6, addr_positional[35475:35472], addr_8868_7);

wire[31:0] addr_8869_7;

Selector_2 s8869_7(wires_2217_6[1], addr_2217_6, addr_positional[35479:35476], addr_8869_7);

wire[31:0] addr_8870_7;

Selector_2 s8870_7(wires_2217_6[2], addr_2217_6, addr_positional[35483:35480], addr_8870_7);

wire[31:0] addr_8871_7;

Selector_2 s8871_7(wires_2217_6[3], addr_2217_6, addr_positional[35487:35484], addr_8871_7);

wire[31:0] addr_8872_7;

Selector_2 s8872_7(wires_2218_6[0], addr_2218_6, addr_positional[35491:35488], addr_8872_7);

wire[31:0] addr_8873_7;

Selector_2 s8873_7(wires_2218_6[1], addr_2218_6, addr_positional[35495:35492], addr_8873_7);

wire[31:0] addr_8874_7;

Selector_2 s8874_7(wires_2218_6[2], addr_2218_6, addr_positional[35499:35496], addr_8874_7);

wire[31:0] addr_8875_7;

Selector_2 s8875_7(wires_2218_6[3], addr_2218_6, addr_positional[35503:35500], addr_8875_7);

wire[31:0] addr_8876_7;

Selector_2 s8876_7(wires_2219_6[0], addr_2219_6, addr_positional[35507:35504], addr_8876_7);

wire[31:0] addr_8877_7;

Selector_2 s8877_7(wires_2219_6[1], addr_2219_6, addr_positional[35511:35508], addr_8877_7);

wire[31:0] addr_8878_7;

Selector_2 s8878_7(wires_2219_6[2], addr_2219_6, addr_positional[35515:35512], addr_8878_7);

wire[31:0] addr_8879_7;

Selector_2 s8879_7(wires_2219_6[3], addr_2219_6, addr_positional[35519:35516], addr_8879_7);

wire[31:0] addr_8880_7;

Selector_2 s8880_7(wires_2220_6[0], addr_2220_6, addr_positional[35523:35520], addr_8880_7);

wire[31:0] addr_8881_7;

Selector_2 s8881_7(wires_2220_6[1], addr_2220_6, addr_positional[35527:35524], addr_8881_7);

wire[31:0] addr_8882_7;

Selector_2 s8882_7(wires_2220_6[2], addr_2220_6, addr_positional[35531:35528], addr_8882_7);

wire[31:0] addr_8883_7;

Selector_2 s8883_7(wires_2220_6[3], addr_2220_6, addr_positional[35535:35532], addr_8883_7);

wire[31:0] addr_8884_7;

Selector_2 s8884_7(wires_2221_6[0], addr_2221_6, addr_positional[35539:35536], addr_8884_7);

wire[31:0] addr_8885_7;

Selector_2 s8885_7(wires_2221_6[1], addr_2221_6, addr_positional[35543:35540], addr_8885_7);

wire[31:0] addr_8886_7;

Selector_2 s8886_7(wires_2221_6[2], addr_2221_6, addr_positional[35547:35544], addr_8886_7);

wire[31:0] addr_8887_7;

Selector_2 s8887_7(wires_2221_6[3], addr_2221_6, addr_positional[35551:35548], addr_8887_7);

wire[31:0] addr_8888_7;

Selector_2 s8888_7(wires_2222_6[0], addr_2222_6, addr_positional[35555:35552], addr_8888_7);

wire[31:0] addr_8889_7;

Selector_2 s8889_7(wires_2222_6[1], addr_2222_6, addr_positional[35559:35556], addr_8889_7);

wire[31:0] addr_8890_7;

Selector_2 s8890_7(wires_2222_6[2], addr_2222_6, addr_positional[35563:35560], addr_8890_7);

wire[31:0] addr_8891_7;

Selector_2 s8891_7(wires_2222_6[3], addr_2222_6, addr_positional[35567:35564], addr_8891_7);

wire[31:0] addr_8892_7;

Selector_2 s8892_7(wires_2223_6[0], addr_2223_6, addr_positional[35571:35568], addr_8892_7);

wire[31:0] addr_8893_7;

Selector_2 s8893_7(wires_2223_6[1], addr_2223_6, addr_positional[35575:35572], addr_8893_7);

wire[31:0] addr_8894_7;

Selector_2 s8894_7(wires_2223_6[2], addr_2223_6, addr_positional[35579:35576], addr_8894_7);

wire[31:0] addr_8895_7;

Selector_2 s8895_7(wires_2223_6[3], addr_2223_6, addr_positional[35583:35580], addr_8895_7);

wire[31:0] addr_8896_7;

Selector_2 s8896_7(wires_2224_6[0], addr_2224_6, addr_positional[35587:35584], addr_8896_7);

wire[31:0] addr_8897_7;

Selector_2 s8897_7(wires_2224_6[1], addr_2224_6, addr_positional[35591:35588], addr_8897_7);

wire[31:0] addr_8898_7;

Selector_2 s8898_7(wires_2224_6[2], addr_2224_6, addr_positional[35595:35592], addr_8898_7);

wire[31:0] addr_8899_7;

Selector_2 s8899_7(wires_2224_6[3], addr_2224_6, addr_positional[35599:35596], addr_8899_7);

wire[31:0] addr_8900_7;

Selector_2 s8900_7(wires_2225_6[0], addr_2225_6, addr_positional[35603:35600], addr_8900_7);

wire[31:0] addr_8901_7;

Selector_2 s8901_7(wires_2225_6[1], addr_2225_6, addr_positional[35607:35604], addr_8901_7);

wire[31:0] addr_8902_7;

Selector_2 s8902_7(wires_2225_6[2], addr_2225_6, addr_positional[35611:35608], addr_8902_7);

wire[31:0] addr_8903_7;

Selector_2 s8903_7(wires_2225_6[3], addr_2225_6, addr_positional[35615:35612], addr_8903_7);

wire[31:0] addr_8904_7;

Selector_2 s8904_7(wires_2226_6[0], addr_2226_6, addr_positional[35619:35616], addr_8904_7);

wire[31:0] addr_8905_7;

Selector_2 s8905_7(wires_2226_6[1], addr_2226_6, addr_positional[35623:35620], addr_8905_7);

wire[31:0] addr_8906_7;

Selector_2 s8906_7(wires_2226_6[2], addr_2226_6, addr_positional[35627:35624], addr_8906_7);

wire[31:0] addr_8907_7;

Selector_2 s8907_7(wires_2226_6[3], addr_2226_6, addr_positional[35631:35628], addr_8907_7);

wire[31:0] addr_8908_7;

Selector_2 s8908_7(wires_2227_6[0], addr_2227_6, addr_positional[35635:35632], addr_8908_7);

wire[31:0] addr_8909_7;

Selector_2 s8909_7(wires_2227_6[1], addr_2227_6, addr_positional[35639:35636], addr_8909_7);

wire[31:0] addr_8910_7;

Selector_2 s8910_7(wires_2227_6[2], addr_2227_6, addr_positional[35643:35640], addr_8910_7);

wire[31:0] addr_8911_7;

Selector_2 s8911_7(wires_2227_6[3], addr_2227_6, addr_positional[35647:35644], addr_8911_7);

wire[31:0] addr_8912_7;

Selector_2 s8912_7(wires_2228_6[0], addr_2228_6, addr_positional[35651:35648], addr_8912_7);

wire[31:0] addr_8913_7;

Selector_2 s8913_7(wires_2228_6[1], addr_2228_6, addr_positional[35655:35652], addr_8913_7);

wire[31:0] addr_8914_7;

Selector_2 s8914_7(wires_2228_6[2], addr_2228_6, addr_positional[35659:35656], addr_8914_7);

wire[31:0] addr_8915_7;

Selector_2 s8915_7(wires_2228_6[3], addr_2228_6, addr_positional[35663:35660], addr_8915_7);

wire[31:0] addr_8916_7;

Selector_2 s8916_7(wires_2229_6[0], addr_2229_6, addr_positional[35667:35664], addr_8916_7);

wire[31:0] addr_8917_7;

Selector_2 s8917_7(wires_2229_6[1], addr_2229_6, addr_positional[35671:35668], addr_8917_7);

wire[31:0] addr_8918_7;

Selector_2 s8918_7(wires_2229_6[2], addr_2229_6, addr_positional[35675:35672], addr_8918_7);

wire[31:0] addr_8919_7;

Selector_2 s8919_7(wires_2229_6[3], addr_2229_6, addr_positional[35679:35676], addr_8919_7);

wire[31:0] addr_8920_7;

Selector_2 s8920_7(wires_2230_6[0], addr_2230_6, addr_positional[35683:35680], addr_8920_7);

wire[31:0] addr_8921_7;

Selector_2 s8921_7(wires_2230_6[1], addr_2230_6, addr_positional[35687:35684], addr_8921_7);

wire[31:0] addr_8922_7;

Selector_2 s8922_7(wires_2230_6[2], addr_2230_6, addr_positional[35691:35688], addr_8922_7);

wire[31:0] addr_8923_7;

Selector_2 s8923_7(wires_2230_6[3], addr_2230_6, addr_positional[35695:35692], addr_8923_7);

wire[31:0] addr_8924_7;

Selector_2 s8924_7(wires_2231_6[0], addr_2231_6, addr_positional[35699:35696], addr_8924_7);

wire[31:0] addr_8925_7;

Selector_2 s8925_7(wires_2231_6[1], addr_2231_6, addr_positional[35703:35700], addr_8925_7);

wire[31:0] addr_8926_7;

Selector_2 s8926_7(wires_2231_6[2], addr_2231_6, addr_positional[35707:35704], addr_8926_7);

wire[31:0] addr_8927_7;

Selector_2 s8927_7(wires_2231_6[3], addr_2231_6, addr_positional[35711:35708], addr_8927_7);

wire[31:0] addr_8928_7;

Selector_2 s8928_7(wires_2232_6[0], addr_2232_6, addr_positional[35715:35712], addr_8928_7);

wire[31:0] addr_8929_7;

Selector_2 s8929_7(wires_2232_6[1], addr_2232_6, addr_positional[35719:35716], addr_8929_7);

wire[31:0] addr_8930_7;

Selector_2 s8930_7(wires_2232_6[2], addr_2232_6, addr_positional[35723:35720], addr_8930_7);

wire[31:0] addr_8931_7;

Selector_2 s8931_7(wires_2232_6[3], addr_2232_6, addr_positional[35727:35724], addr_8931_7);

wire[31:0] addr_8932_7;

Selector_2 s8932_7(wires_2233_6[0], addr_2233_6, addr_positional[35731:35728], addr_8932_7);

wire[31:0] addr_8933_7;

Selector_2 s8933_7(wires_2233_6[1], addr_2233_6, addr_positional[35735:35732], addr_8933_7);

wire[31:0] addr_8934_7;

Selector_2 s8934_7(wires_2233_6[2], addr_2233_6, addr_positional[35739:35736], addr_8934_7);

wire[31:0] addr_8935_7;

Selector_2 s8935_7(wires_2233_6[3], addr_2233_6, addr_positional[35743:35740], addr_8935_7);

wire[31:0] addr_8936_7;

Selector_2 s8936_7(wires_2234_6[0], addr_2234_6, addr_positional[35747:35744], addr_8936_7);

wire[31:0] addr_8937_7;

Selector_2 s8937_7(wires_2234_6[1], addr_2234_6, addr_positional[35751:35748], addr_8937_7);

wire[31:0] addr_8938_7;

Selector_2 s8938_7(wires_2234_6[2], addr_2234_6, addr_positional[35755:35752], addr_8938_7);

wire[31:0] addr_8939_7;

Selector_2 s8939_7(wires_2234_6[3], addr_2234_6, addr_positional[35759:35756], addr_8939_7);

wire[31:0] addr_8940_7;

Selector_2 s8940_7(wires_2235_6[0], addr_2235_6, addr_positional[35763:35760], addr_8940_7);

wire[31:0] addr_8941_7;

Selector_2 s8941_7(wires_2235_6[1], addr_2235_6, addr_positional[35767:35764], addr_8941_7);

wire[31:0] addr_8942_7;

Selector_2 s8942_7(wires_2235_6[2], addr_2235_6, addr_positional[35771:35768], addr_8942_7);

wire[31:0] addr_8943_7;

Selector_2 s8943_7(wires_2235_6[3], addr_2235_6, addr_positional[35775:35772], addr_8943_7);

wire[31:0] addr_8944_7;

Selector_2 s8944_7(wires_2236_6[0], addr_2236_6, addr_positional[35779:35776], addr_8944_7);

wire[31:0] addr_8945_7;

Selector_2 s8945_7(wires_2236_6[1], addr_2236_6, addr_positional[35783:35780], addr_8945_7);

wire[31:0] addr_8946_7;

Selector_2 s8946_7(wires_2236_6[2], addr_2236_6, addr_positional[35787:35784], addr_8946_7);

wire[31:0] addr_8947_7;

Selector_2 s8947_7(wires_2236_6[3], addr_2236_6, addr_positional[35791:35788], addr_8947_7);

wire[31:0] addr_8948_7;

Selector_2 s8948_7(wires_2237_6[0], addr_2237_6, addr_positional[35795:35792], addr_8948_7);

wire[31:0] addr_8949_7;

Selector_2 s8949_7(wires_2237_6[1], addr_2237_6, addr_positional[35799:35796], addr_8949_7);

wire[31:0] addr_8950_7;

Selector_2 s8950_7(wires_2237_6[2], addr_2237_6, addr_positional[35803:35800], addr_8950_7);

wire[31:0] addr_8951_7;

Selector_2 s8951_7(wires_2237_6[3], addr_2237_6, addr_positional[35807:35804], addr_8951_7);

wire[31:0] addr_8952_7;

Selector_2 s8952_7(wires_2238_6[0], addr_2238_6, addr_positional[35811:35808], addr_8952_7);

wire[31:0] addr_8953_7;

Selector_2 s8953_7(wires_2238_6[1], addr_2238_6, addr_positional[35815:35812], addr_8953_7);

wire[31:0] addr_8954_7;

Selector_2 s8954_7(wires_2238_6[2], addr_2238_6, addr_positional[35819:35816], addr_8954_7);

wire[31:0] addr_8955_7;

Selector_2 s8955_7(wires_2238_6[3], addr_2238_6, addr_positional[35823:35820], addr_8955_7);

wire[31:0] addr_8956_7;

Selector_2 s8956_7(wires_2239_6[0], addr_2239_6, addr_positional[35827:35824], addr_8956_7);

wire[31:0] addr_8957_7;

Selector_2 s8957_7(wires_2239_6[1], addr_2239_6, addr_positional[35831:35828], addr_8957_7);

wire[31:0] addr_8958_7;

Selector_2 s8958_7(wires_2239_6[2], addr_2239_6, addr_positional[35835:35832], addr_8958_7);

wire[31:0] addr_8959_7;

Selector_2 s8959_7(wires_2239_6[3], addr_2239_6, addr_positional[35839:35836], addr_8959_7);

wire[31:0] addr_8960_7;

Selector_2 s8960_7(wires_2240_6[0], addr_2240_6, addr_positional[35843:35840], addr_8960_7);

wire[31:0] addr_8961_7;

Selector_2 s8961_7(wires_2240_6[1], addr_2240_6, addr_positional[35847:35844], addr_8961_7);

wire[31:0] addr_8962_7;

Selector_2 s8962_7(wires_2240_6[2], addr_2240_6, addr_positional[35851:35848], addr_8962_7);

wire[31:0] addr_8963_7;

Selector_2 s8963_7(wires_2240_6[3], addr_2240_6, addr_positional[35855:35852], addr_8963_7);

wire[31:0] addr_8964_7;

Selector_2 s8964_7(wires_2241_6[0], addr_2241_6, addr_positional[35859:35856], addr_8964_7);

wire[31:0] addr_8965_7;

Selector_2 s8965_7(wires_2241_6[1], addr_2241_6, addr_positional[35863:35860], addr_8965_7);

wire[31:0] addr_8966_7;

Selector_2 s8966_7(wires_2241_6[2], addr_2241_6, addr_positional[35867:35864], addr_8966_7);

wire[31:0] addr_8967_7;

Selector_2 s8967_7(wires_2241_6[3], addr_2241_6, addr_positional[35871:35868], addr_8967_7);

wire[31:0] addr_8968_7;

Selector_2 s8968_7(wires_2242_6[0], addr_2242_6, addr_positional[35875:35872], addr_8968_7);

wire[31:0] addr_8969_7;

Selector_2 s8969_7(wires_2242_6[1], addr_2242_6, addr_positional[35879:35876], addr_8969_7);

wire[31:0] addr_8970_7;

Selector_2 s8970_7(wires_2242_6[2], addr_2242_6, addr_positional[35883:35880], addr_8970_7);

wire[31:0] addr_8971_7;

Selector_2 s8971_7(wires_2242_6[3], addr_2242_6, addr_positional[35887:35884], addr_8971_7);

wire[31:0] addr_8972_7;

Selector_2 s8972_7(wires_2243_6[0], addr_2243_6, addr_positional[35891:35888], addr_8972_7);

wire[31:0] addr_8973_7;

Selector_2 s8973_7(wires_2243_6[1], addr_2243_6, addr_positional[35895:35892], addr_8973_7);

wire[31:0] addr_8974_7;

Selector_2 s8974_7(wires_2243_6[2], addr_2243_6, addr_positional[35899:35896], addr_8974_7);

wire[31:0] addr_8975_7;

Selector_2 s8975_7(wires_2243_6[3], addr_2243_6, addr_positional[35903:35900], addr_8975_7);

wire[31:0] addr_8976_7;

Selector_2 s8976_7(wires_2244_6[0], addr_2244_6, addr_positional[35907:35904], addr_8976_7);

wire[31:0] addr_8977_7;

Selector_2 s8977_7(wires_2244_6[1], addr_2244_6, addr_positional[35911:35908], addr_8977_7);

wire[31:0] addr_8978_7;

Selector_2 s8978_7(wires_2244_6[2], addr_2244_6, addr_positional[35915:35912], addr_8978_7);

wire[31:0] addr_8979_7;

Selector_2 s8979_7(wires_2244_6[3], addr_2244_6, addr_positional[35919:35916], addr_8979_7);

wire[31:0] addr_8980_7;

Selector_2 s8980_7(wires_2245_6[0], addr_2245_6, addr_positional[35923:35920], addr_8980_7);

wire[31:0] addr_8981_7;

Selector_2 s8981_7(wires_2245_6[1], addr_2245_6, addr_positional[35927:35924], addr_8981_7);

wire[31:0] addr_8982_7;

Selector_2 s8982_7(wires_2245_6[2], addr_2245_6, addr_positional[35931:35928], addr_8982_7);

wire[31:0] addr_8983_7;

Selector_2 s8983_7(wires_2245_6[3], addr_2245_6, addr_positional[35935:35932], addr_8983_7);

wire[31:0] addr_8984_7;

Selector_2 s8984_7(wires_2246_6[0], addr_2246_6, addr_positional[35939:35936], addr_8984_7);

wire[31:0] addr_8985_7;

Selector_2 s8985_7(wires_2246_6[1], addr_2246_6, addr_positional[35943:35940], addr_8985_7);

wire[31:0] addr_8986_7;

Selector_2 s8986_7(wires_2246_6[2], addr_2246_6, addr_positional[35947:35944], addr_8986_7);

wire[31:0] addr_8987_7;

Selector_2 s8987_7(wires_2246_6[3], addr_2246_6, addr_positional[35951:35948], addr_8987_7);

wire[31:0] addr_8988_7;

Selector_2 s8988_7(wires_2247_6[0], addr_2247_6, addr_positional[35955:35952], addr_8988_7);

wire[31:0] addr_8989_7;

Selector_2 s8989_7(wires_2247_6[1], addr_2247_6, addr_positional[35959:35956], addr_8989_7);

wire[31:0] addr_8990_7;

Selector_2 s8990_7(wires_2247_6[2], addr_2247_6, addr_positional[35963:35960], addr_8990_7);

wire[31:0] addr_8991_7;

Selector_2 s8991_7(wires_2247_6[3], addr_2247_6, addr_positional[35967:35964], addr_8991_7);

wire[31:0] addr_8992_7;

Selector_2 s8992_7(wires_2248_6[0], addr_2248_6, addr_positional[35971:35968], addr_8992_7);

wire[31:0] addr_8993_7;

Selector_2 s8993_7(wires_2248_6[1], addr_2248_6, addr_positional[35975:35972], addr_8993_7);

wire[31:0] addr_8994_7;

Selector_2 s8994_7(wires_2248_6[2], addr_2248_6, addr_positional[35979:35976], addr_8994_7);

wire[31:0] addr_8995_7;

Selector_2 s8995_7(wires_2248_6[3], addr_2248_6, addr_positional[35983:35980], addr_8995_7);

wire[31:0] addr_8996_7;

Selector_2 s8996_7(wires_2249_6[0], addr_2249_6, addr_positional[35987:35984], addr_8996_7);

wire[31:0] addr_8997_7;

Selector_2 s8997_7(wires_2249_6[1], addr_2249_6, addr_positional[35991:35988], addr_8997_7);

wire[31:0] addr_8998_7;

Selector_2 s8998_7(wires_2249_6[2], addr_2249_6, addr_positional[35995:35992], addr_8998_7);

wire[31:0] addr_8999_7;

Selector_2 s8999_7(wires_2249_6[3], addr_2249_6, addr_positional[35999:35996], addr_8999_7);

wire[31:0] addr_9000_7;

Selector_2 s9000_7(wires_2250_6[0], addr_2250_6, addr_positional[36003:36000], addr_9000_7);

wire[31:0] addr_9001_7;

Selector_2 s9001_7(wires_2250_6[1], addr_2250_6, addr_positional[36007:36004], addr_9001_7);

wire[31:0] addr_9002_7;

Selector_2 s9002_7(wires_2250_6[2], addr_2250_6, addr_positional[36011:36008], addr_9002_7);

wire[31:0] addr_9003_7;

Selector_2 s9003_7(wires_2250_6[3], addr_2250_6, addr_positional[36015:36012], addr_9003_7);

wire[31:0] addr_9004_7;

Selector_2 s9004_7(wires_2251_6[0], addr_2251_6, addr_positional[36019:36016], addr_9004_7);

wire[31:0] addr_9005_7;

Selector_2 s9005_7(wires_2251_6[1], addr_2251_6, addr_positional[36023:36020], addr_9005_7);

wire[31:0] addr_9006_7;

Selector_2 s9006_7(wires_2251_6[2], addr_2251_6, addr_positional[36027:36024], addr_9006_7);

wire[31:0] addr_9007_7;

Selector_2 s9007_7(wires_2251_6[3], addr_2251_6, addr_positional[36031:36028], addr_9007_7);

wire[31:0] addr_9008_7;

Selector_2 s9008_7(wires_2252_6[0], addr_2252_6, addr_positional[36035:36032], addr_9008_7);

wire[31:0] addr_9009_7;

Selector_2 s9009_7(wires_2252_6[1], addr_2252_6, addr_positional[36039:36036], addr_9009_7);

wire[31:0] addr_9010_7;

Selector_2 s9010_7(wires_2252_6[2], addr_2252_6, addr_positional[36043:36040], addr_9010_7);

wire[31:0] addr_9011_7;

Selector_2 s9011_7(wires_2252_6[3], addr_2252_6, addr_positional[36047:36044], addr_9011_7);

wire[31:0] addr_9012_7;

Selector_2 s9012_7(wires_2253_6[0], addr_2253_6, addr_positional[36051:36048], addr_9012_7);

wire[31:0] addr_9013_7;

Selector_2 s9013_7(wires_2253_6[1], addr_2253_6, addr_positional[36055:36052], addr_9013_7);

wire[31:0] addr_9014_7;

Selector_2 s9014_7(wires_2253_6[2], addr_2253_6, addr_positional[36059:36056], addr_9014_7);

wire[31:0] addr_9015_7;

Selector_2 s9015_7(wires_2253_6[3], addr_2253_6, addr_positional[36063:36060], addr_9015_7);

wire[31:0] addr_9016_7;

Selector_2 s9016_7(wires_2254_6[0], addr_2254_6, addr_positional[36067:36064], addr_9016_7);

wire[31:0] addr_9017_7;

Selector_2 s9017_7(wires_2254_6[1], addr_2254_6, addr_positional[36071:36068], addr_9017_7);

wire[31:0] addr_9018_7;

Selector_2 s9018_7(wires_2254_6[2], addr_2254_6, addr_positional[36075:36072], addr_9018_7);

wire[31:0] addr_9019_7;

Selector_2 s9019_7(wires_2254_6[3], addr_2254_6, addr_positional[36079:36076], addr_9019_7);

wire[31:0] addr_9020_7;

Selector_2 s9020_7(wires_2255_6[0], addr_2255_6, addr_positional[36083:36080], addr_9020_7);

wire[31:0] addr_9021_7;

Selector_2 s9021_7(wires_2255_6[1], addr_2255_6, addr_positional[36087:36084], addr_9021_7);

wire[31:0] addr_9022_7;

Selector_2 s9022_7(wires_2255_6[2], addr_2255_6, addr_positional[36091:36088], addr_9022_7);

wire[31:0] addr_9023_7;

Selector_2 s9023_7(wires_2255_6[3], addr_2255_6, addr_positional[36095:36092], addr_9023_7);

wire[31:0] addr_9024_7;

Selector_2 s9024_7(wires_2256_6[0], addr_2256_6, addr_positional[36099:36096], addr_9024_7);

wire[31:0] addr_9025_7;

Selector_2 s9025_7(wires_2256_6[1], addr_2256_6, addr_positional[36103:36100], addr_9025_7);

wire[31:0] addr_9026_7;

Selector_2 s9026_7(wires_2256_6[2], addr_2256_6, addr_positional[36107:36104], addr_9026_7);

wire[31:0] addr_9027_7;

Selector_2 s9027_7(wires_2256_6[3], addr_2256_6, addr_positional[36111:36108], addr_9027_7);

wire[31:0] addr_9028_7;

Selector_2 s9028_7(wires_2257_6[0], addr_2257_6, addr_positional[36115:36112], addr_9028_7);

wire[31:0] addr_9029_7;

Selector_2 s9029_7(wires_2257_6[1], addr_2257_6, addr_positional[36119:36116], addr_9029_7);

wire[31:0] addr_9030_7;

Selector_2 s9030_7(wires_2257_6[2], addr_2257_6, addr_positional[36123:36120], addr_9030_7);

wire[31:0] addr_9031_7;

Selector_2 s9031_7(wires_2257_6[3], addr_2257_6, addr_positional[36127:36124], addr_9031_7);

wire[31:0] addr_9032_7;

Selector_2 s9032_7(wires_2258_6[0], addr_2258_6, addr_positional[36131:36128], addr_9032_7);

wire[31:0] addr_9033_7;

Selector_2 s9033_7(wires_2258_6[1], addr_2258_6, addr_positional[36135:36132], addr_9033_7);

wire[31:0] addr_9034_7;

Selector_2 s9034_7(wires_2258_6[2], addr_2258_6, addr_positional[36139:36136], addr_9034_7);

wire[31:0] addr_9035_7;

Selector_2 s9035_7(wires_2258_6[3], addr_2258_6, addr_positional[36143:36140], addr_9035_7);

wire[31:0] addr_9036_7;

Selector_2 s9036_7(wires_2259_6[0], addr_2259_6, addr_positional[36147:36144], addr_9036_7);

wire[31:0] addr_9037_7;

Selector_2 s9037_7(wires_2259_6[1], addr_2259_6, addr_positional[36151:36148], addr_9037_7);

wire[31:0] addr_9038_7;

Selector_2 s9038_7(wires_2259_6[2], addr_2259_6, addr_positional[36155:36152], addr_9038_7);

wire[31:0] addr_9039_7;

Selector_2 s9039_7(wires_2259_6[3], addr_2259_6, addr_positional[36159:36156], addr_9039_7);

wire[31:0] addr_9040_7;

Selector_2 s9040_7(wires_2260_6[0], addr_2260_6, addr_positional[36163:36160], addr_9040_7);

wire[31:0] addr_9041_7;

Selector_2 s9041_7(wires_2260_6[1], addr_2260_6, addr_positional[36167:36164], addr_9041_7);

wire[31:0] addr_9042_7;

Selector_2 s9042_7(wires_2260_6[2], addr_2260_6, addr_positional[36171:36168], addr_9042_7);

wire[31:0] addr_9043_7;

Selector_2 s9043_7(wires_2260_6[3], addr_2260_6, addr_positional[36175:36172], addr_9043_7);

wire[31:0] addr_9044_7;

Selector_2 s9044_7(wires_2261_6[0], addr_2261_6, addr_positional[36179:36176], addr_9044_7);

wire[31:0] addr_9045_7;

Selector_2 s9045_7(wires_2261_6[1], addr_2261_6, addr_positional[36183:36180], addr_9045_7);

wire[31:0] addr_9046_7;

Selector_2 s9046_7(wires_2261_6[2], addr_2261_6, addr_positional[36187:36184], addr_9046_7);

wire[31:0] addr_9047_7;

Selector_2 s9047_7(wires_2261_6[3], addr_2261_6, addr_positional[36191:36188], addr_9047_7);

wire[31:0] addr_9048_7;

Selector_2 s9048_7(wires_2262_6[0], addr_2262_6, addr_positional[36195:36192], addr_9048_7);

wire[31:0] addr_9049_7;

Selector_2 s9049_7(wires_2262_6[1], addr_2262_6, addr_positional[36199:36196], addr_9049_7);

wire[31:0] addr_9050_7;

Selector_2 s9050_7(wires_2262_6[2], addr_2262_6, addr_positional[36203:36200], addr_9050_7);

wire[31:0] addr_9051_7;

Selector_2 s9051_7(wires_2262_6[3], addr_2262_6, addr_positional[36207:36204], addr_9051_7);

wire[31:0] addr_9052_7;

Selector_2 s9052_7(wires_2263_6[0], addr_2263_6, addr_positional[36211:36208], addr_9052_7);

wire[31:0] addr_9053_7;

Selector_2 s9053_7(wires_2263_6[1], addr_2263_6, addr_positional[36215:36212], addr_9053_7);

wire[31:0] addr_9054_7;

Selector_2 s9054_7(wires_2263_6[2], addr_2263_6, addr_positional[36219:36216], addr_9054_7);

wire[31:0] addr_9055_7;

Selector_2 s9055_7(wires_2263_6[3], addr_2263_6, addr_positional[36223:36220], addr_9055_7);

wire[31:0] addr_9056_7;

Selector_2 s9056_7(wires_2264_6[0], addr_2264_6, addr_positional[36227:36224], addr_9056_7);

wire[31:0] addr_9057_7;

Selector_2 s9057_7(wires_2264_6[1], addr_2264_6, addr_positional[36231:36228], addr_9057_7);

wire[31:0] addr_9058_7;

Selector_2 s9058_7(wires_2264_6[2], addr_2264_6, addr_positional[36235:36232], addr_9058_7);

wire[31:0] addr_9059_7;

Selector_2 s9059_7(wires_2264_6[3], addr_2264_6, addr_positional[36239:36236], addr_9059_7);

wire[31:0] addr_9060_7;

Selector_2 s9060_7(wires_2265_6[0], addr_2265_6, addr_positional[36243:36240], addr_9060_7);

wire[31:0] addr_9061_7;

Selector_2 s9061_7(wires_2265_6[1], addr_2265_6, addr_positional[36247:36244], addr_9061_7);

wire[31:0] addr_9062_7;

Selector_2 s9062_7(wires_2265_6[2], addr_2265_6, addr_positional[36251:36248], addr_9062_7);

wire[31:0] addr_9063_7;

Selector_2 s9063_7(wires_2265_6[3], addr_2265_6, addr_positional[36255:36252], addr_9063_7);

wire[31:0] addr_9064_7;

Selector_2 s9064_7(wires_2266_6[0], addr_2266_6, addr_positional[36259:36256], addr_9064_7);

wire[31:0] addr_9065_7;

Selector_2 s9065_7(wires_2266_6[1], addr_2266_6, addr_positional[36263:36260], addr_9065_7);

wire[31:0] addr_9066_7;

Selector_2 s9066_7(wires_2266_6[2], addr_2266_6, addr_positional[36267:36264], addr_9066_7);

wire[31:0] addr_9067_7;

Selector_2 s9067_7(wires_2266_6[3], addr_2266_6, addr_positional[36271:36268], addr_9067_7);

wire[31:0] addr_9068_7;

Selector_2 s9068_7(wires_2267_6[0], addr_2267_6, addr_positional[36275:36272], addr_9068_7);

wire[31:0] addr_9069_7;

Selector_2 s9069_7(wires_2267_6[1], addr_2267_6, addr_positional[36279:36276], addr_9069_7);

wire[31:0] addr_9070_7;

Selector_2 s9070_7(wires_2267_6[2], addr_2267_6, addr_positional[36283:36280], addr_9070_7);

wire[31:0] addr_9071_7;

Selector_2 s9071_7(wires_2267_6[3], addr_2267_6, addr_positional[36287:36284], addr_9071_7);

wire[31:0] addr_9072_7;

Selector_2 s9072_7(wires_2268_6[0], addr_2268_6, addr_positional[36291:36288], addr_9072_7);

wire[31:0] addr_9073_7;

Selector_2 s9073_7(wires_2268_6[1], addr_2268_6, addr_positional[36295:36292], addr_9073_7);

wire[31:0] addr_9074_7;

Selector_2 s9074_7(wires_2268_6[2], addr_2268_6, addr_positional[36299:36296], addr_9074_7);

wire[31:0] addr_9075_7;

Selector_2 s9075_7(wires_2268_6[3], addr_2268_6, addr_positional[36303:36300], addr_9075_7);

wire[31:0] addr_9076_7;

Selector_2 s9076_7(wires_2269_6[0], addr_2269_6, addr_positional[36307:36304], addr_9076_7);

wire[31:0] addr_9077_7;

Selector_2 s9077_7(wires_2269_6[1], addr_2269_6, addr_positional[36311:36308], addr_9077_7);

wire[31:0] addr_9078_7;

Selector_2 s9078_7(wires_2269_6[2], addr_2269_6, addr_positional[36315:36312], addr_9078_7);

wire[31:0] addr_9079_7;

Selector_2 s9079_7(wires_2269_6[3], addr_2269_6, addr_positional[36319:36316], addr_9079_7);

wire[31:0] addr_9080_7;

Selector_2 s9080_7(wires_2270_6[0], addr_2270_6, addr_positional[36323:36320], addr_9080_7);

wire[31:0] addr_9081_7;

Selector_2 s9081_7(wires_2270_6[1], addr_2270_6, addr_positional[36327:36324], addr_9081_7);

wire[31:0] addr_9082_7;

Selector_2 s9082_7(wires_2270_6[2], addr_2270_6, addr_positional[36331:36328], addr_9082_7);

wire[31:0] addr_9083_7;

Selector_2 s9083_7(wires_2270_6[3], addr_2270_6, addr_positional[36335:36332], addr_9083_7);

wire[31:0] addr_9084_7;

Selector_2 s9084_7(wires_2271_6[0], addr_2271_6, addr_positional[36339:36336], addr_9084_7);

wire[31:0] addr_9085_7;

Selector_2 s9085_7(wires_2271_6[1], addr_2271_6, addr_positional[36343:36340], addr_9085_7);

wire[31:0] addr_9086_7;

Selector_2 s9086_7(wires_2271_6[2], addr_2271_6, addr_positional[36347:36344], addr_9086_7);

wire[31:0] addr_9087_7;

Selector_2 s9087_7(wires_2271_6[3], addr_2271_6, addr_positional[36351:36348], addr_9087_7);

wire[31:0] addr_9088_7;

Selector_2 s9088_7(wires_2272_6[0], addr_2272_6, addr_positional[36355:36352], addr_9088_7);

wire[31:0] addr_9089_7;

Selector_2 s9089_7(wires_2272_6[1], addr_2272_6, addr_positional[36359:36356], addr_9089_7);

wire[31:0] addr_9090_7;

Selector_2 s9090_7(wires_2272_6[2], addr_2272_6, addr_positional[36363:36360], addr_9090_7);

wire[31:0] addr_9091_7;

Selector_2 s9091_7(wires_2272_6[3], addr_2272_6, addr_positional[36367:36364], addr_9091_7);

wire[31:0] addr_9092_7;

Selector_2 s9092_7(wires_2273_6[0], addr_2273_6, addr_positional[36371:36368], addr_9092_7);

wire[31:0] addr_9093_7;

Selector_2 s9093_7(wires_2273_6[1], addr_2273_6, addr_positional[36375:36372], addr_9093_7);

wire[31:0] addr_9094_7;

Selector_2 s9094_7(wires_2273_6[2], addr_2273_6, addr_positional[36379:36376], addr_9094_7);

wire[31:0] addr_9095_7;

Selector_2 s9095_7(wires_2273_6[3], addr_2273_6, addr_positional[36383:36380], addr_9095_7);

wire[31:0] addr_9096_7;

Selector_2 s9096_7(wires_2274_6[0], addr_2274_6, addr_positional[36387:36384], addr_9096_7);

wire[31:0] addr_9097_7;

Selector_2 s9097_7(wires_2274_6[1], addr_2274_6, addr_positional[36391:36388], addr_9097_7);

wire[31:0] addr_9098_7;

Selector_2 s9098_7(wires_2274_6[2], addr_2274_6, addr_positional[36395:36392], addr_9098_7);

wire[31:0] addr_9099_7;

Selector_2 s9099_7(wires_2274_6[3], addr_2274_6, addr_positional[36399:36396], addr_9099_7);

wire[31:0] addr_9100_7;

Selector_2 s9100_7(wires_2275_6[0], addr_2275_6, addr_positional[36403:36400], addr_9100_7);

wire[31:0] addr_9101_7;

Selector_2 s9101_7(wires_2275_6[1], addr_2275_6, addr_positional[36407:36404], addr_9101_7);

wire[31:0] addr_9102_7;

Selector_2 s9102_7(wires_2275_6[2], addr_2275_6, addr_positional[36411:36408], addr_9102_7);

wire[31:0] addr_9103_7;

Selector_2 s9103_7(wires_2275_6[3], addr_2275_6, addr_positional[36415:36412], addr_9103_7);

wire[31:0] addr_9104_7;

Selector_2 s9104_7(wires_2276_6[0], addr_2276_6, addr_positional[36419:36416], addr_9104_7);

wire[31:0] addr_9105_7;

Selector_2 s9105_7(wires_2276_6[1], addr_2276_6, addr_positional[36423:36420], addr_9105_7);

wire[31:0] addr_9106_7;

Selector_2 s9106_7(wires_2276_6[2], addr_2276_6, addr_positional[36427:36424], addr_9106_7);

wire[31:0] addr_9107_7;

Selector_2 s9107_7(wires_2276_6[3], addr_2276_6, addr_positional[36431:36428], addr_9107_7);

wire[31:0] addr_9108_7;

Selector_2 s9108_7(wires_2277_6[0], addr_2277_6, addr_positional[36435:36432], addr_9108_7);

wire[31:0] addr_9109_7;

Selector_2 s9109_7(wires_2277_6[1], addr_2277_6, addr_positional[36439:36436], addr_9109_7);

wire[31:0] addr_9110_7;

Selector_2 s9110_7(wires_2277_6[2], addr_2277_6, addr_positional[36443:36440], addr_9110_7);

wire[31:0] addr_9111_7;

Selector_2 s9111_7(wires_2277_6[3], addr_2277_6, addr_positional[36447:36444], addr_9111_7);

wire[31:0] addr_9112_7;

Selector_2 s9112_7(wires_2278_6[0], addr_2278_6, addr_positional[36451:36448], addr_9112_7);

wire[31:0] addr_9113_7;

Selector_2 s9113_7(wires_2278_6[1], addr_2278_6, addr_positional[36455:36452], addr_9113_7);

wire[31:0] addr_9114_7;

Selector_2 s9114_7(wires_2278_6[2], addr_2278_6, addr_positional[36459:36456], addr_9114_7);

wire[31:0] addr_9115_7;

Selector_2 s9115_7(wires_2278_6[3], addr_2278_6, addr_positional[36463:36460], addr_9115_7);

wire[31:0] addr_9116_7;

Selector_2 s9116_7(wires_2279_6[0], addr_2279_6, addr_positional[36467:36464], addr_9116_7);

wire[31:0] addr_9117_7;

Selector_2 s9117_7(wires_2279_6[1], addr_2279_6, addr_positional[36471:36468], addr_9117_7);

wire[31:0] addr_9118_7;

Selector_2 s9118_7(wires_2279_6[2], addr_2279_6, addr_positional[36475:36472], addr_9118_7);

wire[31:0] addr_9119_7;

Selector_2 s9119_7(wires_2279_6[3], addr_2279_6, addr_positional[36479:36476], addr_9119_7);

wire[31:0] addr_9120_7;

Selector_2 s9120_7(wires_2280_6[0], addr_2280_6, addr_positional[36483:36480], addr_9120_7);

wire[31:0] addr_9121_7;

Selector_2 s9121_7(wires_2280_6[1], addr_2280_6, addr_positional[36487:36484], addr_9121_7);

wire[31:0] addr_9122_7;

Selector_2 s9122_7(wires_2280_6[2], addr_2280_6, addr_positional[36491:36488], addr_9122_7);

wire[31:0] addr_9123_7;

Selector_2 s9123_7(wires_2280_6[3], addr_2280_6, addr_positional[36495:36492], addr_9123_7);

wire[31:0] addr_9124_7;

Selector_2 s9124_7(wires_2281_6[0], addr_2281_6, addr_positional[36499:36496], addr_9124_7);

wire[31:0] addr_9125_7;

Selector_2 s9125_7(wires_2281_6[1], addr_2281_6, addr_positional[36503:36500], addr_9125_7);

wire[31:0] addr_9126_7;

Selector_2 s9126_7(wires_2281_6[2], addr_2281_6, addr_positional[36507:36504], addr_9126_7);

wire[31:0] addr_9127_7;

Selector_2 s9127_7(wires_2281_6[3], addr_2281_6, addr_positional[36511:36508], addr_9127_7);

wire[31:0] addr_9128_7;

Selector_2 s9128_7(wires_2282_6[0], addr_2282_6, addr_positional[36515:36512], addr_9128_7);

wire[31:0] addr_9129_7;

Selector_2 s9129_7(wires_2282_6[1], addr_2282_6, addr_positional[36519:36516], addr_9129_7);

wire[31:0] addr_9130_7;

Selector_2 s9130_7(wires_2282_6[2], addr_2282_6, addr_positional[36523:36520], addr_9130_7);

wire[31:0] addr_9131_7;

Selector_2 s9131_7(wires_2282_6[3], addr_2282_6, addr_positional[36527:36524], addr_9131_7);

wire[31:0] addr_9132_7;

Selector_2 s9132_7(wires_2283_6[0], addr_2283_6, addr_positional[36531:36528], addr_9132_7);

wire[31:0] addr_9133_7;

Selector_2 s9133_7(wires_2283_6[1], addr_2283_6, addr_positional[36535:36532], addr_9133_7);

wire[31:0] addr_9134_7;

Selector_2 s9134_7(wires_2283_6[2], addr_2283_6, addr_positional[36539:36536], addr_9134_7);

wire[31:0] addr_9135_7;

Selector_2 s9135_7(wires_2283_6[3], addr_2283_6, addr_positional[36543:36540], addr_9135_7);

wire[31:0] addr_9136_7;

Selector_2 s9136_7(wires_2284_6[0], addr_2284_6, addr_positional[36547:36544], addr_9136_7);

wire[31:0] addr_9137_7;

Selector_2 s9137_7(wires_2284_6[1], addr_2284_6, addr_positional[36551:36548], addr_9137_7);

wire[31:0] addr_9138_7;

Selector_2 s9138_7(wires_2284_6[2], addr_2284_6, addr_positional[36555:36552], addr_9138_7);

wire[31:0] addr_9139_7;

Selector_2 s9139_7(wires_2284_6[3], addr_2284_6, addr_positional[36559:36556], addr_9139_7);

wire[31:0] addr_9140_7;

Selector_2 s9140_7(wires_2285_6[0], addr_2285_6, addr_positional[36563:36560], addr_9140_7);

wire[31:0] addr_9141_7;

Selector_2 s9141_7(wires_2285_6[1], addr_2285_6, addr_positional[36567:36564], addr_9141_7);

wire[31:0] addr_9142_7;

Selector_2 s9142_7(wires_2285_6[2], addr_2285_6, addr_positional[36571:36568], addr_9142_7);

wire[31:0] addr_9143_7;

Selector_2 s9143_7(wires_2285_6[3], addr_2285_6, addr_positional[36575:36572], addr_9143_7);

wire[31:0] addr_9144_7;

Selector_2 s9144_7(wires_2286_6[0], addr_2286_6, addr_positional[36579:36576], addr_9144_7);

wire[31:0] addr_9145_7;

Selector_2 s9145_7(wires_2286_6[1], addr_2286_6, addr_positional[36583:36580], addr_9145_7);

wire[31:0] addr_9146_7;

Selector_2 s9146_7(wires_2286_6[2], addr_2286_6, addr_positional[36587:36584], addr_9146_7);

wire[31:0] addr_9147_7;

Selector_2 s9147_7(wires_2286_6[3], addr_2286_6, addr_positional[36591:36588], addr_9147_7);

wire[31:0] addr_9148_7;

Selector_2 s9148_7(wires_2287_6[0], addr_2287_6, addr_positional[36595:36592], addr_9148_7);

wire[31:0] addr_9149_7;

Selector_2 s9149_7(wires_2287_6[1], addr_2287_6, addr_positional[36599:36596], addr_9149_7);

wire[31:0] addr_9150_7;

Selector_2 s9150_7(wires_2287_6[2], addr_2287_6, addr_positional[36603:36600], addr_9150_7);

wire[31:0] addr_9151_7;

Selector_2 s9151_7(wires_2287_6[3], addr_2287_6, addr_positional[36607:36604], addr_9151_7);

wire[31:0] addr_9152_7;

Selector_2 s9152_7(wires_2288_6[0], addr_2288_6, addr_positional[36611:36608], addr_9152_7);

wire[31:0] addr_9153_7;

Selector_2 s9153_7(wires_2288_6[1], addr_2288_6, addr_positional[36615:36612], addr_9153_7);

wire[31:0] addr_9154_7;

Selector_2 s9154_7(wires_2288_6[2], addr_2288_6, addr_positional[36619:36616], addr_9154_7);

wire[31:0] addr_9155_7;

Selector_2 s9155_7(wires_2288_6[3], addr_2288_6, addr_positional[36623:36620], addr_9155_7);

wire[31:0] addr_9156_7;

Selector_2 s9156_7(wires_2289_6[0], addr_2289_6, addr_positional[36627:36624], addr_9156_7);

wire[31:0] addr_9157_7;

Selector_2 s9157_7(wires_2289_6[1], addr_2289_6, addr_positional[36631:36628], addr_9157_7);

wire[31:0] addr_9158_7;

Selector_2 s9158_7(wires_2289_6[2], addr_2289_6, addr_positional[36635:36632], addr_9158_7);

wire[31:0] addr_9159_7;

Selector_2 s9159_7(wires_2289_6[3], addr_2289_6, addr_positional[36639:36636], addr_9159_7);

wire[31:0] addr_9160_7;

Selector_2 s9160_7(wires_2290_6[0], addr_2290_6, addr_positional[36643:36640], addr_9160_7);

wire[31:0] addr_9161_7;

Selector_2 s9161_7(wires_2290_6[1], addr_2290_6, addr_positional[36647:36644], addr_9161_7);

wire[31:0] addr_9162_7;

Selector_2 s9162_7(wires_2290_6[2], addr_2290_6, addr_positional[36651:36648], addr_9162_7);

wire[31:0] addr_9163_7;

Selector_2 s9163_7(wires_2290_6[3], addr_2290_6, addr_positional[36655:36652], addr_9163_7);

wire[31:0] addr_9164_7;

Selector_2 s9164_7(wires_2291_6[0], addr_2291_6, addr_positional[36659:36656], addr_9164_7);

wire[31:0] addr_9165_7;

Selector_2 s9165_7(wires_2291_6[1], addr_2291_6, addr_positional[36663:36660], addr_9165_7);

wire[31:0] addr_9166_7;

Selector_2 s9166_7(wires_2291_6[2], addr_2291_6, addr_positional[36667:36664], addr_9166_7);

wire[31:0] addr_9167_7;

Selector_2 s9167_7(wires_2291_6[3], addr_2291_6, addr_positional[36671:36668], addr_9167_7);

wire[31:0] addr_9168_7;

Selector_2 s9168_7(wires_2292_6[0], addr_2292_6, addr_positional[36675:36672], addr_9168_7);

wire[31:0] addr_9169_7;

Selector_2 s9169_7(wires_2292_6[1], addr_2292_6, addr_positional[36679:36676], addr_9169_7);

wire[31:0] addr_9170_7;

Selector_2 s9170_7(wires_2292_6[2], addr_2292_6, addr_positional[36683:36680], addr_9170_7);

wire[31:0] addr_9171_7;

Selector_2 s9171_7(wires_2292_6[3], addr_2292_6, addr_positional[36687:36684], addr_9171_7);

wire[31:0] addr_9172_7;

Selector_2 s9172_7(wires_2293_6[0], addr_2293_6, addr_positional[36691:36688], addr_9172_7);

wire[31:0] addr_9173_7;

Selector_2 s9173_7(wires_2293_6[1], addr_2293_6, addr_positional[36695:36692], addr_9173_7);

wire[31:0] addr_9174_7;

Selector_2 s9174_7(wires_2293_6[2], addr_2293_6, addr_positional[36699:36696], addr_9174_7);

wire[31:0] addr_9175_7;

Selector_2 s9175_7(wires_2293_6[3], addr_2293_6, addr_positional[36703:36700], addr_9175_7);

wire[31:0] addr_9176_7;

Selector_2 s9176_7(wires_2294_6[0], addr_2294_6, addr_positional[36707:36704], addr_9176_7);

wire[31:0] addr_9177_7;

Selector_2 s9177_7(wires_2294_6[1], addr_2294_6, addr_positional[36711:36708], addr_9177_7);

wire[31:0] addr_9178_7;

Selector_2 s9178_7(wires_2294_6[2], addr_2294_6, addr_positional[36715:36712], addr_9178_7);

wire[31:0] addr_9179_7;

Selector_2 s9179_7(wires_2294_6[3], addr_2294_6, addr_positional[36719:36716], addr_9179_7);

wire[31:0] addr_9180_7;

Selector_2 s9180_7(wires_2295_6[0], addr_2295_6, addr_positional[36723:36720], addr_9180_7);

wire[31:0] addr_9181_7;

Selector_2 s9181_7(wires_2295_6[1], addr_2295_6, addr_positional[36727:36724], addr_9181_7);

wire[31:0] addr_9182_7;

Selector_2 s9182_7(wires_2295_6[2], addr_2295_6, addr_positional[36731:36728], addr_9182_7);

wire[31:0] addr_9183_7;

Selector_2 s9183_7(wires_2295_6[3], addr_2295_6, addr_positional[36735:36732], addr_9183_7);

wire[31:0] addr_9184_7;

Selector_2 s9184_7(wires_2296_6[0], addr_2296_6, addr_positional[36739:36736], addr_9184_7);

wire[31:0] addr_9185_7;

Selector_2 s9185_7(wires_2296_6[1], addr_2296_6, addr_positional[36743:36740], addr_9185_7);

wire[31:0] addr_9186_7;

Selector_2 s9186_7(wires_2296_6[2], addr_2296_6, addr_positional[36747:36744], addr_9186_7);

wire[31:0] addr_9187_7;

Selector_2 s9187_7(wires_2296_6[3], addr_2296_6, addr_positional[36751:36748], addr_9187_7);

wire[31:0] addr_9188_7;

Selector_2 s9188_7(wires_2297_6[0], addr_2297_6, addr_positional[36755:36752], addr_9188_7);

wire[31:0] addr_9189_7;

Selector_2 s9189_7(wires_2297_6[1], addr_2297_6, addr_positional[36759:36756], addr_9189_7);

wire[31:0] addr_9190_7;

Selector_2 s9190_7(wires_2297_6[2], addr_2297_6, addr_positional[36763:36760], addr_9190_7);

wire[31:0] addr_9191_7;

Selector_2 s9191_7(wires_2297_6[3], addr_2297_6, addr_positional[36767:36764], addr_9191_7);

wire[31:0] addr_9192_7;

Selector_2 s9192_7(wires_2298_6[0], addr_2298_6, addr_positional[36771:36768], addr_9192_7);

wire[31:0] addr_9193_7;

Selector_2 s9193_7(wires_2298_6[1], addr_2298_6, addr_positional[36775:36772], addr_9193_7);

wire[31:0] addr_9194_7;

Selector_2 s9194_7(wires_2298_6[2], addr_2298_6, addr_positional[36779:36776], addr_9194_7);

wire[31:0] addr_9195_7;

Selector_2 s9195_7(wires_2298_6[3], addr_2298_6, addr_positional[36783:36780], addr_9195_7);

wire[31:0] addr_9196_7;

Selector_2 s9196_7(wires_2299_6[0], addr_2299_6, addr_positional[36787:36784], addr_9196_7);

wire[31:0] addr_9197_7;

Selector_2 s9197_7(wires_2299_6[1], addr_2299_6, addr_positional[36791:36788], addr_9197_7);

wire[31:0] addr_9198_7;

Selector_2 s9198_7(wires_2299_6[2], addr_2299_6, addr_positional[36795:36792], addr_9198_7);

wire[31:0] addr_9199_7;

Selector_2 s9199_7(wires_2299_6[3], addr_2299_6, addr_positional[36799:36796], addr_9199_7);

wire[31:0] addr_9200_7;

Selector_2 s9200_7(wires_2300_6[0], addr_2300_6, addr_positional[36803:36800], addr_9200_7);

wire[31:0] addr_9201_7;

Selector_2 s9201_7(wires_2300_6[1], addr_2300_6, addr_positional[36807:36804], addr_9201_7);

wire[31:0] addr_9202_7;

Selector_2 s9202_7(wires_2300_6[2], addr_2300_6, addr_positional[36811:36808], addr_9202_7);

wire[31:0] addr_9203_7;

Selector_2 s9203_7(wires_2300_6[3], addr_2300_6, addr_positional[36815:36812], addr_9203_7);

wire[31:0] addr_9204_7;

Selector_2 s9204_7(wires_2301_6[0], addr_2301_6, addr_positional[36819:36816], addr_9204_7);

wire[31:0] addr_9205_7;

Selector_2 s9205_7(wires_2301_6[1], addr_2301_6, addr_positional[36823:36820], addr_9205_7);

wire[31:0] addr_9206_7;

Selector_2 s9206_7(wires_2301_6[2], addr_2301_6, addr_positional[36827:36824], addr_9206_7);

wire[31:0] addr_9207_7;

Selector_2 s9207_7(wires_2301_6[3], addr_2301_6, addr_positional[36831:36828], addr_9207_7);

wire[31:0] addr_9208_7;

Selector_2 s9208_7(wires_2302_6[0], addr_2302_6, addr_positional[36835:36832], addr_9208_7);

wire[31:0] addr_9209_7;

Selector_2 s9209_7(wires_2302_6[1], addr_2302_6, addr_positional[36839:36836], addr_9209_7);

wire[31:0] addr_9210_7;

Selector_2 s9210_7(wires_2302_6[2], addr_2302_6, addr_positional[36843:36840], addr_9210_7);

wire[31:0] addr_9211_7;

Selector_2 s9211_7(wires_2302_6[3], addr_2302_6, addr_positional[36847:36844], addr_9211_7);

wire[31:0] addr_9212_7;

Selector_2 s9212_7(wires_2303_6[0], addr_2303_6, addr_positional[36851:36848], addr_9212_7);

wire[31:0] addr_9213_7;

Selector_2 s9213_7(wires_2303_6[1], addr_2303_6, addr_positional[36855:36852], addr_9213_7);

wire[31:0] addr_9214_7;

Selector_2 s9214_7(wires_2303_6[2], addr_2303_6, addr_positional[36859:36856], addr_9214_7);

wire[31:0] addr_9215_7;

Selector_2 s9215_7(wires_2303_6[3], addr_2303_6, addr_positional[36863:36860], addr_9215_7);

wire[31:0] addr_9216_7;

Selector_2 s9216_7(wires_2304_6[0], addr_2304_6, addr_positional[36867:36864], addr_9216_7);

wire[31:0] addr_9217_7;

Selector_2 s9217_7(wires_2304_6[1], addr_2304_6, addr_positional[36871:36868], addr_9217_7);

wire[31:0] addr_9218_7;

Selector_2 s9218_7(wires_2304_6[2], addr_2304_6, addr_positional[36875:36872], addr_9218_7);

wire[31:0] addr_9219_7;

Selector_2 s9219_7(wires_2304_6[3], addr_2304_6, addr_positional[36879:36876], addr_9219_7);

wire[31:0] addr_9220_7;

Selector_2 s9220_7(wires_2305_6[0], addr_2305_6, addr_positional[36883:36880], addr_9220_7);

wire[31:0] addr_9221_7;

Selector_2 s9221_7(wires_2305_6[1], addr_2305_6, addr_positional[36887:36884], addr_9221_7);

wire[31:0] addr_9222_7;

Selector_2 s9222_7(wires_2305_6[2], addr_2305_6, addr_positional[36891:36888], addr_9222_7);

wire[31:0] addr_9223_7;

Selector_2 s9223_7(wires_2305_6[3], addr_2305_6, addr_positional[36895:36892], addr_9223_7);

wire[31:0] addr_9224_7;

Selector_2 s9224_7(wires_2306_6[0], addr_2306_6, addr_positional[36899:36896], addr_9224_7);

wire[31:0] addr_9225_7;

Selector_2 s9225_7(wires_2306_6[1], addr_2306_6, addr_positional[36903:36900], addr_9225_7);

wire[31:0] addr_9226_7;

Selector_2 s9226_7(wires_2306_6[2], addr_2306_6, addr_positional[36907:36904], addr_9226_7);

wire[31:0] addr_9227_7;

Selector_2 s9227_7(wires_2306_6[3], addr_2306_6, addr_positional[36911:36908], addr_9227_7);

wire[31:0] addr_9228_7;

Selector_2 s9228_7(wires_2307_6[0], addr_2307_6, addr_positional[36915:36912], addr_9228_7);

wire[31:0] addr_9229_7;

Selector_2 s9229_7(wires_2307_6[1], addr_2307_6, addr_positional[36919:36916], addr_9229_7);

wire[31:0] addr_9230_7;

Selector_2 s9230_7(wires_2307_6[2], addr_2307_6, addr_positional[36923:36920], addr_9230_7);

wire[31:0] addr_9231_7;

Selector_2 s9231_7(wires_2307_6[3], addr_2307_6, addr_positional[36927:36924], addr_9231_7);

wire[31:0] addr_9232_7;

Selector_2 s9232_7(wires_2308_6[0], addr_2308_6, addr_positional[36931:36928], addr_9232_7);

wire[31:0] addr_9233_7;

Selector_2 s9233_7(wires_2308_6[1], addr_2308_6, addr_positional[36935:36932], addr_9233_7);

wire[31:0] addr_9234_7;

Selector_2 s9234_7(wires_2308_6[2], addr_2308_6, addr_positional[36939:36936], addr_9234_7);

wire[31:0] addr_9235_7;

Selector_2 s9235_7(wires_2308_6[3], addr_2308_6, addr_positional[36943:36940], addr_9235_7);

wire[31:0] addr_9236_7;

Selector_2 s9236_7(wires_2309_6[0], addr_2309_6, addr_positional[36947:36944], addr_9236_7);

wire[31:0] addr_9237_7;

Selector_2 s9237_7(wires_2309_6[1], addr_2309_6, addr_positional[36951:36948], addr_9237_7);

wire[31:0] addr_9238_7;

Selector_2 s9238_7(wires_2309_6[2], addr_2309_6, addr_positional[36955:36952], addr_9238_7);

wire[31:0] addr_9239_7;

Selector_2 s9239_7(wires_2309_6[3], addr_2309_6, addr_positional[36959:36956], addr_9239_7);

wire[31:0] addr_9240_7;

Selector_2 s9240_7(wires_2310_6[0], addr_2310_6, addr_positional[36963:36960], addr_9240_7);

wire[31:0] addr_9241_7;

Selector_2 s9241_7(wires_2310_6[1], addr_2310_6, addr_positional[36967:36964], addr_9241_7);

wire[31:0] addr_9242_7;

Selector_2 s9242_7(wires_2310_6[2], addr_2310_6, addr_positional[36971:36968], addr_9242_7);

wire[31:0] addr_9243_7;

Selector_2 s9243_7(wires_2310_6[3], addr_2310_6, addr_positional[36975:36972], addr_9243_7);

wire[31:0] addr_9244_7;

Selector_2 s9244_7(wires_2311_6[0], addr_2311_6, addr_positional[36979:36976], addr_9244_7);

wire[31:0] addr_9245_7;

Selector_2 s9245_7(wires_2311_6[1], addr_2311_6, addr_positional[36983:36980], addr_9245_7);

wire[31:0] addr_9246_7;

Selector_2 s9246_7(wires_2311_6[2], addr_2311_6, addr_positional[36987:36984], addr_9246_7);

wire[31:0] addr_9247_7;

Selector_2 s9247_7(wires_2311_6[3], addr_2311_6, addr_positional[36991:36988], addr_9247_7);

wire[31:0] addr_9248_7;

Selector_2 s9248_7(wires_2312_6[0], addr_2312_6, addr_positional[36995:36992], addr_9248_7);

wire[31:0] addr_9249_7;

Selector_2 s9249_7(wires_2312_6[1], addr_2312_6, addr_positional[36999:36996], addr_9249_7);

wire[31:0] addr_9250_7;

Selector_2 s9250_7(wires_2312_6[2], addr_2312_6, addr_positional[37003:37000], addr_9250_7);

wire[31:0] addr_9251_7;

Selector_2 s9251_7(wires_2312_6[3], addr_2312_6, addr_positional[37007:37004], addr_9251_7);

wire[31:0] addr_9252_7;

Selector_2 s9252_7(wires_2313_6[0], addr_2313_6, addr_positional[37011:37008], addr_9252_7);

wire[31:0] addr_9253_7;

Selector_2 s9253_7(wires_2313_6[1], addr_2313_6, addr_positional[37015:37012], addr_9253_7);

wire[31:0] addr_9254_7;

Selector_2 s9254_7(wires_2313_6[2], addr_2313_6, addr_positional[37019:37016], addr_9254_7);

wire[31:0] addr_9255_7;

Selector_2 s9255_7(wires_2313_6[3], addr_2313_6, addr_positional[37023:37020], addr_9255_7);

wire[31:0] addr_9256_7;

Selector_2 s9256_7(wires_2314_6[0], addr_2314_6, addr_positional[37027:37024], addr_9256_7);

wire[31:0] addr_9257_7;

Selector_2 s9257_7(wires_2314_6[1], addr_2314_6, addr_positional[37031:37028], addr_9257_7);

wire[31:0] addr_9258_7;

Selector_2 s9258_7(wires_2314_6[2], addr_2314_6, addr_positional[37035:37032], addr_9258_7);

wire[31:0] addr_9259_7;

Selector_2 s9259_7(wires_2314_6[3], addr_2314_6, addr_positional[37039:37036], addr_9259_7);

wire[31:0] addr_9260_7;

Selector_2 s9260_7(wires_2315_6[0], addr_2315_6, addr_positional[37043:37040], addr_9260_7);

wire[31:0] addr_9261_7;

Selector_2 s9261_7(wires_2315_6[1], addr_2315_6, addr_positional[37047:37044], addr_9261_7);

wire[31:0] addr_9262_7;

Selector_2 s9262_7(wires_2315_6[2], addr_2315_6, addr_positional[37051:37048], addr_9262_7);

wire[31:0] addr_9263_7;

Selector_2 s9263_7(wires_2315_6[3], addr_2315_6, addr_positional[37055:37052], addr_9263_7);

wire[31:0] addr_9264_7;

Selector_2 s9264_7(wires_2316_6[0], addr_2316_6, addr_positional[37059:37056], addr_9264_7);

wire[31:0] addr_9265_7;

Selector_2 s9265_7(wires_2316_6[1], addr_2316_6, addr_positional[37063:37060], addr_9265_7);

wire[31:0] addr_9266_7;

Selector_2 s9266_7(wires_2316_6[2], addr_2316_6, addr_positional[37067:37064], addr_9266_7);

wire[31:0] addr_9267_7;

Selector_2 s9267_7(wires_2316_6[3], addr_2316_6, addr_positional[37071:37068], addr_9267_7);

wire[31:0] addr_9268_7;

Selector_2 s9268_7(wires_2317_6[0], addr_2317_6, addr_positional[37075:37072], addr_9268_7);

wire[31:0] addr_9269_7;

Selector_2 s9269_7(wires_2317_6[1], addr_2317_6, addr_positional[37079:37076], addr_9269_7);

wire[31:0] addr_9270_7;

Selector_2 s9270_7(wires_2317_6[2], addr_2317_6, addr_positional[37083:37080], addr_9270_7);

wire[31:0] addr_9271_7;

Selector_2 s9271_7(wires_2317_6[3], addr_2317_6, addr_positional[37087:37084], addr_9271_7);

wire[31:0] addr_9272_7;

Selector_2 s9272_7(wires_2318_6[0], addr_2318_6, addr_positional[37091:37088], addr_9272_7);

wire[31:0] addr_9273_7;

Selector_2 s9273_7(wires_2318_6[1], addr_2318_6, addr_positional[37095:37092], addr_9273_7);

wire[31:0] addr_9274_7;

Selector_2 s9274_7(wires_2318_6[2], addr_2318_6, addr_positional[37099:37096], addr_9274_7);

wire[31:0] addr_9275_7;

Selector_2 s9275_7(wires_2318_6[3], addr_2318_6, addr_positional[37103:37100], addr_9275_7);

wire[31:0] addr_9276_7;

Selector_2 s9276_7(wires_2319_6[0], addr_2319_6, addr_positional[37107:37104], addr_9276_7);

wire[31:0] addr_9277_7;

Selector_2 s9277_7(wires_2319_6[1], addr_2319_6, addr_positional[37111:37108], addr_9277_7);

wire[31:0] addr_9278_7;

Selector_2 s9278_7(wires_2319_6[2], addr_2319_6, addr_positional[37115:37112], addr_9278_7);

wire[31:0] addr_9279_7;

Selector_2 s9279_7(wires_2319_6[3], addr_2319_6, addr_positional[37119:37116], addr_9279_7);

wire[31:0] addr_9280_7;

Selector_2 s9280_7(wires_2320_6[0], addr_2320_6, addr_positional[37123:37120], addr_9280_7);

wire[31:0] addr_9281_7;

Selector_2 s9281_7(wires_2320_6[1], addr_2320_6, addr_positional[37127:37124], addr_9281_7);

wire[31:0] addr_9282_7;

Selector_2 s9282_7(wires_2320_6[2], addr_2320_6, addr_positional[37131:37128], addr_9282_7);

wire[31:0] addr_9283_7;

Selector_2 s9283_7(wires_2320_6[3], addr_2320_6, addr_positional[37135:37132], addr_9283_7);

wire[31:0] addr_9284_7;

Selector_2 s9284_7(wires_2321_6[0], addr_2321_6, addr_positional[37139:37136], addr_9284_7);

wire[31:0] addr_9285_7;

Selector_2 s9285_7(wires_2321_6[1], addr_2321_6, addr_positional[37143:37140], addr_9285_7);

wire[31:0] addr_9286_7;

Selector_2 s9286_7(wires_2321_6[2], addr_2321_6, addr_positional[37147:37144], addr_9286_7);

wire[31:0] addr_9287_7;

Selector_2 s9287_7(wires_2321_6[3], addr_2321_6, addr_positional[37151:37148], addr_9287_7);

wire[31:0] addr_9288_7;

Selector_2 s9288_7(wires_2322_6[0], addr_2322_6, addr_positional[37155:37152], addr_9288_7);

wire[31:0] addr_9289_7;

Selector_2 s9289_7(wires_2322_6[1], addr_2322_6, addr_positional[37159:37156], addr_9289_7);

wire[31:0] addr_9290_7;

Selector_2 s9290_7(wires_2322_6[2], addr_2322_6, addr_positional[37163:37160], addr_9290_7);

wire[31:0] addr_9291_7;

Selector_2 s9291_7(wires_2322_6[3], addr_2322_6, addr_positional[37167:37164], addr_9291_7);

wire[31:0] addr_9292_7;

Selector_2 s9292_7(wires_2323_6[0], addr_2323_6, addr_positional[37171:37168], addr_9292_7);

wire[31:0] addr_9293_7;

Selector_2 s9293_7(wires_2323_6[1], addr_2323_6, addr_positional[37175:37172], addr_9293_7);

wire[31:0] addr_9294_7;

Selector_2 s9294_7(wires_2323_6[2], addr_2323_6, addr_positional[37179:37176], addr_9294_7);

wire[31:0] addr_9295_7;

Selector_2 s9295_7(wires_2323_6[3], addr_2323_6, addr_positional[37183:37180], addr_9295_7);

wire[31:0] addr_9296_7;

Selector_2 s9296_7(wires_2324_6[0], addr_2324_6, addr_positional[37187:37184], addr_9296_7);

wire[31:0] addr_9297_7;

Selector_2 s9297_7(wires_2324_6[1], addr_2324_6, addr_positional[37191:37188], addr_9297_7);

wire[31:0] addr_9298_7;

Selector_2 s9298_7(wires_2324_6[2], addr_2324_6, addr_positional[37195:37192], addr_9298_7);

wire[31:0] addr_9299_7;

Selector_2 s9299_7(wires_2324_6[3], addr_2324_6, addr_positional[37199:37196], addr_9299_7);

wire[31:0] addr_9300_7;

Selector_2 s9300_7(wires_2325_6[0], addr_2325_6, addr_positional[37203:37200], addr_9300_7);

wire[31:0] addr_9301_7;

Selector_2 s9301_7(wires_2325_6[1], addr_2325_6, addr_positional[37207:37204], addr_9301_7);

wire[31:0] addr_9302_7;

Selector_2 s9302_7(wires_2325_6[2], addr_2325_6, addr_positional[37211:37208], addr_9302_7);

wire[31:0] addr_9303_7;

Selector_2 s9303_7(wires_2325_6[3], addr_2325_6, addr_positional[37215:37212], addr_9303_7);

wire[31:0] addr_9304_7;

Selector_2 s9304_7(wires_2326_6[0], addr_2326_6, addr_positional[37219:37216], addr_9304_7);

wire[31:0] addr_9305_7;

Selector_2 s9305_7(wires_2326_6[1], addr_2326_6, addr_positional[37223:37220], addr_9305_7);

wire[31:0] addr_9306_7;

Selector_2 s9306_7(wires_2326_6[2], addr_2326_6, addr_positional[37227:37224], addr_9306_7);

wire[31:0] addr_9307_7;

Selector_2 s9307_7(wires_2326_6[3], addr_2326_6, addr_positional[37231:37228], addr_9307_7);

wire[31:0] addr_9308_7;

Selector_2 s9308_7(wires_2327_6[0], addr_2327_6, addr_positional[37235:37232], addr_9308_7);

wire[31:0] addr_9309_7;

Selector_2 s9309_7(wires_2327_6[1], addr_2327_6, addr_positional[37239:37236], addr_9309_7);

wire[31:0] addr_9310_7;

Selector_2 s9310_7(wires_2327_6[2], addr_2327_6, addr_positional[37243:37240], addr_9310_7);

wire[31:0] addr_9311_7;

Selector_2 s9311_7(wires_2327_6[3], addr_2327_6, addr_positional[37247:37244], addr_9311_7);

wire[31:0] addr_9312_7;

Selector_2 s9312_7(wires_2328_6[0], addr_2328_6, addr_positional[37251:37248], addr_9312_7);

wire[31:0] addr_9313_7;

Selector_2 s9313_7(wires_2328_6[1], addr_2328_6, addr_positional[37255:37252], addr_9313_7);

wire[31:0] addr_9314_7;

Selector_2 s9314_7(wires_2328_6[2], addr_2328_6, addr_positional[37259:37256], addr_9314_7);

wire[31:0] addr_9315_7;

Selector_2 s9315_7(wires_2328_6[3], addr_2328_6, addr_positional[37263:37260], addr_9315_7);

wire[31:0] addr_9316_7;

Selector_2 s9316_7(wires_2329_6[0], addr_2329_6, addr_positional[37267:37264], addr_9316_7);

wire[31:0] addr_9317_7;

Selector_2 s9317_7(wires_2329_6[1], addr_2329_6, addr_positional[37271:37268], addr_9317_7);

wire[31:0] addr_9318_7;

Selector_2 s9318_7(wires_2329_6[2], addr_2329_6, addr_positional[37275:37272], addr_9318_7);

wire[31:0] addr_9319_7;

Selector_2 s9319_7(wires_2329_6[3], addr_2329_6, addr_positional[37279:37276], addr_9319_7);

wire[31:0] addr_9320_7;

Selector_2 s9320_7(wires_2330_6[0], addr_2330_6, addr_positional[37283:37280], addr_9320_7);

wire[31:0] addr_9321_7;

Selector_2 s9321_7(wires_2330_6[1], addr_2330_6, addr_positional[37287:37284], addr_9321_7);

wire[31:0] addr_9322_7;

Selector_2 s9322_7(wires_2330_6[2], addr_2330_6, addr_positional[37291:37288], addr_9322_7);

wire[31:0] addr_9323_7;

Selector_2 s9323_7(wires_2330_6[3], addr_2330_6, addr_positional[37295:37292], addr_9323_7);

wire[31:0] addr_9324_7;

Selector_2 s9324_7(wires_2331_6[0], addr_2331_6, addr_positional[37299:37296], addr_9324_7);

wire[31:0] addr_9325_7;

Selector_2 s9325_7(wires_2331_6[1], addr_2331_6, addr_positional[37303:37300], addr_9325_7);

wire[31:0] addr_9326_7;

Selector_2 s9326_7(wires_2331_6[2], addr_2331_6, addr_positional[37307:37304], addr_9326_7);

wire[31:0] addr_9327_7;

Selector_2 s9327_7(wires_2331_6[3], addr_2331_6, addr_positional[37311:37308], addr_9327_7);

wire[31:0] addr_9328_7;

Selector_2 s9328_7(wires_2332_6[0], addr_2332_6, addr_positional[37315:37312], addr_9328_7);

wire[31:0] addr_9329_7;

Selector_2 s9329_7(wires_2332_6[1], addr_2332_6, addr_positional[37319:37316], addr_9329_7);

wire[31:0] addr_9330_7;

Selector_2 s9330_7(wires_2332_6[2], addr_2332_6, addr_positional[37323:37320], addr_9330_7);

wire[31:0] addr_9331_7;

Selector_2 s9331_7(wires_2332_6[3], addr_2332_6, addr_positional[37327:37324], addr_9331_7);

wire[31:0] addr_9332_7;

Selector_2 s9332_7(wires_2333_6[0], addr_2333_6, addr_positional[37331:37328], addr_9332_7);

wire[31:0] addr_9333_7;

Selector_2 s9333_7(wires_2333_6[1], addr_2333_6, addr_positional[37335:37332], addr_9333_7);

wire[31:0] addr_9334_7;

Selector_2 s9334_7(wires_2333_6[2], addr_2333_6, addr_positional[37339:37336], addr_9334_7);

wire[31:0] addr_9335_7;

Selector_2 s9335_7(wires_2333_6[3], addr_2333_6, addr_positional[37343:37340], addr_9335_7);

wire[31:0] addr_9336_7;

Selector_2 s9336_7(wires_2334_6[0], addr_2334_6, addr_positional[37347:37344], addr_9336_7);

wire[31:0] addr_9337_7;

Selector_2 s9337_7(wires_2334_6[1], addr_2334_6, addr_positional[37351:37348], addr_9337_7);

wire[31:0] addr_9338_7;

Selector_2 s9338_7(wires_2334_6[2], addr_2334_6, addr_positional[37355:37352], addr_9338_7);

wire[31:0] addr_9339_7;

Selector_2 s9339_7(wires_2334_6[3], addr_2334_6, addr_positional[37359:37356], addr_9339_7);

wire[31:0] addr_9340_7;

Selector_2 s9340_7(wires_2335_6[0], addr_2335_6, addr_positional[37363:37360], addr_9340_7);

wire[31:0] addr_9341_7;

Selector_2 s9341_7(wires_2335_6[1], addr_2335_6, addr_positional[37367:37364], addr_9341_7);

wire[31:0] addr_9342_7;

Selector_2 s9342_7(wires_2335_6[2], addr_2335_6, addr_positional[37371:37368], addr_9342_7);

wire[31:0] addr_9343_7;

Selector_2 s9343_7(wires_2335_6[3], addr_2335_6, addr_positional[37375:37372], addr_9343_7);

wire[31:0] addr_9344_7;

Selector_2 s9344_7(wires_2336_6[0], addr_2336_6, addr_positional[37379:37376], addr_9344_7);

wire[31:0] addr_9345_7;

Selector_2 s9345_7(wires_2336_6[1], addr_2336_6, addr_positional[37383:37380], addr_9345_7);

wire[31:0] addr_9346_7;

Selector_2 s9346_7(wires_2336_6[2], addr_2336_6, addr_positional[37387:37384], addr_9346_7);

wire[31:0] addr_9347_7;

Selector_2 s9347_7(wires_2336_6[3], addr_2336_6, addr_positional[37391:37388], addr_9347_7);

wire[31:0] addr_9348_7;

Selector_2 s9348_7(wires_2337_6[0], addr_2337_6, addr_positional[37395:37392], addr_9348_7);

wire[31:0] addr_9349_7;

Selector_2 s9349_7(wires_2337_6[1], addr_2337_6, addr_positional[37399:37396], addr_9349_7);

wire[31:0] addr_9350_7;

Selector_2 s9350_7(wires_2337_6[2], addr_2337_6, addr_positional[37403:37400], addr_9350_7);

wire[31:0] addr_9351_7;

Selector_2 s9351_7(wires_2337_6[3], addr_2337_6, addr_positional[37407:37404], addr_9351_7);

wire[31:0] addr_9352_7;

Selector_2 s9352_7(wires_2338_6[0], addr_2338_6, addr_positional[37411:37408], addr_9352_7);

wire[31:0] addr_9353_7;

Selector_2 s9353_7(wires_2338_6[1], addr_2338_6, addr_positional[37415:37412], addr_9353_7);

wire[31:0] addr_9354_7;

Selector_2 s9354_7(wires_2338_6[2], addr_2338_6, addr_positional[37419:37416], addr_9354_7);

wire[31:0] addr_9355_7;

Selector_2 s9355_7(wires_2338_6[3], addr_2338_6, addr_positional[37423:37420], addr_9355_7);

wire[31:0] addr_9356_7;

Selector_2 s9356_7(wires_2339_6[0], addr_2339_6, addr_positional[37427:37424], addr_9356_7);

wire[31:0] addr_9357_7;

Selector_2 s9357_7(wires_2339_6[1], addr_2339_6, addr_positional[37431:37428], addr_9357_7);

wire[31:0] addr_9358_7;

Selector_2 s9358_7(wires_2339_6[2], addr_2339_6, addr_positional[37435:37432], addr_9358_7);

wire[31:0] addr_9359_7;

Selector_2 s9359_7(wires_2339_6[3], addr_2339_6, addr_positional[37439:37436], addr_9359_7);

wire[31:0] addr_9360_7;

Selector_2 s9360_7(wires_2340_6[0], addr_2340_6, addr_positional[37443:37440], addr_9360_7);

wire[31:0] addr_9361_7;

Selector_2 s9361_7(wires_2340_6[1], addr_2340_6, addr_positional[37447:37444], addr_9361_7);

wire[31:0] addr_9362_7;

Selector_2 s9362_7(wires_2340_6[2], addr_2340_6, addr_positional[37451:37448], addr_9362_7);

wire[31:0] addr_9363_7;

Selector_2 s9363_7(wires_2340_6[3], addr_2340_6, addr_positional[37455:37452], addr_9363_7);

wire[31:0] addr_9364_7;

Selector_2 s9364_7(wires_2341_6[0], addr_2341_6, addr_positional[37459:37456], addr_9364_7);

wire[31:0] addr_9365_7;

Selector_2 s9365_7(wires_2341_6[1], addr_2341_6, addr_positional[37463:37460], addr_9365_7);

wire[31:0] addr_9366_7;

Selector_2 s9366_7(wires_2341_6[2], addr_2341_6, addr_positional[37467:37464], addr_9366_7);

wire[31:0] addr_9367_7;

Selector_2 s9367_7(wires_2341_6[3], addr_2341_6, addr_positional[37471:37468], addr_9367_7);

wire[31:0] addr_9368_7;

Selector_2 s9368_7(wires_2342_6[0], addr_2342_6, addr_positional[37475:37472], addr_9368_7);

wire[31:0] addr_9369_7;

Selector_2 s9369_7(wires_2342_6[1], addr_2342_6, addr_positional[37479:37476], addr_9369_7);

wire[31:0] addr_9370_7;

Selector_2 s9370_7(wires_2342_6[2], addr_2342_6, addr_positional[37483:37480], addr_9370_7);

wire[31:0] addr_9371_7;

Selector_2 s9371_7(wires_2342_6[3], addr_2342_6, addr_positional[37487:37484], addr_9371_7);

wire[31:0] addr_9372_7;

Selector_2 s9372_7(wires_2343_6[0], addr_2343_6, addr_positional[37491:37488], addr_9372_7);

wire[31:0] addr_9373_7;

Selector_2 s9373_7(wires_2343_6[1], addr_2343_6, addr_positional[37495:37492], addr_9373_7);

wire[31:0] addr_9374_7;

Selector_2 s9374_7(wires_2343_6[2], addr_2343_6, addr_positional[37499:37496], addr_9374_7);

wire[31:0] addr_9375_7;

Selector_2 s9375_7(wires_2343_6[3], addr_2343_6, addr_positional[37503:37500], addr_9375_7);

wire[31:0] addr_9376_7;

Selector_2 s9376_7(wires_2344_6[0], addr_2344_6, addr_positional[37507:37504], addr_9376_7);

wire[31:0] addr_9377_7;

Selector_2 s9377_7(wires_2344_6[1], addr_2344_6, addr_positional[37511:37508], addr_9377_7);

wire[31:0] addr_9378_7;

Selector_2 s9378_7(wires_2344_6[2], addr_2344_6, addr_positional[37515:37512], addr_9378_7);

wire[31:0] addr_9379_7;

Selector_2 s9379_7(wires_2344_6[3], addr_2344_6, addr_positional[37519:37516], addr_9379_7);

wire[31:0] addr_9380_7;

Selector_2 s9380_7(wires_2345_6[0], addr_2345_6, addr_positional[37523:37520], addr_9380_7);

wire[31:0] addr_9381_7;

Selector_2 s9381_7(wires_2345_6[1], addr_2345_6, addr_positional[37527:37524], addr_9381_7);

wire[31:0] addr_9382_7;

Selector_2 s9382_7(wires_2345_6[2], addr_2345_6, addr_positional[37531:37528], addr_9382_7);

wire[31:0] addr_9383_7;

Selector_2 s9383_7(wires_2345_6[3], addr_2345_6, addr_positional[37535:37532], addr_9383_7);

wire[31:0] addr_9384_7;

Selector_2 s9384_7(wires_2346_6[0], addr_2346_6, addr_positional[37539:37536], addr_9384_7);

wire[31:0] addr_9385_7;

Selector_2 s9385_7(wires_2346_6[1], addr_2346_6, addr_positional[37543:37540], addr_9385_7);

wire[31:0] addr_9386_7;

Selector_2 s9386_7(wires_2346_6[2], addr_2346_6, addr_positional[37547:37544], addr_9386_7);

wire[31:0] addr_9387_7;

Selector_2 s9387_7(wires_2346_6[3], addr_2346_6, addr_positional[37551:37548], addr_9387_7);

wire[31:0] addr_9388_7;

Selector_2 s9388_7(wires_2347_6[0], addr_2347_6, addr_positional[37555:37552], addr_9388_7);

wire[31:0] addr_9389_7;

Selector_2 s9389_7(wires_2347_6[1], addr_2347_6, addr_positional[37559:37556], addr_9389_7);

wire[31:0] addr_9390_7;

Selector_2 s9390_7(wires_2347_6[2], addr_2347_6, addr_positional[37563:37560], addr_9390_7);

wire[31:0] addr_9391_7;

Selector_2 s9391_7(wires_2347_6[3], addr_2347_6, addr_positional[37567:37564], addr_9391_7);

wire[31:0] addr_9392_7;

Selector_2 s9392_7(wires_2348_6[0], addr_2348_6, addr_positional[37571:37568], addr_9392_7);

wire[31:0] addr_9393_7;

Selector_2 s9393_7(wires_2348_6[1], addr_2348_6, addr_positional[37575:37572], addr_9393_7);

wire[31:0] addr_9394_7;

Selector_2 s9394_7(wires_2348_6[2], addr_2348_6, addr_positional[37579:37576], addr_9394_7);

wire[31:0] addr_9395_7;

Selector_2 s9395_7(wires_2348_6[3], addr_2348_6, addr_positional[37583:37580], addr_9395_7);

wire[31:0] addr_9396_7;

Selector_2 s9396_7(wires_2349_6[0], addr_2349_6, addr_positional[37587:37584], addr_9396_7);

wire[31:0] addr_9397_7;

Selector_2 s9397_7(wires_2349_6[1], addr_2349_6, addr_positional[37591:37588], addr_9397_7);

wire[31:0] addr_9398_7;

Selector_2 s9398_7(wires_2349_6[2], addr_2349_6, addr_positional[37595:37592], addr_9398_7);

wire[31:0] addr_9399_7;

Selector_2 s9399_7(wires_2349_6[3], addr_2349_6, addr_positional[37599:37596], addr_9399_7);

wire[31:0] addr_9400_7;

Selector_2 s9400_7(wires_2350_6[0], addr_2350_6, addr_positional[37603:37600], addr_9400_7);

wire[31:0] addr_9401_7;

Selector_2 s9401_7(wires_2350_6[1], addr_2350_6, addr_positional[37607:37604], addr_9401_7);

wire[31:0] addr_9402_7;

Selector_2 s9402_7(wires_2350_6[2], addr_2350_6, addr_positional[37611:37608], addr_9402_7);

wire[31:0] addr_9403_7;

Selector_2 s9403_7(wires_2350_6[3], addr_2350_6, addr_positional[37615:37612], addr_9403_7);

wire[31:0] addr_9404_7;

Selector_2 s9404_7(wires_2351_6[0], addr_2351_6, addr_positional[37619:37616], addr_9404_7);

wire[31:0] addr_9405_7;

Selector_2 s9405_7(wires_2351_6[1], addr_2351_6, addr_positional[37623:37620], addr_9405_7);

wire[31:0] addr_9406_7;

Selector_2 s9406_7(wires_2351_6[2], addr_2351_6, addr_positional[37627:37624], addr_9406_7);

wire[31:0] addr_9407_7;

Selector_2 s9407_7(wires_2351_6[3], addr_2351_6, addr_positional[37631:37628], addr_9407_7);

wire[31:0] addr_9408_7;

Selector_2 s9408_7(wires_2352_6[0], addr_2352_6, addr_positional[37635:37632], addr_9408_7);

wire[31:0] addr_9409_7;

Selector_2 s9409_7(wires_2352_6[1], addr_2352_6, addr_positional[37639:37636], addr_9409_7);

wire[31:0] addr_9410_7;

Selector_2 s9410_7(wires_2352_6[2], addr_2352_6, addr_positional[37643:37640], addr_9410_7);

wire[31:0] addr_9411_7;

Selector_2 s9411_7(wires_2352_6[3], addr_2352_6, addr_positional[37647:37644], addr_9411_7);

wire[31:0] addr_9412_7;

Selector_2 s9412_7(wires_2353_6[0], addr_2353_6, addr_positional[37651:37648], addr_9412_7);

wire[31:0] addr_9413_7;

Selector_2 s9413_7(wires_2353_6[1], addr_2353_6, addr_positional[37655:37652], addr_9413_7);

wire[31:0] addr_9414_7;

Selector_2 s9414_7(wires_2353_6[2], addr_2353_6, addr_positional[37659:37656], addr_9414_7);

wire[31:0] addr_9415_7;

Selector_2 s9415_7(wires_2353_6[3], addr_2353_6, addr_positional[37663:37660], addr_9415_7);

wire[31:0] addr_9416_7;

Selector_2 s9416_7(wires_2354_6[0], addr_2354_6, addr_positional[37667:37664], addr_9416_7);

wire[31:0] addr_9417_7;

Selector_2 s9417_7(wires_2354_6[1], addr_2354_6, addr_positional[37671:37668], addr_9417_7);

wire[31:0] addr_9418_7;

Selector_2 s9418_7(wires_2354_6[2], addr_2354_6, addr_positional[37675:37672], addr_9418_7);

wire[31:0] addr_9419_7;

Selector_2 s9419_7(wires_2354_6[3], addr_2354_6, addr_positional[37679:37676], addr_9419_7);

wire[31:0] addr_9420_7;

Selector_2 s9420_7(wires_2355_6[0], addr_2355_6, addr_positional[37683:37680], addr_9420_7);

wire[31:0] addr_9421_7;

Selector_2 s9421_7(wires_2355_6[1], addr_2355_6, addr_positional[37687:37684], addr_9421_7);

wire[31:0] addr_9422_7;

Selector_2 s9422_7(wires_2355_6[2], addr_2355_6, addr_positional[37691:37688], addr_9422_7);

wire[31:0] addr_9423_7;

Selector_2 s9423_7(wires_2355_6[3], addr_2355_6, addr_positional[37695:37692], addr_9423_7);

wire[31:0] addr_9424_7;

Selector_2 s9424_7(wires_2356_6[0], addr_2356_6, addr_positional[37699:37696], addr_9424_7);

wire[31:0] addr_9425_7;

Selector_2 s9425_7(wires_2356_6[1], addr_2356_6, addr_positional[37703:37700], addr_9425_7);

wire[31:0] addr_9426_7;

Selector_2 s9426_7(wires_2356_6[2], addr_2356_6, addr_positional[37707:37704], addr_9426_7);

wire[31:0] addr_9427_7;

Selector_2 s9427_7(wires_2356_6[3], addr_2356_6, addr_positional[37711:37708], addr_9427_7);

wire[31:0] addr_9428_7;

Selector_2 s9428_7(wires_2357_6[0], addr_2357_6, addr_positional[37715:37712], addr_9428_7);

wire[31:0] addr_9429_7;

Selector_2 s9429_7(wires_2357_6[1], addr_2357_6, addr_positional[37719:37716], addr_9429_7);

wire[31:0] addr_9430_7;

Selector_2 s9430_7(wires_2357_6[2], addr_2357_6, addr_positional[37723:37720], addr_9430_7);

wire[31:0] addr_9431_7;

Selector_2 s9431_7(wires_2357_6[3], addr_2357_6, addr_positional[37727:37724], addr_9431_7);

wire[31:0] addr_9432_7;

Selector_2 s9432_7(wires_2358_6[0], addr_2358_6, addr_positional[37731:37728], addr_9432_7);

wire[31:0] addr_9433_7;

Selector_2 s9433_7(wires_2358_6[1], addr_2358_6, addr_positional[37735:37732], addr_9433_7);

wire[31:0] addr_9434_7;

Selector_2 s9434_7(wires_2358_6[2], addr_2358_6, addr_positional[37739:37736], addr_9434_7);

wire[31:0] addr_9435_7;

Selector_2 s9435_7(wires_2358_6[3], addr_2358_6, addr_positional[37743:37740], addr_9435_7);

wire[31:0] addr_9436_7;

Selector_2 s9436_7(wires_2359_6[0], addr_2359_6, addr_positional[37747:37744], addr_9436_7);

wire[31:0] addr_9437_7;

Selector_2 s9437_7(wires_2359_6[1], addr_2359_6, addr_positional[37751:37748], addr_9437_7);

wire[31:0] addr_9438_7;

Selector_2 s9438_7(wires_2359_6[2], addr_2359_6, addr_positional[37755:37752], addr_9438_7);

wire[31:0] addr_9439_7;

Selector_2 s9439_7(wires_2359_6[3], addr_2359_6, addr_positional[37759:37756], addr_9439_7);

wire[31:0] addr_9440_7;

Selector_2 s9440_7(wires_2360_6[0], addr_2360_6, addr_positional[37763:37760], addr_9440_7);

wire[31:0] addr_9441_7;

Selector_2 s9441_7(wires_2360_6[1], addr_2360_6, addr_positional[37767:37764], addr_9441_7);

wire[31:0] addr_9442_7;

Selector_2 s9442_7(wires_2360_6[2], addr_2360_6, addr_positional[37771:37768], addr_9442_7);

wire[31:0] addr_9443_7;

Selector_2 s9443_7(wires_2360_6[3], addr_2360_6, addr_positional[37775:37772], addr_9443_7);

wire[31:0] addr_9444_7;

Selector_2 s9444_7(wires_2361_6[0], addr_2361_6, addr_positional[37779:37776], addr_9444_7);

wire[31:0] addr_9445_7;

Selector_2 s9445_7(wires_2361_6[1], addr_2361_6, addr_positional[37783:37780], addr_9445_7);

wire[31:0] addr_9446_7;

Selector_2 s9446_7(wires_2361_6[2], addr_2361_6, addr_positional[37787:37784], addr_9446_7);

wire[31:0] addr_9447_7;

Selector_2 s9447_7(wires_2361_6[3], addr_2361_6, addr_positional[37791:37788], addr_9447_7);

wire[31:0] addr_9448_7;

Selector_2 s9448_7(wires_2362_6[0], addr_2362_6, addr_positional[37795:37792], addr_9448_7);

wire[31:0] addr_9449_7;

Selector_2 s9449_7(wires_2362_6[1], addr_2362_6, addr_positional[37799:37796], addr_9449_7);

wire[31:0] addr_9450_7;

Selector_2 s9450_7(wires_2362_6[2], addr_2362_6, addr_positional[37803:37800], addr_9450_7);

wire[31:0] addr_9451_7;

Selector_2 s9451_7(wires_2362_6[3], addr_2362_6, addr_positional[37807:37804], addr_9451_7);

wire[31:0] addr_9452_7;

Selector_2 s9452_7(wires_2363_6[0], addr_2363_6, addr_positional[37811:37808], addr_9452_7);

wire[31:0] addr_9453_7;

Selector_2 s9453_7(wires_2363_6[1], addr_2363_6, addr_positional[37815:37812], addr_9453_7);

wire[31:0] addr_9454_7;

Selector_2 s9454_7(wires_2363_6[2], addr_2363_6, addr_positional[37819:37816], addr_9454_7);

wire[31:0] addr_9455_7;

Selector_2 s9455_7(wires_2363_6[3], addr_2363_6, addr_positional[37823:37820], addr_9455_7);

wire[31:0] addr_9456_7;

Selector_2 s9456_7(wires_2364_6[0], addr_2364_6, addr_positional[37827:37824], addr_9456_7);

wire[31:0] addr_9457_7;

Selector_2 s9457_7(wires_2364_6[1], addr_2364_6, addr_positional[37831:37828], addr_9457_7);

wire[31:0] addr_9458_7;

Selector_2 s9458_7(wires_2364_6[2], addr_2364_6, addr_positional[37835:37832], addr_9458_7);

wire[31:0] addr_9459_7;

Selector_2 s9459_7(wires_2364_6[3], addr_2364_6, addr_positional[37839:37836], addr_9459_7);

wire[31:0] addr_9460_7;

Selector_2 s9460_7(wires_2365_6[0], addr_2365_6, addr_positional[37843:37840], addr_9460_7);

wire[31:0] addr_9461_7;

Selector_2 s9461_7(wires_2365_6[1], addr_2365_6, addr_positional[37847:37844], addr_9461_7);

wire[31:0] addr_9462_7;

Selector_2 s9462_7(wires_2365_6[2], addr_2365_6, addr_positional[37851:37848], addr_9462_7);

wire[31:0] addr_9463_7;

Selector_2 s9463_7(wires_2365_6[3], addr_2365_6, addr_positional[37855:37852], addr_9463_7);

wire[31:0] addr_9464_7;

Selector_2 s9464_7(wires_2366_6[0], addr_2366_6, addr_positional[37859:37856], addr_9464_7);

wire[31:0] addr_9465_7;

Selector_2 s9465_7(wires_2366_6[1], addr_2366_6, addr_positional[37863:37860], addr_9465_7);

wire[31:0] addr_9466_7;

Selector_2 s9466_7(wires_2366_6[2], addr_2366_6, addr_positional[37867:37864], addr_9466_7);

wire[31:0] addr_9467_7;

Selector_2 s9467_7(wires_2366_6[3], addr_2366_6, addr_positional[37871:37868], addr_9467_7);

wire[31:0] addr_9468_7;

Selector_2 s9468_7(wires_2367_6[0], addr_2367_6, addr_positional[37875:37872], addr_9468_7);

wire[31:0] addr_9469_7;

Selector_2 s9469_7(wires_2367_6[1], addr_2367_6, addr_positional[37879:37876], addr_9469_7);

wire[31:0] addr_9470_7;

Selector_2 s9470_7(wires_2367_6[2], addr_2367_6, addr_positional[37883:37880], addr_9470_7);

wire[31:0] addr_9471_7;

Selector_2 s9471_7(wires_2367_6[3], addr_2367_6, addr_positional[37887:37884], addr_9471_7);

wire[31:0] addr_9472_7;

Selector_2 s9472_7(wires_2368_6[0], addr_2368_6, addr_positional[37891:37888], addr_9472_7);

wire[31:0] addr_9473_7;

Selector_2 s9473_7(wires_2368_6[1], addr_2368_6, addr_positional[37895:37892], addr_9473_7);

wire[31:0] addr_9474_7;

Selector_2 s9474_7(wires_2368_6[2], addr_2368_6, addr_positional[37899:37896], addr_9474_7);

wire[31:0] addr_9475_7;

Selector_2 s9475_7(wires_2368_6[3], addr_2368_6, addr_positional[37903:37900], addr_9475_7);

wire[31:0] addr_9476_7;

Selector_2 s9476_7(wires_2369_6[0], addr_2369_6, addr_positional[37907:37904], addr_9476_7);

wire[31:0] addr_9477_7;

Selector_2 s9477_7(wires_2369_6[1], addr_2369_6, addr_positional[37911:37908], addr_9477_7);

wire[31:0] addr_9478_7;

Selector_2 s9478_7(wires_2369_6[2], addr_2369_6, addr_positional[37915:37912], addr_9478_7);

wire[31:0] addr_9479_7;

Selector_2 s9479_7(wires_2369_6[3], addr_2369_6, addr_positional[37919:37916], addr_9479_7);

wire[31:0] addr_9480_7;

Selector_2 s9480_7(wires_2370_6[0], addr_2370_6, addr_positional[37923:37920], addr_9480_7);

wire[31:0] addr_9481_7;

Selector_2 s9481_7(wires_2370_6[1], addr_2370_6, addr_positional[37927:37924], addr_9481_7);

wire[31:0] addr_9482_7;

Selector_2 s9482_7(wires_2370_6[2], addr_2370_6, addr_positional[37931:37928], addr_9482_7);

wire[31:0] addr_9483_7;

Selector_2 s9483_7(wires_2370_6[3], addr_2370_6, addr_positional[37935:37932], addr_9483_7);

wire[31:0] addr_9484_7;

Selector_2 s9484_7(wires_2371_6[0], addr_2371_6, addr_positional[37939:37936], addr_9484_7);

wire[31:0] addr_9485_7;

Selector_2 s9485_7(wires_2371_6[1], addr_2371_6, addr_positional[37943:37940], addr_9485_7);

wire[31:0] addr_9486_7;

Selector_2 s9486_7(wires_2371_6[2], addr_2371_6, addr_positional[37947:37944], addr_9486_7);

wire[31:0] addr_9487_7;

Selector_2 s9487_7(wires_2371_6[3], addr_2371_6, addr_positional[37951:37948], addr_9487_7);

wire[31:0] addr_9488_7;

Selector_2 s9488_7(wires_2372_6[0], addr_2372_6, addr_positional[37955:37952], addr_9488_7);

wire[31:0] addr_9489_7;

Selector_2 s9489_7(wires_2372_6[1], addr_2372_6, addr_positional[37959:37956], addr_9489_7);

wire[31:0] addr_9490_7;

Selector_2 s9490_7(wires_2372_6[2], addr_2372_6, addr_positional[37963:37960], addr_9490_7);

wire[31:0] addr_9491_7;

Selector_2 s9491_7(wires_2372_6[3], addr_2372_6, addr_positional[37967:37964], addr_9491_7);

wire[31:0] addr_9492_7;

Selector_2 s9492_7(wires_2373_6[0], addr_2373_6, addr_positional[37971:37968], addr_9492_7);

wire[31:0] addr_9493_7;

Selector_2 s9493_7(wires_2373_6[1], addr_2373_6, addr_positional[37975:37972], addr_9493_7);

wire[31:0] addr_9494_7;

Selector_2 s9494_7(wires_2373_6[2], addr_2373_6, addr_positional[37979:37976], addr_9494_7);

wire[31:0] addr_9495_7;

Selector_2 s9495_7(wires_2373_6[3], addr_2373_6, addr_positional[37983:37980], addr_9495_7);

wire[31:0] addr_9496_7;

Selector_2 s9496_7(wires_2374_6[0], addr_2374_6, addr_positional[37987:37984], addr_9496_7);

wire[31:0] addr_9497_7;

Selector_2 s9497_7(wires_2374_6[1], addr_2374_6, addr_positional[37991:37988], addr_9497_7);

wire[31:0] addr_9498_7;

Selector_2 s9498_7(wires_2374_6[2], addr_2374_6, addr_positional[37995:37992], addr_9498_7);

wire[31:0] addr_9499_7;

Selector_2 s9499_7(wires_2374_6[3], addr_2374_6, addr_positional[37999:37996], addr_9499_7);

wire[31:0] addr_9500_7;

Selector_2 s9500_7(wires_2375_6[0], addr_2375_6, addr_positional[38003:38000], addr_9500_7);

wire[31:0] addr_9501_7;

Selector_2 s9501_7(wires_2375_6[1], addr_2375_6, addr_positional[38007:38004], addr_9501_7);

wire[31:0] addr_9502_7;

Selector_2 s9502_7(wires_2375_6[2], addr_2375_6, addr_positional[38011:38008], addr_9502_7);

wire[31:0] addr_9503_7;

Selector_2 s9503_7(wires_2375_6[3], addr_2375_6, addr_positional[38015:38012], addr_9503_7);

wire[31:0] addr_9504_7;

Selector_2 s9504_7(wires_2376_6[0], addr_2376_6, addr_positional[38019:38016], addr_9504_7);

wire[31:0] addr_9505_7;

Selector_2 s9505_7(wires_2376_6[1], addr_2376_6, addr_positional[38023:38020], addr_9505_7);

wire[31:0] addr_9506_7;

Selector_2 s9506_7(wires_2376_6[2], addr_2376_6, addr_positional[38027:38024], addr_9506_7);

wire[31:0] addr_9507_7;

Selector_2 s9507_7(wires_2376_6[3], addr_2376_6, addr_positional[38031:38028], addr_9507_7);

wire[31:0] addr_9508_7;

Selector_2 s9508_7(wires_2377_6[0], addr_2377_6, addr_positional[38035:38032], addr_9508_7);

wire[31:0] addr_9509_7;

Selector_2 s9509_7(wires_2377_6[1], addr_2377_6, addr_positional[38039:38036], addr_9509_7);

wire[31:0] addr_9510_7;

Selector_2 s9510_7(wires_2377_6[2], addr_2377_6, addr_positional[38043:38040], addr_9510_7);

wire[31:0] addr_9511_7;

Selector_2 s9511_7(wires_2377_6[3], addr_2377_6, addr_positional[38047:38044], addr_9511_7);

wire[31:0] addr_9512_7;

Selector_2 s9512_7(wires_2378_6[0], addr_2378_6, addr_positional[38051:38048], addr_9512_7);

wire[31:0] addr_9513_7;

Selector_2 s9513_7(wires_2378_6[1], addr_2378_6, addr_positional[38055:38052], addr_9513_7);

wire[31:0] addr_9514_7;

Selector_2 s9514_7(wires_2378_6[2], addr_2378_6, addr_positional[38059:38056], addr_9514_7);

wire[31:0] addr_9515_7;

Selector_2 s9515_7(wires_2378_6[3], addr_2378_6, addr_positional[38063:38060], addr_9515_7);

wire[31:0] addr_9516_7;

Selector_2 s9516_7(wires_2379_6[0], addr_2379_6, addr_positional[38067:38064], addr_9516_7);

wire[31:0] addr_9517_7;

Selector_2 s9517_7(wires_2379_6[1], addr_2379_6, addr_positional[38071:38068], addr_9517_7);

wire[31:0] addr_9518_7;

Selector_2 s9518_7(wires_2379_6[2], addr_2379_6, addr_positional[38075:38072], addr_9518_7);

wire[31:0] addr_9519_7;

Selector_2 s9519_7(wires_2379_6[3], addr_2379_6, addr_positional[38079:38076], addr_9519_7);

wire[31:0] addr_9520_7;

Selector_2 s9520_7(wires_2380_6[0], addr_2380_6, addr_positional[38083:38080], addr_9520_7);

wire[31:0] addr_9521_7;

Selector_2 s9521_7(wires_2380_6[1], addr_2380_6, addr_positional[38087:38084], addr_9521_7);

wire[31:0] addr_9522_7;

Selector_2 s9522_7(wires_2380_6[2], addr_2380_6, addr_positional[38091:38088], addr_9522_7);

wire[31:0] addr_9523_7;

Selector_2 s9523_7(wires_2380_6[3], addr_2380_6, addr_positional[38095:38092], addr_9523_7);

wire[31:0] addr_9524_7;

Selector_2 s9524_7(wires_2381_6[0], addr_2381_6, addr_positional[38099:38096], addr_9524_7);

wire[31:0] addr_9525_7;

Selector_2 s9525_7(wires_2381_6[1], addr_2381_6, addr_positional[38103:38100], addr_9525_7);

wire[31:0] addr_9526_7;

Selector_2 s9526_7(wires_2381_6[2], addr_2381_6, addr_positional[38107:38104], addr_9526_7);

wire[31:0] addr_9527_7;

Selector_2 s9527_7(wires_2381_6[3], addr_2381_6, addr_positional[38111:38108], addr_9527_7);

wire[31:0] addr_9528_7;

Selector_2 s9528_7(wires_2382_6[0], addr_2382_6, addr_positional[38115:38112], addr_9528_7);

wire[31:0] addr_9529_7;

Selector_2 s9529_7(wires_2382_6[1], addr_2382_6, addr_positional[38119:38116], addr_9529_7);

wire[31:0] addr_9530_7;

Selector_2 s9530_7(wires_2382_6[2], addr_2382_6, addr_positional[38123:38120], addr_9530_7);

wire[31:0] addr_9531_7;

Selector_2 s9531_7(wires_2382_6[3], addr_2382_6, addr_positional[38127:38124], addr_9531_7);

wire[31:0] addr_9532_7;

Selector_2 s9532_7(wires_2383_6[0], addr_2383_6, addr_positional[38131:38128], addr_9532_7);

wire[31:0] addr_9533_7;

Selector_2 s9533_7(wires_2383_6[1], addr_2383_6, addr_positional[38135:38132], addr_9533_7);

wire[31:0] addr_9534_7;

Selector_2 s9534_7(wires_2383_6[2], addr_2383_6, addr_positional[38139:38136], addr_9534_7);

wire[31:0] addr_9535_7;

Selector_2 s9535_7(wires_2383_6[3], addr_2383_6, addr_positional[38143:38140], addr_9535_7);

wire[31:0] addr_9536_7;

Selector_2 s9536_7(wires_2384_6[0], addr_2384_6, addr_positional[38147:38144], addr_9536_7);

wire[31:0] addr_9537_7;

Selector_2 s9537_7(wires_2384_6[1], addr_2384_6, addr_positional[38151:38148], addr_9537_7);

wire[31:0] addr_9538_7;

Selector_2 s9538_7(wires_2384_6[2], addr_2384_6, addr_positional[38155:38152], addr_9538_7);

wire[31:0] addr_9539_7;

Selector_2 s9539_7(wires_2384_6[3], addr_2384_6, addr_positional[38159:38156], addr_9539_7);

wire[31:0] addr_9540_7;

Selector_2 s9540_7(wires_2385_6[0], addr_2385_6, addr_positional[38163:38160], addr_9540_7);

wire[31:0] addr_9541_7;

Selector_2 s9541_7(wires_2385_6[1], addr_2385_6, addr_positional[38167:38164], addr_9541_7);

wire[31:0] addr_9542_7;

Selector_2 s9542_7(wires_2385_6[2], addr_2385_6, addr_positional[38171:38168], addr_9542_7);

wire[31:0] addr_9543_7;

Selector_2 s9543_7(wires_2385_6[3], addr_2385_6, addr_positional[38175:38172], addr_9543_7);

wire[31:0] addr_9544_7;

Selector_2 s9544_7(wires_2386_6[0], addr_2386_6, addr_positional[38179:38176], addr_9544_7);

wire[31:0] addr_9545_7;

Selector_2 s9545_7(wires_2386_6[1], addr_2386_6, addr_positional[38183:38180], addr_9545_7);

wire[31:0] addr_9546_7;

Selector_2 s9546_7(wires_2386_6[2], addr_2386_6, addr_positional[38187:38184], addr_9546_7);

wire[31:0] addr_9547_7;

Selector_2 s9547_7(wires_2386_6[3], addr_2386_6, addr_positional[38191:38188], addr_9547_7);

wire[31:0] addr_9548_7;

Selector_2 s9548_7(wires_2387_6[0], addr_2387_6, addr_positional[38195:38192], addr_9548_7);

wire[31:0] addr_9549_7;

Selector_2 s9549_7(wires_2387_6[1], addr_2387_6, addr_positional[38199:38196], addr_9549_7);

wire[31:0] addr_9550_7;

Selector_2 s9550_7(wires_2387_6[2], addr_2387_6, addr_positional[38203:38200], addr_9550_7);

wire[31:0] addr_9551_7;

Selector_2 s9551_7(wires_2387_6[3], addr_2387_6, addr_positional[38207:38204], addr_9551_7);

wire[31:0] addr_9552_7;

Selector_2 s9552_7(wires_2388_6[0], addr_2388_6, addr_positional[38211:38208], addr_9552_7);

wire[31:0] addr_9553_7;

Selector_2 s9553_7(wires_2388_6[1], addr_2388_6, addr_positional[38215:38212], addr_9553_7);

wire[31:0] addr_9554_7;

Selector_2 s9554_7(wires_2388_6[2], addr_2388_6, addr_positional[38219:38216], addr_9554_7);

wire[31:0] addr_9555_7;

Selector_2 s9555_7(wires_2388_6[3], addr_2388_6, addr_positional[38223:38220], addr_9555_7);

wire[31:0] addr_9556_7;

Selector_2 s9556_7(wires_2389_6[0], addr_2389_6, addr_positional[38227:38224], addr_9556_7);

wire[31:0] addr_9557_7;

Selector_2 s9557_7(wires_2389_6[1], addr_2389_6, addr_positional[38231:38228], addr_9557_7);

wire[31:0] addr_9558_7;

Selector_2 s9558_7(wires_2389_6[2], addr_2389_6, addr_positional[38235:38232], addr_9558_7);

wire[31:0] addr_9559_7;

Selector_2 s9559_7(wires_2389_6[3], addr_2389_6, addr_positional[38239:38236], addr_9559_7);

wire[31:0] addr_9560_7;

Selector_2 s9560_7(wires_2390_6[0], addr_2390_6, addr_positional[38243:38240], addr_9560_7);

wire[31:0] addr_9561_7;

Selector_2 s9561_7(wires_2390_6[1], addr_2390_6, addr_positional[38247:38244], addr_9561_7);

wire[31:0] addr_9562_7;

Selector_2 s9562_7(wires_2390_6[2], addr_2390_6, addr_positional[38251:38248], addr_9562_7);

wire[31:0] addr_9563_7;

Selector_2 s9563_7(wires_2390_6[3], addr_2390_6, addr_positional[38255:38252], addr_9563_7);

wire[31:0] addr_9564_7;

Selector_2 s9564_7(wires_2391_6[0], addr_2391_6, addr_positional[38259:38256], addr_9564_7);

wire[31:0] addr_9565_7;

Selector_2 s9565_7(wires_2391_6[1], addr_2391_6, addr_positional[38263:38260], addr_9565_7);

wire[31:0] addr_9566_7;

Selector_2 s9566_7(wires_2391_6[2], addr_2391_6, addr_positional[38267:38264], addr_9566_7);

wire[31:0] addr_9567_7;

Selector_2 s9567_7(wires_2391_6[3], addr_2391_6, addr_positional[38271:38268], addr_9567_7);

wire[31:0] addr_9568_7;

Selector_2 s9568_7(wires_2392_6[0], addr_2392_6, addr_positional[38275:38272], addr_9568_7);

wire[31:0] addr_9569_7;

Selector_2 s9569_7(wires_2392_6[1], addr_2392_6, addr_positional[38279:38276], addr_9569_7);

wire[31:0] addr_9570_7;

Selector_2 s9570_7(wires_2392_6[2], addr_2392_6, addr_positional[38283:38280], addr_9570_7);

wire[31:0] addr_9571_7;

Selector_2 s9571_7(wires_2392_6[3], addr_2392_6, addr_positional[38287:38284], addr_9571_7);

wire[31:0] addr_9572_7;

Selector_2 s9572_7(wires_2393_6[0], addr_2393_6, addr_positional[38291:38288], addr_9572_7);

wire[31:0] addr_9573_7;

Selector_2 s9573_7(wires_2393_6[1], addr_2393_6, addr_positional[38295:38292], addr_9573_7);

wire[31:0] addr_9574_7;

Selector_2 s9574_7(wires_2393_6[2], addr_2393_6, addr_positional[38299:38296], addr_9574_7);

wire[31:0] addr_9575_7;

Selector_2 s9575_7(wires_2393_6[3], addr_2393_6, addr_positional[38303:38300], addr_9575_7);

wire[31:0] addr_9576_7;

Selector_2 s9576_7(wires_2394_6[0], addr_2394_6, addr_positional[38307:38304], addr_9576_7);

wire[31:0] addr_9577_7;

Selector_2 s9577_7(wires_2394_6[1], addr_2394_6, addr_positional[38311:38308], addr_9577_7);

wire[31:0] addr_9578_7;

Selector_2 s9578_7(wires_2394_6[2], addr_2394_6, addr_positional[38315:38312], addr_9578_7);

wire[31:0] addr_9579_7;

Selector_2 s9579_7(wires_2394_6[3], addr_2394_6, addr_positional[38319:38316], addr_9579_7);

wire[31:0] addr_9580_7;

Selector_2 s9580_7(wires_2395_6[0], addr_2395_6, addr_positional[38323:38320], addr_9580_7);

wire[31:0] addr_9581_7;

Selector_2 s9581_7(wires_2395_6[1], addr_2395_6, addr_positional[38327:38324], addr_9581_7);

wire[31:0] addr_9582_7;

Selector_2 s9582_7(wires_2395_6[2], addr_2395_6, addr_positional[38331:38328], addr_9582_7);

wire[31:0] addr_9583_7;

Selector_2 s9583_7(wires_2395_6[3], addr_2395_6, addr_positional[38335:38332], addr_9583_7);

wire[31:0] addr_9584_7;

Selector_2 s9584_7(wires_2396_6[0], addr_2396_6, addr_positional[38339:38336], addr_9584_7);

wire[31:0] addr_9585_7;

Selector_2 s9585_7(wires_2396_6[1], addr_2396_6, addr_positional[38343:38340], addr_9585_7);

wire[31:0] addr_9586_7;

Selector_2 s9586_7(wires_2396_6[2], addr_2396_6, addr_positional[38347:38344], addr_9586_7);

wire[31:0] addr_9587_7;

Selector_2 s9587_7(wires_2396_6[3], addr_2396_6, addr_positional[38351:38348], addr_9587_7);

wire[31:0] addr_9588_7;

Selector_2 s9588_7(wires_2397_6[0], addr_2397_6, addr_positional[38355:38352], addr_9588_7);

wire[31:0] addr_9589_7;

Selector_2 s9589_7(wires_2397_6[1], addr_2397_6, addr_positional[38359:38356], addr_9589_7);

wire[31:0] addr_9590_7;

Selector_2 s9590_7(wires_2397_6[2], addr_2397_6, addr_positional[38363:38360], addr_9590_7);

wire[31:0] addr_9591_7;

Selector_2 s9591_7(wires_2397_6[3], addr_2397_6, addr_positional[38367:38364], addr_9591_7);

wire[31:0] addr_9592_7;

Selector_2 s9592_7(wires_2398_6[0], addr_2398_6, addr_positional[38371:38368], addr_9592_7);

wire[31:0] addr_9593_7;

Selector_2 s9593_7(wires_2398_6[1], addr_2398_6, addr_positional[38375:38372], addr_9593_7);

wire[31:0] addr_9594_7;

Selector_2 s9594_7(wires_2398_6[2], addr_2398_6, addr_positional[38379:38376], addr_9594_7);

wire[31:0] addr_9595_7;

Selector_2 s9595_7(wires_2398_6[3], addr_2398_6, addr_positional[38383:38380], addr_9595_7);

wire[31:0] addr_9596_7;

Selector_2 s9596_7(wires_2399_6[0], addr_2399_6, addr_positional[38387:38384], addr_9596_7);

wire[31:0] addr_9597_7;

Selector_2 s9597_7(wires_2399_6[1], addr_2399_6, addr_positional[38391:38388], addr_9597_7);

wire[31:0] addr_9598_7;

Selector_2 s9598_7(wires_2399_6[2], addr_2399_6, addr_positional[38395:38392], addr_9598_7);

wire[31:0] addr_9599_7;

Selector_2 s9599_7(wires_2399_6[3], addr_2399_6, addr_positional[38399:38396], addr_9599_7);

wire[31:0] addr_9600_7;

Selector_2 s9600_7(wires_2400_6[0], addr_2400_6, addr_positional[38403:38400], addr_9600_7);

wire[31:0] addr_9601_7;

Selector_2 s9601_7(wires_2400_6[1], addr_2400_6, addr_positional[38407:38404], addr_9601_7);

wire[31:0] addr_9602_7;

Selector_2 s9602_7(wires_2400_6[2], addr_2400_6, addr_positional[38411:38408], addr_9602_7);

wire[31:0] addr_9603_7;

Selector_2 s9603_7(wires_2400_6[3], addr_2400_6, addr_positional[38415:38412], addr_9603_7);

wire[31:0] addr_9604_7;

Selector_2 s9604_7(wires_2401_6[0], addr_2401_6, addr_positional[38419:38416], addr_9604_7);

wire[31:0] addr_9605_7;

Selector_2 s9605_7(wires_2401_6[1], addr_2401_6, addr_positional[38423:38420], addr_9605_7);

wire[31:0] addr_9606_7;

Selector_2 s9606_7(wires_2401_6[2], addr_2401_6, addr_positional[38427:38424], addr_9606_7);

wire[31:0] addr_9607_7;

Selector_2 s9607_7(wires_2401_6[3], addr_2401_6, addr_positional[38431:38428], addr_9607_7);

wire[31:0] addr_9608_7;

Selector_2 s9608_7(wires_2402_6[0], addr_2402_6, addr_positional[38435:38432], addr_9608_7);

wire[31:0] addr_9609_7;

Selector_2 s9609_7(wires_2402_6[1], addr_2402_6, addr_positional[38439:38436], addr_9609_7);

wire[31:0] addr_9610_7;

Selector_2 s9610_7(wires_2402_6[2], addr_2402_6, addr_positional[38443:38440], addr_9610_7);

wire[31:0] addr_9611_7;

Selector_2 s9611_7(wires_2402_6[3], addr_2402_6, addr_positional[38447:38444], addr_9611_7);

wire[31:0] addr_9612_7;

Selector_2 s9612_7(wires_2403_6[0], addr_2403_6, addr_positional[38451:38448], addr_9612_7);

wire[31:0] addr_9613_7;

Selector_2 s9613_7(wires_2403_6[1], addr_2403_6, addr_positional[38455:38452], addr_9613_7);

wire[31:0] addr_9614_7;

Selector_2 s9614_7(wires_2403_6[2], addr_2403_6, addr_positional[38459:38456], addr_9614_7);

wire[31:0] addr_9615_7;

Selector_2 s9615_7(wires_2403_6[3], addr_2403_6, addr_positional[38463:38460], addr_9615_7);

wire[31:0] addr_9616_7;

Selector_2 s9616_7(wires_2404_6[0], addr_2404_6, addr_positional[38467:38464], addr_9616_7);

wire[31:0] addr_9617_7;

Selector_2 s9617_7(wires_2404_6[1], addr_2404_6, addr_positional[38471:38468], addr_9617_7);

wire[31:0] addr_9618_7;

Selector_2 s9618_7(wires_2404_6[2], addr_2404_6, addr_positional[38475:38472], addr_9618_7);

wire[31:0] addr_9619_7;

Selector_2 s9619_7(wires_2404_6[3], addr_2404_6, addr_positional[38479:38476], addr_9619_7);

wire[31:0] addr_9620_7;

Selector_2 s9620_7(wires_2405_6[0], addr_2405_6, addr_positional[38483:38480], addr_9620_7);

wire[31:0] addr_9621_7;

Selector_2 s9621_7(wires_2405_6[1], addr_2405_6, addr_positional[38487:38484], addr_9621_7);

wire[31:0] addr_9622_7;

Selector_2 s9622_7(wires_2405_6[2], addr_2405_6, addr_positional[38491:38488], addr_9622_7);

wire[31:0] addr_9623_7;

Selector_2 s9623_7(wires_2405_6[3], addr_2405_6, addr_positional[38495:38492], addr_9623_7);

wire[31:0] addr_9624_7;

Selector_2 s9624_7(wires_2406_6[0], addr_2406_6, addr_positional[38499:38496], addr_9624_7);

wire[31:0] addr_9625_7;

Selector_2 s9625_7(wires_2406_6[1], addr_2406_6, addr_positional[38503:38500], addr_9625_7);

wire[31:0] addr_9626_7;

Selector_2 s9626_7(wires_2406_6[2], addr_2406_6, addr_positional[38507:38504], addr_9626_7);

wire[31:0] addr_9627_7;

Selector_2 s9627_7(wires_2406_6[3], addr_2406_6, addr_positional[38511:38508], addr_9627_7);

wire[31:0] addr_9628_7;

Selector_2 s9628_7(wires_2407_6[0], addr_2407_6, addr_positional[38515:38512], addr_9628_7);

wire[31:0] addr_9629_7;

Selector_2 s9629_7(wires_2407_6[1], addr_2407_6, addr_positional[38519:38516], addr_9629_7);

wire[31:0] addr_9630_7;

Selector_2 s9630_7(wires_2407_6[2], addr_2407_6, addr_positional[38523:38520], addr_9630_7);

wire[31:0] addr_9631_7;

Selector_2 s9631_7(wires_2407_6[3], addr_2407_6, addr_positional[38527:38524], addr_9631_7);

wire[31:0] addr_9632_7;

Selector_2 s9632_7(wires_2408_6[0], addr_2408_6, addr_positional[38531:38528], addr_9632_7);

wire[31:0] addr_9633_7;

Selector_2 s9633_7(wires_2408_6[1], addr_2408_6, addr_positional[38535:38532], addr_9633_7);

wire[31:0] addr_9634_7;

Selector_2 s9634_7(wires_2408_6[2], addr_2408_6, addr_positional[38539:38536], addr_9634_7);

wire[31:0] addr_9635_7;

Selector_2 s9635_7(wires_2408_6[3], addr_2408_6, addr_positional[38543:38540], addr_9635_7);

wire[31:0] addr_9636_7;

Selector_2 s9636_7(wires_2409_6[0], addr_2409_6, addr_positional[38547:38544], addr_9636_7);

wire[31:0] addr_9637_7;

Selector_2 s9637_7(wires_2409_6[1], addr_2409_6, addr_positional[38551:38548], addr_9637_7);

wire[31:0] addr_9638_7;

Selector_2 s9638_7(wires_2409_6[2], addr_2409_6, addr_positional[38555:38552], addr_9638_7);

wire[31:0] addr_9639_7;

Selector_2 s9639_7(wires_2409_6[3], addr_2409_6, addr_positional[38559:38556], addr_9639_7);

wire[31:0] addr_9640_7;

Selector_2 s9640_7(wires_2410_6[0], addr_2410_6, addr_positional[38563:38560], addr_9640_7);

wire[31:0] addr_9641_7;

Selector_2 s9641_7(wires_2410_6[1], addr_2410_6, addr_positional[38567:38564], addr_9641_7);

wire[31:0] addr_9642_7;

Selector_2 s9642_7(wires_2410_6[2], addr_2410_6, addr_positional[38571:38568], addr_9642_7);

wire[31:0] addr_9643_7;

Selector_2 s9643_7(wires_2410_6[3], addr_2410_6, addr_positional[38575:38572], addr_9643_7);

wire[31:0] addr_9644_7;

Selector_2 s9644_7(wires_2411_6[0], addr_2411_6, addr_positional[38579:38576], addr_9644_7);

wire[31:0] addr_9645_7;

Selector_2 s9645_7(wires_2411_6[1], addr_2411_6, addr_positional[38583:38580], addr_9645_7);

wire[31:0] addr_9646_7;

Selector_2 s9646_7(wires_2411_6[2], addr_2411_6, addr_positional[38587:38584], addr_9646_7);

wire[31:0] addr_9647_7;

Selector_2 s9647_7(wires_2411_6[3], addr_2411_6, addr_positional[38591:38588], addr_9647_7);

wire[31:0] addr_9648_7;

Selector_2 s9648_7(wires_2412_6[0], addr_2412_6, addr_positional[38595:38592], addr_9648_7);

wire[31:0] addr_9649_7;

Selector_2 s9649_7(wires_2412_6[1], addr_2412_6, addr_positional[38599:38596], addr_9649_7);

wire[31:0] addr_9650_7;

Selector_2 s9650_7(wires_2412_6[2], addr_2412_6, addr_positional[38603:38600], addr_9650_7);

wire[31:0] addr_9651_7;

Selector_2 s9651_7(wires_2412_6[3], addr_2412_6, addr_positional[38607:38604], addr_9651_7);

wire[31:0] addr_9652_7;

Selector_2 s9652_7(wires_2413_6[0], addr_2413_6, addr_positional[38611:38608], addr_9652_7);

wire[31:0] addr_9653_7;

Selector_2 s9653_7(wires_2413_6[1], addr_2413_6, addr_positional[38615:38612], addr_9653_7);

wire[31:0] addr_9654_7;

Selector_2 s9654_7(wires_2413_6[2], addr_2413_6, addr_positional[38619:38616], addr_9654_7);

wire[31:0] addr_9655_7;

Selector_2 s9655_7(wires_2413_6[3], addr_2413_6, addr_positional[38623:38620], addr_9655_7);

wire[31:0] addr_9656_7;

Selector_2 s9656_7(wires_2414_6[0], addr_2414_6, addr_positional[38627:38624], addr_9656_7);

wire[31:0] addr_9657_7;

Selector_2 s9657_7(wires_2414_6[1], addr_2414_6, addr_positional[38631:38628], addr_9657_7);

wire[31:0] addr_9658_7;

Selector_2 s9658_7(wires_2414_6[2], addr_2414_6, addr_positional[38635:38632], addr_9658_7);

wire[31:0] addr_9659_7;

Selector_2 s9659_7(wires_2414_6[3], addr_2414_6, addr_positional[38639:38636], addr_9659_7);

wire[31:0] addr_9660_7;

Selector_2 s9660_7(wires_2415_6[0], addr_2415_6, addr_positional[38643:38640], addr_9660_7);

wire[31:0] addr_9661_7;

Selector_2 s9661_7(wires_2415_6[1], addr_2415_6, addr_positional[38647:38644], addr_9661_7);

wire[31:0] addr_9662_7;

Selector_2 s9662_7(wires_2415_6[2], addr_2415_6, addr_positional[38651:38648], addr_9662_7);

wire[31:0] addr_9663_7;

Selector_2 s9663_7(wires_2415_6[3], addr_2415_6, addr_positional[38655:38652], addr_9663_7);

wire[31:0] addr_9664_7;

Selector_2 s9664_7(wires_2416_6[0], addr_2416_6, addr_positional[38659:38656], addr_9664_7);

wire[31:0] addr_9665_7;

Selector_2 s9665_7(wires_2416_6[1], addr_2416_6, addr_positional[38663:38660], addr_9665_7);

wire[31:0] addr_9666_7;

Selector_2 s9666_7(wires_2416_6[2], addr_2416_6, addr_positional[38667:38664], addr_9666_7);

wire[31:0] addr_9667_7;

Selector_2 s9667_7(wires_2416_6[3], addr_2416_6, addr_positional[38671:38668], addr_9667_7);

wire[31:0] addr_9668_7;

Selector_2 s9668_7(wires_2417_6[0], addr_2417_6, addr_positional[38675:38672], addr_9668_7);

wire[31:0] addr_9669_7;

Selector_2 s9669_7(wires_2417_6[1], addr_2417_6, addr_positional[38679:38676], addr_9669_7);

wire[31:0] addr_9670_7;

Selector_2 s9670_7(wires_2417_6[2], addr_2417_6, addr_positional[38683:38680], addr_9670_7);

wire[31:0] addr_9671_7;

Selector_2 s9671_7(wires_2417_6[3], addr_2417_6, addr_positional[38687:38684], addr_9671_7);

wire[31:0] addr_9672_7;

Selector_2 s9672_7(wires_2418_6[0], addr_2418_6, addr_positional[38691:38688], addr_9672_7);

wire[31:0] addr_9673_7;

Selector_2 s9673_7(wires_2418_6[1], addr_2418_6, addr_positional[38695:38692], addr_9673_7);

wire[31:0] addr_9674_7;

Selector_2 s9674_7(wires_2418_6[2], addr_2418_6, addr_positional[38699:38696], addr_9674_7);

wire[31:0] addr_9675_7;

Selector_2 s9675_7(wires_2418_6[3], addr_2418_6, addr_positional[38703:38700], addr_9675_7);

wire[31:0] addr_9676_7;

Selector_2 s9676_7(wires_2419_6[0], addr_2419_6, addr_positional[38707:38704], addr_9676_7);

wire[31:0] addr_9677_7;

Selector_2 s9677_7(wires_2419_6[1], addr_2419_6, addr_positional[38711:38708], addr_9677_7);

wire[31:0] addr_9678_7;

Selector_2 s9678_7(wires_2419_6[2], addr_2419_6, addr_positional[38715:38712], addr_9678_7);

wire[31:0] addr_9679_7;

Selector_2 s9679_7(wires_2419_6[3], addr_2419_6, addr_positional[38719:38716], addr_9679_7);

wire[31:0] addr_9680_7;

Selector_2 s9680_7(wires_2420_6[0], addr_2420_6, addr_positional[38723:38720], addr_9680_7);

wire[31:0] addr_9681_7;

Selector_2 s9681_7(wires_2420_6[1], addr_2420_6, addr_positional[38727:38724], addr_9681_7);

wire[31:0] addr_9682_7;

Selector_2 s9682_7(wires_2420_6[2], addr_2420_6, addr_positional[38731:38728], addr_9682_7);

wire[31:0] addr_9683_7;

Selector_2 s9683_7(wires_2420_6[3], addr_2420_6, addr_positional[38735:38732], addr_9683_7);

wire[31:0] addr_9684_7;

Selector_2 s9684_7(wires_2421_6[0], addr_2421_6, addr_positional[38739:38736], addr_9684_7);

wire[31:0] addr_9685_7;

Selector_2 s9685_7(wires_2421_6[1], addr_2421_6, addr_positional[38743:38740], addr_9685_7);

wire[31:0] addr_9686_7;

Selector_2 s9686_7(wires_2421_6[2], addr_2421_6, addr_positional[38747:38744], addr_9686_7);

wire[31:0] addr_9687_7;

Selector_2 s9687_7(wires_2421_6[3], addr_2421_6, addr_positional[38751:38748], addr_9687_7);

wire[31:0] addr_9688_7;

Selector_2 s9688_7(wires_2422_6[0], addr_2422_6, addr_positional[38755:38752], addr_9688_7);

wire[31:0] addr_9689_7;

Selector_2 s9689_7(wires_2422_6[1], addr_2422_6, addr_positional[38759:38756], addr_9689_7);

wire[31:0] addr_9690_7;

Selector_2 s9690_7(wires_2422_6[2], addr_2422_6, addr_positional[38763:38760], addr_9690_7);

wire[31:0] addr_9691_7;

Selector_2 s9691_7(wires_2422_6[3], addr_2422_6, addr_positional[38767:38764], addr_9691_7);

wire[31:0] addr_9692_7;

Selector_2 s9692_7(wires_2423_6[0], addr_2423_6, addr_positional[38771:38768], addr_9692_7);

wire[31:0] addr_9693_7;

Selector_2 s9693_7(wires_2423_6[1], addr_2423_6, addr_positional[38775:38772], addr_9693_7);

wire[31:0] addr_9694_7;

Selector_2 s9694_7(wires_2423_6[2], addr_2423_6, addr_positional[38779:38776], addr_9694_7);

wire[31:0] addr_9695_7;

Selector_2 s9695_7(wires_2423_6[3], addr_2423_6, addr_positional[38783:38780], addr_9695_7);

wire[31:0] addr_9696_7;

Selector_2 s9696_7(wires_2424_6[0], addr_2424_6, addr_positional[38787:38784], addr_9696_7);

wire[31:0] addr_9697_7;

Selector_2 s9697_7(wires_2424_6[1], addr_2424_6, addr_positional[38791:38788], addr_9697_7);

wire[31:0] addr_9698_7;

Selector_2 s9698_7(wires_2424_6[2], addr_2424_6, addr_positional[38795:38792], addr_9698_7);

wire[31:0] addr_9699_7;

Selector_2 s9699_7(wires_2424_6[3], addr_2424_6, addr_positional[38799:38796], addr_9699_7);

wire[31:0] addr_9700_7;

Selector_2 s9700_7(wires_2425_6[0], addr_2425_6, addr_positional[38803:38800], addr_9700_7);

wire[31:0] addr_9701_7;

Selector_2 s9701_7(wires_2425_6[1], addr_2425_6, addr_positional[38807:38804], addr_9701_7);

wire[31:0] addr_9702_7;

Selector_2 s9702_7(wires_2425_6[2], addr_2425_6, addr_positional[38811:38808], addr_9702_7);

wire[31:0] addr_9703_7;

Selector_2 s9703_7(wires_2425_6[3], addr_2425_6, addr_positional[38815:38812], addr_9703_7);

wire[31:0] addr_9704_7;

Selector_2 s9704_7(wires_2426_6[0], addr_2426_6, addr_positional[38819:38816], addr_9704_7);

wire[31:0] addr_9705_7;

Selector_2 s9705_7(wires_2426_6[1], addr_2426_6, addr_positional[38823:38820], addr_9705_7);

wire[31:0] addr_9706_7;

Selector_2 s9706_7(wires_2426_6[2], addr_2426_6, addr_positional[38827:38824], addr_9706_7);

wire[31:0] addr_9707_7;

Selector_2 s9707_7(wires_2426_6[3], addr_2426_6, addr_positional[38831:38828], addr_9707_7);

wire[31:0] addr_9708_7;

Selector_2 s9708_7(wires_2427_6[0], addr_2427_6, addr_positional[38835:38832], addr_9708_7);

wire[31:0] addr_9709_7;

Selector_2 s9709_7(wires_2427_6[1], addr_2427_6, addr_positional[38839:38836], addr_9709_7);

wire[31:0] addr_9710_7;

Selector_2 s9710_7(wires_2427_6[2], addr_2427_6, addr_positional[38843:38840], addr_9710_7);

wire[31:0] addr_9711_7;

Selector_2 s9711_7(wires_2427_6[3], addr_2427_6, addr_positional[38847:38844], addr_9711_7);

wire[31:0] addr_9712_7;

Selector_2 s9712_7(wires_2428_6[0], addr_2428_6, addr_positional[38851:38848], addr_9712_7);

wire[31:0] addr_9713_7;

Selector_2 s9713_7(wires_2428_6[1], addr_2428_6, addr_positional[38855:38852], addr_9713_7);

wire[31:0] addr_9714_7;

Selector_2 s9714_7(wires_2428_6[2], addr_2428_6, addr_positional[38859:38856], addr_9714_7);

wire[31:0] addr_9715_7;

Selector_2 s9715_7(wires_2428_6[3], addr_2428_6, addr_positional[38863:38860], addr_9715_7);

wire[31:0] addr_9716_7;

Selector_2 s9716_7(wires_2429_6[0], addr_2429_6, addr_positional[38867:38864], addr_9716_7);

wire[31:0] addr_9717_7;

Selector_2 s9717_7(wires_2429_6[1], addr_2429_6, addr_positional[38871:38868], addr_9717_7);

wire[31:0] addr_9718_7;

Selector_2 s9718_7(wires_2429_6[2], addr_2429_6, addr_positional[38875:38872], addr_9718_7);

wire[31:0] addr_9719_7;

Selector_2 s9719_7(wires_2429_6[3], addr_2429_6, addr_positional[38879:38876], addr_9719_7);

wire[31:0] addr_9720_7;

Selector_2 s9720_7(wires_2430_6[0], addr_2430_6, addr_positional[38883:38880], addr_9720_7);

wire[31:0] addr_9721_7;

Selector_2 s9721_7(wires_2430_6[1], addr_2430_6, addr_positional[38887:38884], addr_9721_7);

wire[31:0] addr_9722_7;

Selector_2 s9722_7(wires_2430_6[2], addr_2430_6, addr_positional[38891:38888], addr_9722_7);

wire[31:0] addr_9723_7;

Selector_2 s9723_7(wires_2430_6[3], addr_2430_6, addr_positional[38895:38892], addr_9723_7);

wire[31:0] addr_9724_7;

Selector_2 s9724_7(wires_2431_6[0], addr_2431_6, addr_positional[38899:38896], addr_9724_7);

wire[31:0] addr_9725_7;

Selector_2 s9725_7(wires_2431_6[1], addr_2431_6, addr_positional[38903:38900], addr_9725_7);

wire[31:0] addr_9726_7;

Selector_2 s9726_7(wires_2431_6[2], addr_2431_6, addr_positional[38907:38904], addr_9726_7);

wire[31:0] addr_9727_7;

Selector_2 s9727_7(wires_2431_6[3], addr_2431_6, addr_positional[38911:38908], addr_9727_7);

wire[31:0] addr_9728_7;

Selector_2 s9728_7(wires_2432_6[0], addr_2432_6, addr_positional[38915:38912], addr_9728_7);

wire[31:0] addr_9729_7;

Selector_2 s9729_7(wires_2432_6[1], addr_2432_6, addr_positional[38919:38916], addr_9729_7);

wire[31:0] addr_9730_7;

Selector_2 s9730_7(wires_2432_6[2], addr_2432_6, addr_positional[38923:38920], addr_9730_7);

wire[31:0] addr_9731_7;

Selector_2 s9731_7(wires_2432_6[3], addr_2432_6, addr_positional[38927:38924], addr_9731_7);

wire[31:0] addr_9732_7;

Selector_2 s9732_7(wires_2433_6[0], addr_2433_6, addr_positional[38931:38928], addr_9732_7);

wire[31:0] addr_9733_7;

Selector_2 s9733_7(wires_2433_6[1], addr_2433_6, addr_positional[38935:38932], addr_9733_7);

wire[31:0] addr_9734_7;

Selector_2 s9734_7(wires_2433_6[2], addr_2433_6, addr_positional[38939:38936], addr_9734_7);

wire[31:0] addr_9735_7;

Selector_2 s9735_7(wires_2433_6[3], addr_2433_6, addr_positional[38943:38940], addr_9735_7);

wire[31:0] addr_9736_7;

Selector_2 s9736_7(wires_2434_6[0], addr_2434_6, addr_positional[38947:38944], addr_9736_7);

wire[31:0] addr_9737_7;

Selector_2 s9737_7(wires_2434_6[1], addr_2434_6, addr_positional[38951:38948], addr_9737_7);

wire[31:0] addr_9738_7;

Selector_2 s9738_7(wires_2434_6[2], addr_2434_6, addr_positional[38955:38952], addr_9738_7);

wire[31:0] addr_9739_7;

Selector_2 s9739_7(wires_2434_6[3], addr_2434_6, addr_positional[38959:38956], addr_9739_7);

wire[31:0] addr_9740_7;

Selector_2 s9740_7(wires_2435_6[0], addr_2435_6, addr_positional[38963:38960], addr_9740_7);

wire[31:0] addr_9741_7;

Selector_2 s9741_7(wires_2435_6[1], addr_2435_6, addr_positional[38967:38964], addr_9741_7);

wire[31:0] addr_9742_7;

Selector_2 s9742_7(wires_2435_6[2], addr_2435_6, addr_positional[38971:38968], addr_9742_7);

wire[31:0] addr_9743_7;

Selector_2 s9743_7(wires_2435_6[3], addr_2435_6, addr_positional[38975:38972], addr_9743_7);

wire[31:0] addr_9744_7;

Selector_2 s9744_7(wires_2436_6[0], addr_2436_6, addr_positional[38979:38976], addr_9744_7);

wire[31:0] addr_9745_7;

Selector_2 s9745_7(wires_2436_6[1], addr_2436_6, addr_positional[38983:38980], addr_9745_7);

wire[31:0] addr_9746_7;

Selector_2 s9746_7(wires_2436_6[2], addr_2436_6, addr_positional[38987:38984], addr_9746_7);

wire[31:0] addr_9747_7;

Selector_2 s9747_7(wires_2436_6[3], addr_2436_6, addr_positional[38991:38988], addr_9747_7);

wire[31:0] addr_9748_7;

Selector_2 s9748_7(wires_2437_6[0], addr_2437_6, addr_positional[38995:38992], addr_9748_7);

wire[31:0] addr_9749_7;

Selector_2 s9749_7(wires_2437_6[1], addr_2437_6, addr_positional[38999:38996], addr_9749_7);

wire[31:0] addr_9750_7;

Selector_2 s9750_7(wires_2437_6[2], addr_2437_6, addr_positional[39003:39000], addr_9750_7);

wire[31:0] addr_9751_7;

Selector_2 s9751_7(wires_2437_6[3], addr_2437_6, addr_positional[39007:39004], addr_9751_7);

wire[31:0] addr_9752_7;

Selector_2 s9752_7(wires_2438_6[0], addr_2438_6, addr_positional[39011:39008], addr_9752_7);

wire[31:0] addr_9753_7;

Selector_2 s9753_7(wires_2438_6[1], addr_2438_6, addr_positional[39015:39012], addr_9753_7);

wire[31:0] addr_9754_7;

Selector_2 s9754_7(wires_2438_6[2], addr_2438_6, addr_positional[39019:39016], addr_9754_7);

wire[31:0] addr_9755_7;

Selector_2 s9755_7(wires_2438_6[3], addr_2438_6, addr_positional[39023:39020], addr_9755_7);

wire[31:0] addr_9756_7;

Selector_2 s9756_7(wires_2439_6[0], addr_2439_6, addr_positional[39027:39024], addr_9756_7);

wire[31:0] addr_9757_7;

Selector_2 s9757_7(wires_2439_6[1], addr_2439_6, addr_positional[39031:39028], addr_9757_7);

wire[31:0] addr_9758_7;

Selector_2 s9758_7(wires_2439_6[2], addr_2439_6, addr_positional[39035:39032], addr_9758_7);

wire[31:0] addr_9759_7;

Selector_2 s9759_7(wires_2439_6[3], addr_2439_6, addr_positional[39039:39036], addr_9759_7);

wire[31:0] addr_9760_7;

Selector_2 s9760_7(wires_2440_6[0], addr_2440_6, addr_positional[39043:39040], addr_9760_7);

wire[31:0] addr_9761_7;

Selector_2 s9761_7(wires_2440_6[1], addr_2440_6, addr_positional[39047:39044], addr_9761_7);

wire[31:0] addr_9762_7;

Selector_2 s9762_7(wires_2440_6[2], addr_2440_6, addr_positional[39051:39048], addr_9762_7);

wire[31:0] addr_9763_7;

Selector_2 s9763_7(wires_2440_6[3], addr_2440_6, addr_positional[39055:39052], addr_9763_7);

wire[31:0] addr_9764_7;

Selector_2 s9764_7(wires_2441_6[0], addr_2441_6, addr_positional[39059:39056], addr_9764_7);

wire[31:0] addr_9765_7;

Selector_2 s9765_7(wires_2441_6[1], addr_2441_6, addr_positional[39063:39060], addr_9765_7);

wire[31:0] addr_9766_7;

Selector_2 s9766_7(wires_2441_6[2], addr_2441_6, addr_positional[39067:39064], addr_9766_7);

wire[31:0] addr_9767_7;

Selector_2 s9767_7(wires_2441_6[3], addr_2441_6, addr_positional[39071:39068], addr_9767_7);

wire[31:0] addr_9768_7;

Selector_2 s9768_7(wires_2442_6[0], addr_2442_6, addr_positional[39075:39072], addr_9768_7);

wire[31:0] addr_9769_7;

Selector_2 s9769_7(wires_2442_6[1], addr_2442_6, addr_positional[39079:39076], addr_9769_7);

wire[31:0] addr_9770_7;

Selector_2 s9770_7(wires_2442_6[2], addr_2442_6, addr_positional[39083:39080], addr_9770_7);

wire[31:0] addr_9771_7;

Selector_2 s9771_7(wires_2442_6[3], addr_2442_6, addr_positional[39087:39084], addr_9771_7);

wire[31:0] addr_9772_7;

Selector_2 s9772_7(wires_2443_6[0], addr_2443_6, addr_positional[39091:39088], addr_9772_7);

wire[31:0] addr_9773_7;

Selector_2 s9773_7(wires_2443_6[1], addr_2443_6, addr_positional[39095:39092], addr_9773_7);

wire[31:0] addr_9774_7;

Selector_2 s9774_7(wires_2443_6[2], addr_2443_6, addr_positional[39099:39096], addr_9774_7);

wire[31:0] addr_9775_7;

Selector_2 s9775_7(wires_2443_6[3], addr_2443_6, addr_positional[39103:39100], addr_9775_7);

wire[31:0] addr_9776_7;

Selector_2 s9776_7(wires_2444_6[0], addr_2444_6, addr_positional[39107:39104], addr_9776_7);

wire[31:0] addr_9777_7;

Selector_2 s9777_7(wires_2444_6[1], addr_2444_6, addr_positional[39111:39108], addr_9777_7);

wire[31:0] addr_9778_7;

Selector_2 s9778_7(wires_2444_6[2], addr_2444_6, addr_positional[39115:39112], addr_9778_7);

wire[31:0] addr_9779_7;

Selector_2 s9779_7(wires_2444_6[3], addr_2444_6, addr_positional[39119:39116], addr_9779_7);

wire[31:0] addr_9780_7;

Selector_2 s9780_7(wires_2445_6[0], addr_2445_6, addr_positional[39123:39120], addr_9780_7);

wire[31:0] addr_9781_7;

Selector_2 s9781_7(wires_2445_6[1], addr_2445_6, addr_positional[39127:39124], addr_9781_7);

wire[31:0] addr_9782_7;

Selector_2 s9782_7(wires_2445_6[2], addr_2445_6, addr_positional[39131:39128], addr_9782_7);

wire[31:0] addr_9783_7;

Selector_2 s9783_7(wires_2445_6[3], addr_2445_6, addr_positional[39135:39132], addr_9783_7);

wire[31:0] addr_9784_7;

Selector_2 s9784_7(wires_2446_6[0], addr_2446_6, addr_positional[39139:39136], addr_9784_7);

wire[31:0] addr_9785_7;

Selector_2 s9785_7(wires_2446_6[1], addr_2446_6, addr_positional[39143:39140], addr_9785_7);

wire[31:0] addr_9786_7;

Selector_2 s9786_7(wires_2446_6[2], addr_2446_6, addr_positional[39147:39144], addr_9786_7);

wire[31:0] addr_9787_7;

Selector_2 s9787_7(wires_2446_6[3], addr_2446_6, addr_positional[39151:39148], addr_9787_7);

wire[31:0] addr_9788_7;

Selector_2 s9788_7(wires_2447_6[0], addr_2447_6, addr_positional[39155:39152], addr_9788_7);

wire[31:0] addr_9789_7;

Selector_2 s9789_7(wires_2447_6[1], addr_2447_6, addr_positional[39159:39156], addr_9789_7);

wire[31:0] addr_9790_7;

Selector_2 s9790_7(wires_2447_6[2], addr_2447_6, addr_positional[39163:39160], addr_9790_7);

wire[31:0] addr_9791_7;

Selector_2 s9791_7(wires_2447_6[3], addr_2447_6, addr_positional[39167:39164], addr_9791_7);

wire[31:0] addr_9792_7;

Selector_2 s9792_7(wires_2448_6[0], addr_2448_6, addr_positional[39171:39168], addr_9792_7);

wire[31:0] addr_9793_7;

Selector_2 s9793_7(wires_2448_6[1], addr_2448_6, addr_positional[39175:39172], addr_9793_7);

wire[31:0] addr_9794_7;

Selector_2 s9794_7(wires_2448_6[2], addr_2448_6, addr_positional[39179:39176], addr_9794_7);

wire[31:0] addr_9795_7;

Selector_2 s9795_7(wires_2448_6[3], addr_2448_6, addr_positional[39183:39180], addr_9795_7);

wire[31:0] addr_9796_7;

Selector_2 s9796_7(wires_2449_6[0], addr_2449_6, addr_positional[39187:39184], addr_9796_7);

wire[31:0] addr_9797_7;

Selector_2 s9797_7(wires_2449_6[1], addr_2449_6, addr_positional[39191:39188], addr_9797_7);

wire[31:0] addr_9798_7;

Selector_2 s9798_7(wires_2449_6[2], addr_2449_6, addr_positional[39195:39192], addr_9798_7);

wire[31:0] addr_9799_7;

Selector_2 s9799_7(wires_2449_6[3], addr_2449_6, addr_positional[39199:39196], addr_9799_7);

wire[31:0] addr_9800_7;

Selector_2 s9800_7(wires_2450_6[0], addr_2450_6, addr_positional[39203:39200], addr_9800_7);

wire[31:0] addr_9801_7;

Selector_2 s9801_7(wires_2450_6[1], addr_2450_6, addr_positional[39207:39204], addr_9801_7);

wire[31:0] addr_9802_7;

Selector_2 s9802_7(wires_2450_6[2], addr_2450_6, addr_positional[39211:39208], addr_9802_7);

wire[31:0] addr_9803_7;

Selector_2 s9803_7(wires_2450_6[3], addr_2450_6, addr_positional[39215:39212], addr_9803_7);

wire[31:0] addr_9804_7;

Selector_2 s9804_7(wires_2451_6[0], addr_2451_6, addr_positional[39219:39216], addr_9804_7);

wire[31:0] addr_9805_7;

Selector_2 s9805_7(wires_2451_6[1], addr_2451_6, addr_positional[39223:39220], addr_9805_7);

wire[31:0] addr_9806_7;

Selector_2 s9806_7(wires_2451_6[2], addr_2451_6, addr_positional[39227:39224], addr_9806_7);

wire[31:0] addr_9807_7;

Selector_2 s9807_7(wires_2451_6[3], addr_2451_6, addr_positional[39231:39228], addr_9807_7);

wire[31:0] addr_9808_7;

Selector_2 s9808_7(wires_2452_6[0], addr_2452_6, addr_positional[39235:39232], addr_9808_7);

wire[31:0] addr_9809_7;

Selector_2 s9809_7(wires_2452_6[1], addr_2452_6, addr_positional[39239:39236], addr_9809_7);

wire[31:0] addr_9810_7;

Selector_2 s9810_7(wires_2452_6[2], addr_2452_6, addr_positional[39243:39240], addr_9810_7);

wire[31:0] addr_9811_7;

Selector_2 s9811_7(wires_2452_6[3], addr_2452_6, addr_positional[39247:39244], addr_9811_7);

wire[31:0] addr_9812_7;

Selector_2 s9812_7(wires_2453_6[0], addr_2453_6, addr_positional[39251:39248], addr_9812_7);

wire[31:0] addr_9813_7;

Selector_2 s9813_7(wires_2453_6[1], addr_2453_6, addr_positional[39255:39252], addr_9813_7);

wire[31:0] addr_9814_7;

Selector_2 s9814_7(wires_2453_6[2], addr_2453_6, addr_positional[39259:39256], addr_9814_7);

wire[31:0] addr_9815_7;

Selector_2 s9815_7(wires_2453_6[3], addr_2453_6, addr_positional[39263:39260], addr_9815_7);

wire[31:0] addr_9816_7;

Selector_2 s9816_7(wires_2454_6[0], addr_2454_6, addr_positional[39267:39264], addr_9816_7);

wire[31:0] addr_9817_7;

Selector_2 s9817_7(wires_2454_6[1], addr_2454_6, addr_positional[39271:39268], addr_9817_7);

wire[31:0] addr_9818_7;

Selector_2 s9818_7(wires_2454_6[2], addr_2454_6, addr_positional[39275:39272], addr_9818_7);

wire[31:0] addr_9819_7;

Selector_2 s9819_7(wires_2454_6[3], addr_2454_6, addr_positional[39279:39276], addr_9819_7);

wire[31:0] addr_9820_7;

Selector_2 s9820_7(wires_2455_6[0], addr_2455_6, addr_positional[39283:39280], addr_9820_7);

wire[31:0] addr_9821_7;

Selector_2 s9821_7(wires_2455_6[1], addr_2455_6, addr_positional[39287:39284], addr_9821_7);

wire[31:0] addr_9822_7;

Selector_2 s9822_7(wires_2455_6[2], addr_2455_6, addr_positional[39291:39288], addr_9822_7);

wire[31:0] addr_9823_7;

Selector_2 s9823_7(wires_2455_6[3], addr_2455_6, addr_positional[39295:39292], addr_9823_7);

wire[31:0] addr_9824_7;

Selector_2 s9824_7(wires_2456_6[0], addr_2456_6, addr_positional[39299:39296], addr_9824_7);

wire[31:0] addr_9825_7;

Selector_2 s9825_7(wires_2456_6[1], addr_2456_6, addr_positional[39303:39300], addr_9825_7);

wire[31:0] addr_9826_7;

Selector_2 s9826_7(wires_2456_6[2], addr_2456_6, addr_positional[39307:39304], addr_9826_7);

wire[31:0] addr_9827_7;

Selector_2 s9827_7(wires_2456_6[3], addr_2456_6, addr_positional[39311:39308], addr_9827_7);

wire[31:0] addr_9828_7;

Selector_2 s9828_7(wires_2457_6[0], addr_2457_6, addr_positional[39315:39312], addr_9828_7);

wire[31:0] addr_9829_7;

Selector_2 s9829_7(wires_2457_6[1], addr_2457_6, addr_positional[39319:39316], addr_9829_7);

wire[31:0] addr_9830_7;

Selector_2 s9830_7(wires_2457_6[2], addr_2457_6, addr_positional[39323:39320], addr_9830_7);

wire[31:0] addr_9831_7;

Selector_2 s9831_7(wires_2457_6[3], addr_2457_6, addr_positional[39327:39324], addr_9831_7);

wire[31:0] addr_9832_7;

Selector_2 s9832_7(wires_2458_6[0], addr_2458_6, addr_positional[39331:39328], addr_9832_7);

wire[31:0] addr_9833_7;

Selector_2 s9833_7(wires_2458_6[1], addr_2458_6, addr_positional[39335:39332], addr_9833_7);

wire[31:0] addr_9834_7;

Selector_2 s9834_7(wires_2458_6[2], addr_2458_6, addr_positional[39339:39336], addr_9834_7);

wire[31:0] addr_9835_7;

Selector_2 s9835_7(wires_2458_6[3], addr_2458_6, addr_positional[39343:39340], addr_9835_7);

wire[31:0] addr_9836_7;

Selector_2 s9836_7(wires_2459_6[0], addr_2459_6, addr_positional[39347:39344], addr_9836_7);

wire[31:0] addr_9837_7;

Selector_2 s9837_7(wires_2459_6[1], addr_2459_6, addr_positional[39351:39348], addr_9837_7);

wire[31:0] addr_9838_7;

Selector_2 s9838_7(wires_2459_6[2], addr_2459_6, addr_positional[39355:39352], addr_9838_7);

wire[31:0] addr_9839_7;

Selector_2 s9839_7(wires_2459_6[3], addr_2459_6, addr_positional[39359:39356], addr_9839_7);

wire[31:0] addr_9840_7;

Selector_2 s9840_7(wires_2460_6[0], addr_2460_6, addr_positional[39363:39360], addr_9840_7);

wire[31:0] addr_9841_7;

Selector_2 s9841_7(wires_2460_6[1], addr_2460_6, addr_positional[39367:39364], addr_9841_7);

wire[31:0] addr_9842_7;

Selector_2 s9842_7(wires_2460_6[2], addr_2460_6, addr_positional[39371:39368], addr_9842_7);

wire[31:0] addr_9843_7;

Selector_2 s9843_7(wires_2460_6[3], addr_2460_6, addr_positional[39375:39372], addr_9843_7);

wire[31:0] addr_9844_7;

Selector_2 s9844_7(wires_2461_6[0], addr_2461_6, addr_positional[39379:39376], addr_9844_7);

wire[31:0] addr_9845_7;

Selector_2 s9845_7(wires_2461_6[1], addr_2461_6, addr_positional[39383:39380], addr_9845_7);

wire[31:0] addr_9846_7;

Selector_2 s9846_7(wires_2461_6[2], addr_2461_6, addr_positional[39387:39384], addr_9846_7);

wire[31:0] addr_9847_7;

Selector_2 s9847_7(wires_2461_6[3], addr_2461_6, addr_positional[39391:39388], addr_9847_7);

wire[31:0] addr_9848_7;

Selector_2 s9848_7(wires_2462_6[0], addr_2462_6, addr_positional[39395:39392], addr_9848_7);

wire[31:0] addr_9849_7;

Selector_2 s9849_7(wires_2462_6[1], addr_2462_6, addr_positional[39399:39396], addr_9849_7);

wire[31:0] addr_9850_7;

Selector_2 s9850_7(wires_2462_6[2], addr_2462_6, addr_positional[39403:39400], addr_9850_7);

wire[31:0] addr_9851_7;

Selector_2 s9851_7(wires_2462_6[3], addr_2462_6, addr_positional[39407:39404], addr_9851_7);

wire[31:0] addr_9852_7;

Selector_2 s9852_7(wires_2463_6[0], addr_2463_6, addr_positional[39411:39408], addr_9852_7);

wire[31:0] addr_9853_7;

Selector_2 s9853_7(wires_2463_6[1], addr_2463_6, addr_positional[39415:39412], addr_9853_7);

wire[31:0] addr_9854_7;

Selector_2 s9854_7(wires_2463_6[2], addr_2463_6, addr_positional[39419:39416], addr_9854_7);

wire[31:0] addr_9855_7;

Selector_2 s9855_7(wires_2463_6[3], addr_2463_6, addr_positional[39423:39420], addr_9855_7);

wire[31:0] addr_9856_7;

Selector_2 s9856_7(wires_2464_6[0], addr_2464_6, addr_positional[39427:39424], addr_9856_7);

wire[31:0] addr_9857_7;

Selector_2 s9857_7(wires_2464_6[1], addr_2464_6, addr_positional[39431:39428], addr_9857_7);

wire[31:0] addr_9858_7;

Selector_2 s9858_7(wires_2464_6[2], addr_2464_6, addr_positional[39435:39432], addr_9858_7);

wire[31:0] addr_9859_7;

Selector_2 s9859_7(wires_2464_6[3], addr_2464_6, addr_positional[39439:39436], addr_9859_7);

wire[31:0] addr_9860_7;

Selector_2 s9860_7(wires_2465_6[0], addr_2465_6, addr_positional[39443:39440], addr_9860_7);

wire[31:0] addr_9861_7;

Selector_2 s9861_7(wires_2465_6[1], addr_2465_6, addr_positional[39447:39444], addr_9861_7);

wire[31:0] addr_9862_7;

Selector_2 s9862_7(wires_2465_6[2], addr_2465_6, addr_positional[39451:39448], addr_9862_7);

wire[31:0] addr_9863_7;

Selector_2 s9863_7(wires_2465_6[3], addr_2465_6, addr_positional[39455:39452], addr_9863_7);

wire[31:0] addr_9864_7;

Selector_2 s9864_7(wires_2466_6[0], addr_2466_6, addr_positional[39459:39456], addr_9864_7);

wire[31:0] addr_9865_7;

Selector_2 s9865_7(wires_2466_6[1], addr_2466_6, addr_positional[39463:39460], addr_9865_7);

wire[31:0] addr_9866_7;

Selector_2 s9866_7(wires_2466_6[2], addr_2466_6, addr_positional[39467:39464], addr_9866_7);

wire[31:0] addr_9867_7;

Selector_2 s9867_7(wires_2466_6[3], addr_2466_6, addr_positional[39471:39468], addr_9867_7);

wire[31:0] addr_9868_7;

Selector_2 s9868_7(wires_2467_6[0], addr_2467_6, addr_positional[39475:39472], addr_9868_7);

wire[31:0] addr_9869_7;

Selector_2 s9869_7(wires_2467_6[1], addr_2467_6, addr_positional[39479:39476], addr_9869_7);

wire[31:0] addr_9870_7;

Selector_2 s9870_7(wires_2467_6[2], addr_2467_6, addr_positional[39483:39480], addr_9870_7);

wire[31:0] addr_9871_7;

Selector_2 s9871_7(wires_2467_6[3], addr_2467_6, addr_positional[39487:39484], addr_9871_7);

wire[31:0] addr_9872_7;

Selector_2 s9872_7(wires_2468_6[0], addr_2468_6, addr_positional[39491:39488], addr_9872_7);

wire[31:0] addr_9873_7;

Selector_2 s9873_7(wires_2468_6[1], addr_2468_6, addr_positional[39495:39492], addr_9873_7);

wire[31:0] addr_9874_7;

Selector_2 s9874_7(wires_2468_6[2], addr_2468_6, addr_positional[39499:39496], addr_9874_7);

wire[31:0] addr_9875_7;

Selector_2 s9875_7(wires_2468_6[3], addr_2468_6, addr_positional[39503:39500], addr_9875_7);

wire[31:0] addr_9876_7;

Selector_2 s9876_7(wires_2469_6[0], addr_2469_6, addr_positional[39507:39504], addr_9876_7);

wire[31:0] addr_9877_7;

Selector_2 s9877_7(wires_2469_6[1], addr_2469_6, addr_positional[39511:39508], addr_9877_7);

wire[31:0] addr_9878_7;

Selector_2 s9878_7(wires_2469_6[2], addr_2469_6, addr_positional[39515:39512], addr_9878_7);

wire[31:0] addr_9879_7;

Selector_2 s9879_7(wires_2469_6[3], addr_2469_6, addr_positional[39519:39516], addr_9879_7);

wire[31:0] addr_9880_7;

Selector_2 s9880_7(wires_2470_6[0], addr_2470_6, addr_positional[39523:39520], addr_9880_7);

wire[31:0] addr_9881_7;

Selector_2 s9881_7(wires_2470_6[1], addr_2470_6, addr_positional[39527:39524], addr_9881_7);

wire[31:0] addr_9882_7;

Selector_2 s9882_7(wires_2470_6[2], addr_2470_6, addr_positional[39531:39528], addr_9882_7);

wire[31:0] addr_9883_7;

Selector_2 s9883_7(wires_2470_6[3], addr_2470_6, addr_positional[39535:39532], addr_9883_7);

wire[31:0] addr_9884_7;

Selector_2 s9884_7(wires_2471_6[0], addr_2471_6, addr_positional[39539:39536], addr_9884_7);

wire[31:0] addr_9885_7;

Selector_2 s9885_7(wires_2471_6[1], addr_2471_6, addr_positional[39543:39540], addr_9885_7);

wire[31:0] addr_9886_7;

Selector_2 s9886_7(wires_2471_6[2], addr_2471_6, addr_positional[39547:39544], addr_9886_7);

wire[31:0] addr_9887_7;

Selector_2 s9887_7(wires_2471_6[3], addr_2471_6, addr_positional[39551:39548], addr_9887_7);

wire[31:0] addr_9888_7;

Selector_2 s9888_7(wires_2472_6[0], addr_2472_6, addr_positional[39555:39552], addr_9888_7);

wire[31:0] addr_9889_7;

Selector_2 s9889_7(wires_2472_6[1], addr_2472_6, addr_positional[39559:39556], addr_9889_7);

wire[31:0] addr_9890_7;

Selector_2 s9890_7(wires_2472_6[2], addr_2472_6, addr_positional[39563:39560], addr_9890_7);

wire[31:0] addr_9891_7;

Selector_2 s9891_7(wires_2472_6[3], addr_2472_6, addr_positional[39567:39564], addr_9891_7);

wire[31:0] addr_9892_7;

Selector_2 s9892_7(wires_2473_6[0], addr_2473_6, addr_positional[39571:39568], addr_9892_7);

wire[31:0] addr_9893_7;

Selector_2 s9893_7(wires_2473_6[1], addr_2473_6, addr_positional[39575:39572], addr_9893_7);

wire[31:0] addr_9894_7;

Selector_2 s9894_7(wires_2473_6[2], addr_2473_6, addr_positional[39579:39576], addr_9894_7);

wire[31:0] addr_9895_7;

Selector_2 s9895_7(wires_2473_6[3], addr_2473_6, addr_positional[39583:39580], addr_9895_7);

wire[31:0] addr_9896_7;

Selector_2 s9896_7(wires_2474_6[0], addr_2474_6, addr_positional[39587:39584], addr_9896_7);

wire[31:0] addr_9897_7;

Selector_2 s9897_7(wires_2474_6[1], addr_2474_6, addr_positional[39591:39588], addr_9897_7);

wire[31:0] addr_9898_7;

Selector_2 s9898_7(wires_2474_6[2], addr_2474_6, addr_positional[39595:39592], addr_9898_7);

wire[31:0] addr_9899_7;

Selector_2 s9899_7(wires_2474_6[3], addr_2474_6, addr_positional[39599:39596], addr_9899_7);

wire[31:0] addr_9900_7;

Selector_2 s9900_7(wires_2475_6[0], addr_2475_6, addr_positional[39603:39600], addr_9900_7);

wire[31:0] addr_9901_7;

Selector_2 s9901_7(wires_2475_6[1], addr_2475_6, addr_positional[39607:39604], addr_9901_7);

wire[31:0] addr_9902_7;

Selector_2 s9902_7(wires_2475_6[2], addr_2475_6, addr_positional[39611:39608], addr_9902_7);

wire[31:0] addr_9903_7;

Selector_2 s9903_7(wires_2475_6[3], addr_2475_6, addr_positional[39615:39612], addr_9903_7);

wire[31:0] addr_9904_7;

Selector_2 s9904_7(wires_2476_6[0], addr_2476_6, addr_positional[39619:39616], addr_9904_7);

wire[31:0] addr_9905_7;

Selector_2 s9905_7(wires_2476_6[1], addr_2476_6, addr_positional[39623:39620], addr_9905_7);

wire[31:0] addr_9906_7;

Selector_2 s9906_7(wires_2476_6[2], addr_2476_6, addr_positional[39627:39624], addr_9906_7);

wire[31:0] addr_9907_7;

Selector_2 s9907_7(wires_2476_6[3], addr_2476_6, addr_positional[39631:39628], addr_9907_7);

wire[31:0] addr_9908_7;

Selector_2 s9908_7(wires_2477_6[0], addr_2477_6, addr_positional[39635:39632], addr_9908_7);

wire[31:0] addr_9909_7;

Selector_2 s9909_7(wires_2477_6[1], addr_2477_6, addr_positional[39639:39636], addr_9909_7);

wire[31:0] addr_9910_7;

Selector_2 s9910_7(wires_2477_6[2], addr_2477_6, addr_positional[39643:39640], addr_9910_7);

wire[31:0] addr_9911_7;

Selector_2 s9911_7(wires_2477_6[3], addr_2477_6, addr_positional[39647:39644], addr_9911_7);

wire[31:0] addr_9912_7;

Selector_2 s9912_7(wires_2478_6[0], addr_2478_6, addr_positional[39651:39648], addr_9912_7);

wire[31:0] addr_9913_7;

Selector_2 s9913_7(wires_2478_6[1], addr_2478_6, addr_positional[39655:39652], addr_9913_7);

wire[31:0] addr_9914_7;

Selector_2 s9914_7(wires_2478_6[2], addr_2478_6, addr_positional[39659:39656], addr_9914_7);

wire[31:0] addr_9915_7;

Selector_2 s9915_7(wires_2478_6[3], addr_2478_6, addr_positional[39663:39660], addr_9915_7);

wire[31:0] addr_9916_7;

Selector_2 s9916_7(wires_2479_6[0], addr_2479_6, addr_positional[39667:39664], addr_9916_7);

wire[31:0] addr_9917_7;

Selector_2 s9917_7(wires_2479_6[1], addr_2479_6, addr_positional[39671:39668], addr_9917_7);

wire[31:0] addr_9918_7;

Selector_2 s9918_7(wires_2479_6[2], addr_2479_6, addr_positional[39675:39672], addr_9918_7);

wire[31:0] addr_9919_7;

Selector_2 s9919_7(wires_2479_6[3], addr_2479_6, addr_positional[39679:39676], addr_9919_7);

wire[31:0] addr_9920_7;

Selector_2 s9920_7(wires_2480_6[0], addr_2480_6, addr_positional[39683:39680], addr_9920_7);

wire[31:0] addr_9921_7;

Selector_2 s9921_7(wires_2480_6[1], addr_2480_6, addr_positional[39687:39684], addr_9921_7);

wire[31:0] addr_9922_7;

Selector_2 s9922_7(wires_2480_6[2], addr_2480_6, addr_positional[39691:39688], addr_9922_7);

wire[31:0] addr_9923_7;

Selector_2 s9923_7(wires_2480_6[3], addr_2480_6, addr_positional[39695:39692], addr_9923_7);

wire[31:0] addr_9924_7;

Selector_2 s9924_7(wires_2481_6[0], addr_2481_6, addr_positional[39699:39696], addr_9924_7);

wire[31:0] addr_9925_7;

Selector_2 s9925_7(wires_2481_6[1], addr_2481_6, addr_positional[39703:39700], addr_9925_7);

wire[31:0] addr_9926_7;

Selector_2 s9926_7(wires_2481_6[2], addr_2481_6, addr_positional[39707:39704], addr_9926_7);

wire[31:0] addr_9927_7;

Selector_2 s9927_7(wires_2481_6[3], addr_2481_6, addr_positional[39711:39708], addr_9927_7);

wire[31:0] addr_9928_7;

Selector_2 s9928_7(wires_2482_6[0], addr_2482_6, addr_positional[39715:39712], addr_9928_7);

wire[31:0] addr_9929_7;

Selector_2 s9929_7(wires_2482_6[1], addr_2482_6, addr_positional[39719:39716], addr_9929_7);

wire[31:0] addr_9930_7;

Selector_2 s9930_7(wires_2482_6[2], addr_2482_6, addr_positional[39723:39720], addr_9930_7);

wire[31:0] addr_9931_7;

Selector_2 s9931_7(wires_2482_6[3], addr_2482_6, addr_positional[39727:39724], addr_9931_7);

wire[31:0] addr_9932_7;

Selector_2 s9932_7(wires_2483_6[0], addr_2483_6, addr_positional[39731:39728], addr_9932_7);

wire[31:0] addr_9933_7;

Selector_2 s9933_7(wires_2483_6[1], addr_2483_6, addr_positional[39735:39732], addr_9933_7);

wire[31:0] addr_9934_7;

Selector_2 s9934_7(wires_2483_6[2], addr_2483_6, addr_positional[39739:39736], addr_9934_7);

wire[31:0] addr_9935_7;

Selector_2 s9935_7(wires_2483_6[3], addr_2483_6, addr_positional[39743:39740], addr_9935_7);

wire[31:0] addr_9936_7;

Selector_2 s9936_7(wires_2484_6[0], addr_2484_6, addr_positional[39747:39744], addr_9936_7);

wire[31:0] addr_9937_7;

Selector_2 s9937_7(wires_2484_6[1], addr_2484_6, addr_positional[39751:39748], addr_9937_7);

wire[31:0] addr_9938_7;

Selector_2 s9938_7(wires_2484_6[2], addr_2484_6, addr_positional[39755:39752], addr_9938_7);

wire[31:0] addr_9939_7;

Selector_2 s9939_7(wires_2484_6[3], addr_2484_6, addr_positional[39759:39756], addr_9939_7);

wire[31:0] addr_9940_7;

Selector_2 s9940_7(wires_2485_6[0], addr_2485_6, addr_positional[39763:39760], addr_9940_7);

wire[31:0] addr_9941_7;

Selector_2 s9941_7(wires_2485_6[1], addr_2485_6, addr_positional[39767:39764], addr_9941_7);

wire[31:0] addr_9942_7;

Selector_2 s9942_7(wires_2485_6[2], addr_2485_6, addr_positional[39771:39768], addr_9942_7);

wire[31:0] addr_9943_7;

Selector_2 s9943_7(wires_2485_6[3], addr_2485_6, addr_positional[39775:39772], addr_9943_7);

wire[31:0] addr_9944_7;

Selector_2 s9944_7(wires_2486_6[0], addr_2486_6, addr_positional[39779:39776], addr_9944_7);

wire[31:0] addr_9945_7;

Selector_2 s9945_7(wires_2486_6[1], addr_2486_6, addr_positional[39783:39780], addr_9945_7);

wire[31:0] addr_9946_7;

Selector_2 s9946_7(wires_2486_6[2], addr_2486_6, addr_positional[39787:39784], addr_9946_7);

wire[31:0] addr_9947_7;

Selector_2 s9947_7(wires_2486_6[3], addr_2486_6, addr_positional[39791:39788], addr_9947_7);

wire[31:0] addr_9948_7;

Selector_2 s9948_7(wires_2487_6[0], addr_2487_6, addr_positional[39795:39792], addr_9948_7);

wire[31:0] addr_9949_7;

Selector_2 s9949_7(wires_2487_6[1], addr_2487_6, addr_positional[39799:39796], addr_9949_7);

wire[31:0] addr_9950_7;

Selector_2 s9950_7(wires_2487_6[2], addr_2487_6, addr_positional[39803:39800], addr_9950_7);

wire[31:0] addr_9951_7;

Selector_2 s9951_7(wires_2487_6[3], addr_2487_6, addr_positional[39807:39804], addr_9951_7);

wire[31:0] addr_9952_7;

Selector_2 s9952_7(wires_2488_6[0], addr_2488_6, addr_positional[39811:39808], addr_9952_7);

wire[31:0] addr_9953_7;

Selector_2 s9953_7(wires_2488_6[1], addr_2488_6, addr_positional[39815:39812], addr_9953_7);

wire[31:0] addr_9954_7;

Selector_2 s9954_7(wires_2488_6[2], addr_2488_6, addr_positional[39819:39816], addr_9954_7);

wire[31:0] addr_9955_7;

Selector_2 s9955_7(wires_2488_6[3], addr_2488_6, addr_positional[39823:39820], addr_9955_7);

wire[31:0] addr_9956_7;

Selector_2 s9956_7(wires_2489_6[0], addr_2489_6, addr_positional[39827:39824], addr_9956_7);

wire[31:0] addr_9957_7;

Selector_2 s9957_7(wires_2489_6[1], addr_2489_6, addr_positional[39831:39828], addr_9957_7);

wire[31:0] addr_9958_7;

Selector_2 s9958_7(wires_2489_6[2], addr_2489_6, addr_positional[39835:39832], addr_9958_7);

wire[31:0] addr_9959_7;

Selector_2 s9959_7(wires_2489_6[3], addr_2489_6, addr_positional[39839:39836], addr_9959_7);

wire[31:0] addr_9960_7;

Selector_2 s9960_7(wires_2490_6[0], addr_2490_6, addr_positional[39843:39840], addr_9960_7);

wire[31:0] addr_9961_7;

Selector_2 s9961_7(wires_2490_6[1], addr_2490_6, addr_positional[39847:39844], addr_9961_7);

wire[31:0] addr_9962_7;

Selector_2 s9962_7(wires_2490_6[2], addr_2490_6, addr_positional[39851:39848], addr_9962_7);

wire[31:0] addr_9963_7;

Selector_2 s9963_7(wires_2490_6[3], addr_2490_6, addr_positional[39855:39852], addr_9963_7);

wire[31:0] addr_9964_7;

Selector_2 s9964_7(wires_2491_6[0], addr_2491_6, addr_positional[39859:39856], addr_9964_7);

wire[31:0] addr_9965_7;

Selector_2 s9965_7(wires_2491_6[1], addr_2491_6, addr_positional[39863:39860], addr_9965_7);

wire[31:0] addr_9966_7;

Selector_2 s9966_7(wires_2491_6[2], addr_2491_6, addr_positional[39867:39864], addr_9966_7);

wire[31:0] addr_9967_7;

Selector_2 s9967_7(wires_2491_6[3], addr_2491_6, addr_positional[39871:39868], addr_9967_7);

wire[31:0] addr_9968_7;

Selector_2 s9968_7(wires_2492_6[0], addr_2492_6, addr_positional[39875:39872], addr_9968_7);

wire[31:0] addr_9969_7;

Selector_2 s9969_7(wires_2492_6[1], addr_2492_6, addr_positional[39879:39876], addr_9969_7);

wire[31:0] addr_9970_7;

Selector_2 s9970_7(wires_2492_6[2], addr_2492_6, addr_positional[39883:39880], addr_9970_7);

wire[31:0] addr_9971_7;

Selector_2 s9971_7(wires_2492_6[3], addr_2492_6, addr_positional[39887:39884], addr_9971_7);

wire[31:0] addr_9972_7;

Selector_2 s9972_7(wires_2493_6[0], addr_2493_6, addr_positional[39891:39888], addr_9972_7);

wire[31:0] addr_9973_7;

Selector_2 s9973_7(wires_2493_6[1], addr_2493_6, addr_positional[39895:39892], addr_9973_7);

wire[31:0] addr_9974_7;

Selector_2 s9974_7(wires_2493_6[2], addr_2493_6, addr_positional[39899:39896], addr_9974_7);

wire[31:0] addr_9975_7;

Selector_2 s9975_7(wires_2493_6[3], addr_2493_6, addr_positional[39903:39900], addr_9975_7);

wire[31:0] addr_9976_7;

Selector_2 s9976_7(wires_2494_6[0], addr_2494_6, addr_positional[39907:39904], addr_9976_7);

wire[31:0] addr_9977_7;

Selector_2 s9977_7(wires_2494_6[1], addr_2494_6, addr_positional[39911:39908], addr_9977_7);

wire[31:0] addr_9978_7;

Selector_2 s9978_7(wires_2494_6[2], addr_2494_6, addr_positional[39915:39912], addr_9978_7);

wire[31:0] addr_9979_7;

Selector_2 s9979_7(wires_2494_6[3], addr_2494_6, addr_positional[39919:39916], addr_9979_7);

wire[31:0] addr_9980_7;

Selector_2 s9980_7(wires_2495_6[0], addr_2495_6, addr_positional[39923:39920], addr_9980_7);

wire[31:0] addr_9981_7;

Selector_2 s9981_7(wires_2495_6[1], addr_2495_6, addr_positional[39927:39924], addr_9981_7);

wire[31:0] addr_9982_7;

Selector_2 s9982_7(wires_2495_6[2], addr_2495_6, addr_positional[39931:39928], addr_9982_7);

wire[31:0] addr_9983_7;

Selector_2 s9983_7(wires_2495_6[3], addr_2495_6, addr_positional[39935:39932], addr_9983_7);

wire[31:0] addr_9984_7;

Selector_2 s9984_7(wires_2496_6[0], addr_2496_6, addr_positional[39939:39936], addr_9984_7);

wire[31:0] addr_9985_7;

Selector_2 s9985_7(wires_2496_6[1], addr_2496_6, addr_positional[39943:39940], addr_9985_7);

wire[31:0] addr_9986_7;

Selector_2 s9986_7(wires_2496_6[2], addr_2496_6, addr_positional[39947:39944], addr_9986_7);

wire[31:0] addr_9987_7;

Selector_2 s9987_7(wires_2496_6[3], addr_2496_6, addr_positional[39951:39948], addr_9987_7);

wire[31:0] addr_9988_7;

Selector_2 s9988_7(wires_2497_6[0], addr_2497_6, addr_positional[39955:39952], addr_9988_7);

wire[31:0] addr_9989_7;

Selector_2 s9989_7(wires_2497_6[1], addr_2497_6, addr_positional[39959:39956], addr_9989_7);

wire[31:0] addr_9990_7;

Selector_2 s9990_7(wires_2497_6[2], addr_2497_6, addr_positional[39963:39960], addr_9990_7);

wire[31:0] addr_9991_7;

Selector_2 s9991_7(wires_2497_6[3], addr_2497_6, addr_positional[39967:39964], addr_9991_7);

wire[31:0] addr_9992_7;

Selector_2 s9992_7(wires_2498_6[0], addr_2498_6, addr_positional[39971:39968], addr_9992_7);

wire[31:0] addr_9993_7;

Selector_2 s9993_7(wires_2498_6[1], addr_2498_6, addr_positional[39975:39972], addr_9993_7);

wire[31:0] addr_9994_7;

Selector_2 s9994_7(wires_2498_6[2], addr_2498_6, addr_positional[39979:39976], addr_9994_7);

wire[31:0] addr_9995_7;

Selector_2 s9995_7(wires_2498_6[3], addr_2498_6, addr_positional[39983:39980], addr_9995_7);

wire[31:0] addr_9996_7;

Selector_2 s9996_7(wires_2499_6[0], addr_2499_6, addr_positional[39987:39984], addr_9996_7);

wire[31:0] addr_9997_7;

Selector_2 s9997_7(wires_2499_6[1], addr_2499_6, addr_positional[39991:39988], addr_9997_7);

wire[31:0] addr_9998_7;

Selector_2 s9998_7(wires_2499_6[2], addr_2499_6, addr_positional[39995:39992], addr_9998_7);

wire[31:0] addr_9999_7;

Selector_2 s9999_7(wires_2499_6[3], addr_2499_6, addr_positional[39999:39996], addr_9999_7);

wire[31:0] addr_10000_7;

Selector_2 s10000_7(wires_2500_6[0], addr_2500_6, addr_positional[40003:40000], addr_10000_7);

wire[31:0] addr_10001_7;

Selector_2 s10001_7(wires_2500_6[1], addr_2500_6, addr_positional[40007:40004], addr_10001_7);

wire[31:0] addr_10002_7;

Selector_2 s10002_7(wires_2500_6[2], addr_2500_6, addr_positional[40011:40008], addr_10002_7);

wire[31:0] addr_10003_7;

Selector_2 s10003_7(wires_2500_6[3], addr_2500_6, addr_positional[40015:40012], addr_10003_7);

wire[31:0] addr_10004_7;

Selector_2 s10004_7(wires_2501_6[0], addr_2501_6, addr_positional[40019:40016], addr_10004_7);

wire[31:0] addr_10005_7;

Selector_2 s10005_7(wires_2501_6[1], addr_2501_6, addr_positional[40023:40020], addr_10005_7);

wire[31:0] addr_10006_7;

Selector_2 s10006_7(wires_2501_6[2], addr_2501_6, addr_positional[40027:40024], addr_10006_7);

wire[31:0] addr_10007_7;

Selector_2 s10007_7(wires_2501_6[3], addr_2501_6, addr_positional[40031:40028], addr_10007_7);

wire[31:0] addr_10008_7;

Selector_2 s10008_7(wires_2502_6[0], addr_2502_6, addr_positional[40035:40032], addr_10008_7);

wire[31:0] addr_10009_7;

Selector_2 s10009_7(wires_2502_6[1], addr_2502_6, addr_positional[40039:40036], addr_10009_7);

wire[31:0] addr_10010_7;

Selector_2 s10010_7(wires_2502_6[2], addr_2502_6, addr_positional[40043:40040], addr_10010_7);

wire[31:0] addr_10011_7;

Selector_2 s10011_7(wires_2502_6[3], addr_2502_6, addr_positional[40047:40044], addr_10011_7);

wire[31:0] addr_10012_7;

Selector_2 s10012_7(wires_2503_6[0], addr_2503_6, addr_positional[40051:40048], addr_10012_7);

wire[31:0] addr_10013_7;

Selector_2 s10013_7(wires_2503_6[1], addr_2503_6, addr_positional[40055:40052], addr_10013_7);

wire[31:0] addr_10014_7;

Selector_2 s10014_7(wires_2503_6[2], addr_2503_6, addr_positional[40059:40056], addr_10014_7);

wire[31:0] addr_10015_7;

Selector_2 s10015_7(wires_2503_6[3], addr_2503_6, addr_positional[40063:40060], addr_10015_7);

wire[31:0] addr_10016_7;

Selector_2 s10016_7(wires_2504_6[0], addr_2504_6, addr_positional[40067:40064], addr_10016_7);

wire[31:0] addr_10017_7;

Selector_2 s10017_7(wires_2504_6[1], addr_2504_6, addr_positional[40071:40068], addr_10017_7);

wire[31:0] addr_10018_7;

Selector_2 s10018_7(wires_2504_6[2], addr_2504_6, addr_positional[40075:40072], addr_10018_7);

wire[31:0] addr_10019_7;

Selector_2 s10019_7(wires_2504_6[3], addr_2504_6, addr_positional[40079:40076], addr_10019_7);

wire[31:0] addr_10020_7;

Selector_2 s10020_7(wires_2505_6[0], addr_2505_6, addr_positional[40083:40080], addr_10020_7);

wire[31:0] addr_10021_7;

Selector_2 s10021_7(wires_2505_6[1], addr_2505_6, addr_positional[40087:40084], addr_10021_7);

wire[31:0] addr_10022_7;

Selector_2 s10022_7(wires_2505_6[2], addr_2505_6, addr_positional[40091:40088], addr_10022_7);

wire[31:0] addr_10023_7;

Selector_2 s10023_7(wires_2505_6[3], addr_2505_6, addr_positional[40095:40092], addr_10023_7);

wire[31:0] addr_10024_7;

Selector_2 s10024_7(wires_2506_6[0], addr_2506_6, addr_positional[40099:40096], addr_10024_7);

wire[31:0] addr_10025_7;

Selector_2 s10025_7(wires_2506_6[1], addr_2506_6, addr_positional[40103:40100], addr_10025_7);

wire[31:0] addr_10026_7;

Selector_2 s10026_7(wires_2506_6[2], addr_2506_6, addr_positional[40107:40104], addr_10026_7);

wire[31:0] addr_10027_7;

Selector_2 s10027_7(wires_2506_6[3], addr_2506_6, addr_positional[40111:40108], addr_10027_7);

wire[31:0] addr_10028_7;

Selector_2 s10028_7(wires_2507_6[0], addr_2507_6, addr_positional[40115:40112], addr_10028_7);

wire[31:0] addr_10029_7;

Selector_2 s10029_7(wires_2507_6[1], addr_2507_6, addr_positional[40119:40116], addr_10029_7);

wire[31:0] addr_10030_7;

Selector_2 s10030_7(wires_2507_6[2], addr_2507_6, addr_positional[40123:40120], addr_10030_7);

wire[31:0] addr_10031_7;

Selector_2 s10031_7(wires_2507_6[3], addr_2507_6, addr_positional[40127:40124], addr_10031_7);

wire[31:0] addr_10032_7;

Selector_2 s10032_7(wires_2508_6[0], addr_2508_6, addr_positional[40131:40128], addr_10032_7);

wire[31:0] addr_10033_7;

Selector_2 s10033_7(wires_2508_6[1], addr_2508_6, addr_positional[40135:40132], addr_10033_7);

wire[31:0] addr_10034_7;

Selector_2 s10034_7(wires_2508_6[2], addr_2508_6, addr_positional[40139:40136], addr_10034_7);

wire[31:0] addr_10035_7;

Selector_2 s10035_7(wires_2508_6[3], addr_2508_6, addr_positional[40143:40140], addr_10035_7);

wire[31:0] addr_10036_7;

Selector_2 s10036_7(wires_2509_6[0], addr_2509_6, addr_positional[40147:40144], addr_10036_7);

wire[31:0] addr_10037_7;

Selector_2 s10037_7(wires_2509_6[1], addr_2509_6, addr_positional[40151:40148], addr_10037_7);

wire[31:0] addr_10038_7;

Selector_2 s10038_7(wires_2509_6[2], addr_2509_6, addr_positional[40155:40152], addr_10038_7);

wire[31:0] addr_10039_7;

Selector_2 s10039_7(wires_2509_6[3], addr_2509_6, addr_positional[40159:40156], addr_10039_7);

wire[31:0] addr_10040_7;

Selector_2 s10040_7(wires_2510_6[0], addr_2510_6, addr_positional[40163:40160], addr_10040_7);

wire[31:0] addr_10041_7;

Selector_2 s10041_7(wires_2510_6[1], addr_2510_6, addr_positional[40167:40164], addr_10041_7);

wire[31:0] addr_10042_7;

Selector_2 s10042_7(wires_2510_6[2], addr_2510_6, addr_positional[40171:40168], addr_10042_7);

wire[31:0] addr_10043_7;

Selector_2 s10043_7(wires_2510_6[3], addr_2510_6, addr_positional[40175:40172], addr_10043_7);

wire[31:0] addr_10044_7;

Selector_2 s10044_7(wires_2511_6[0], addr_2511_6, addr_positional[40179:40176], addr_10044_7);

wire[31:0] addr_10045_7;

Selector_2 s10045_7(wires_2511_6[1], addr_2511_6, addr_positional[40183:40180], addr_10045_7);

wire[31:0] addr_10046_7;

Selector_2 s10046_7(wires_2511_6[2], addr_2511_6, addr_positional[40187:40184], addr_10046_7);

wire[31:0] addr_10047_7;

Selector_2 s10047_7(wires_2511_6[3], addr_2511_6, addr_positional[40191:40188], addr_10047_7);

wire[31:0] addr_10048_7;

Selector_2 s10048_7(wires_2512_6[0], addr_2512_6, addr_positional[40195:40192], addr_10048_7);

wire[31:0] addr_10049_7;

Selector_2 s10049_7(wires_2512_6[1], addr_2512_6, addr_positional[40199:40196], addr_10049_7);

wire[31:0] addr_10050_7;

Selector_2 s10050_7(wires_2512_6[2], addr_2512_6, addr_positional[40203:40200], addr_10050_7);

wire[31:0] addr_10051_7;

Selector_2 s10051_7(wires_2512_6[3], addr_2512_6, addr_positional[40207:40204], addr_10051_7);

wire[31:0] addr_10052_7;

Selector_2 s10052_7(wires_2513_6[0], addr_2513_6, addr_positional[40211:40208], addr_10052_7);

wire[31:0] addr_10053_7;

Selector_2 s10053_7(wires_2513_6[1], addr_2513_6, addr_positional[40215:40212], addr_10053_7);

wire[31:0] addr_10054_7;

Selector_2 s10054_7(wires_2513_6[2], addr_2513_6, addr_positional[40219:40216], addr_10054_7);

wire[31:0] addr_10055_7;

Selector_2 s10055_7(wires_2513_6[3], addr_2513_6, addr_positional[40223:40220], addr_10055_7);

wire[31:0] addr_10056_7;

Selector_2 s10056_7(wires_2514_6[0], addr_2514_6, addr_positional[40227:40224], addr_10056_7);

wire[31:0] addr_10057_7;

Selector_2 s10057_7(wires_2514_6[1], addr_2514_6, addr_positional[40231:40228], addr_10057_7);

wire[31:0] addr_10058_7;

Selector_2 s10058_7(wires_2514_6[2], addr_2514_6, addr_positional[40235:40232], addr_10058_7);

wire[31:0] addr_10059_7;

Selector_2 s10059_7(wires_2514_6[3], addr_2514_6, addr_positional[40239:40236], addr_10059_7);

wire[31:0] addr_10060_7;

Selector_2 s10060_7(wires_2515_6[0], addr_2515_6, addr_positional[40243:40240], addr_10060_7);

wire[31:0] addr_10061_7;

Selector_2 s10061_7(wires_2515_6[1], addr_2515_6, addr_positional[40247:40244], addr_10061_7);

wire[31:0] addr_10062_7;

Selector_2 s10062_7(wires_2515_6[2], addr_2515_6, addr_positional[40251:40248], addr_10062_7);

wire[31:0] addr_10063_7;

Selector_2 s10063_7(wires_2515_6[3], addr_2515_6, addr_positional[40255:40252], addr_10063_7);

wire[31:0] addr_10064_7;

Selector_2 s10064_7(wires_2516_6[0], addr_2516_6, addr_positional[40259:40256], addr_10064_7);

wire[31:0] addr_10065_7;

Selector_2 s10065_7(wires_2516_6[1], addr_2516_6, addr_positional[40263:40260], addr_10065_7);

wire[31:0] addr_10066_7;

Selector_2 s10066_7(wires_2516_6[2], addr_2516_6, addr_positional[40267:40264], addr_10066_7);

wire[31:0] addr_10067_7;

Selector_2 s10067_7(wires_2516_6[3], addr_2516_6, addr_positional[40271:40268], addr_10067_7);

wire[31:0] addr_10068_7;

Selector_2 s10068_7(wires_2517_6[0], addr_2517_6, addr_positional[40275:40272], addr_10068_7);

wire[31:0] addr_10069_7;

Selector_2 s10069_7(wires_2517_6[1], addr_2517_6, addr_positional[40279:40276], addr_10069_7);

wire[31:0] addr_10070_7;

Selector_2 s10070_7(wires_2517_6[2], addr_2517_6, addr_positional[40283:40280], addr_10070_7);

wire[31:0] addr_10071_7;

Selector_2 s10071_7(wires_2517_6[3], addr_2517_6, addr_positional[40287:40284], addr_10071_7);

wire[31:0] addr_10072_7;

Selector_2 s10072_7(wires_2518_6[0], addr_2518_6, addr_positional[40291:40288], addr_10072_7);

wire[31:0] addr_10073_7;

Selector_2 s10073_7(wires_2518_6[1], addr_2518_6, addr_positional[40295:40292], addr_10073_7);

wire[31:0] addr_10074_7;

Selector_2 s10074_7(wires_2518_6[2], addr_2518_6, addr_positional[40299:40296], addr_10074_7);

wire[31:0] addr_10075_7;

Selector_2 s10075_7(wires_2518_6[3], addr_2518_6, addr_positional[40303:40300], addr_10075_7);

wire[31:0] addr_10076_7;

Selector_2 s10076_7(wires_2519_6[0], addr_2519_6, addr_positional[40307:40304], addr_10076_7);

wire[31:0] addr_10077_7;

Selector_2 s10077_7(wires_2519_6[1], addr_2519_6, addr_positional[40311:40308], addr_10077_7);

wire[31:0] addr_10078_7;

Selector_2 s10078_7(wires_2519_6[2], addr_2519_6, addr_positional[40315:40312], addr_10078_7);

wire[31:0] addr_10079_7;

Selector_2 s10079_7(wires_2519_6[3], addr_2519_6, addr_positional[40319:40316], addr_10079_7);

wire[31:0] addr_10080_7;

Selector_2 s10080_7(wires_2520_6[0], addr_2520_6, addr_positional[40323:40320], addr_10080_7);

wire[31:0] addr_10081_7;

Selector_2 s10081_7(wires_2520_6[1], addr_2520_6, addr_positional[40327:40324], addr_10081_7);

wire[31:0] addr_10082_7;

Selector_2 s10082_7(wires_2520_6[2], addr_2520_6, addr_positional[40331:40328], addr_10082_7);

wire[31:0] addr_10083_7;

Selector_2 s10083_7(wires_2520_6[3], addr_2520_6, addr_positional[40335:40332], addr_10083_7);

wire[31:0] addr_10084_7;

Selector_2 s10084_7(wires_2521_6[0], addr_2521_6, addr_positional[40339:40336], addr_10084_7);

wire[31:0] addr_10085_7;

Selector_2 s10085_7(wires_2521_6[1], addr_2521_6, addr_positional[40343:40340], addr_10085_7);

wire[31:0] addr_10086_7;

Selector_2 s10086_7(wires_2521_6[2], addr_2521_6, addr_positional[40347:40344], addr_10086_7);

wire[31:0] addr_10087_7;

Selector_2 s10087_7(wires_2521_6[3], addr_2521_6, addr_positional[40351:40348], addr_10087_7);

wire[31:0] addr_10088_7;

Selector_2 s10088_7(wires_2522_6[0], addr_2522_6, addr_positional[40355:40352], addr_10088_7);

wire[31:0] addr_10089_7;

Selector_2 s10089_7(wires_2522_6[1], addr_2522_6, addr_positional[40359:40356], addr_10089_7);

wire[31:0] addr_10090_7;

Selector_2 s10090_7(wires_2522_6[2], addr_2522_6, addr_positional[40363:40360], addr_10090_7);

wire[31:0] addr_10091_7;

Selector_2 s10091_7(wires_2522_6[3], addr_2522_6, addr_positional[40367:40364], addr_10091_7);

wire[31:0] addr_10092_7;

Selector_2 s10092_7(wires_2523_6[0], addr_2523_6, addr_positional[40371:40368], addr_10092_7);

wire[31:0] addr_10093_7;

Selector_2 s10093_7(wires_2523_6[1], addr_2523_6, addr_positional[40375:40372], addr_10093_7);

wire[31:0] addr_10094_7;

Selector_2 s10094_7(wires_2523_6[2], addr_2523_6, addr_positional[40379:40376], addr_10094_7);

wire[31:0] addr_10095_7;

Selector_2 s10095_7(wires_2523_6[3], addr_2523_6, addr_positional[40383:40380], addr_10095_7);

wire[31:0] addr_10096_7;

Selector_2 s10096_7(wires_2524_6[0], addr_2524_6, addr_positional[40387:40384], addr_10096_7);

wire[31:0] addr_10097_7;

Selector_2 s10097_7(wires_2524_6[1], addr_2524_6, addr_positional[40391:40388], addr_10097_7);

wire[31:0] addr_10098_7;

Selector_2 s10098_7(wires_2524_6[2], addr_2524_6, addr_positional[40395:40392], addr_10098_7);

wire[31:0] addr_10099_7;

Selector_2 s10099_7(wires_2524_6[3], addr_2524_6, addr_positional[40399:40396], addr_10099_7);

wire[31:0] addr_10100_7;

Selector_2 s10100_7(wires_2525_6[0], addr_2525_6, addr_positional[40403:40400], addr_10100_7);

wire[31:0] addr_10101_7;

Selector_2 s10101_7(wires_2525_6[1], addr_2525_6, addr_positional[40407:40404], addr_10101_7);

wire[31:0] addr_10102_7;

Selector_2 s10102_7(wires_2525_6[2], addr_2525_6, addr_positional[40411:40408], addr_10102_7);

wire[31:0] addr_10103_7;

Selector_2 s10103_7(wires_2525_6[3], addr_2525_6, addr_positional[40415:40412], addr_10103_7);

wire[31:0] addr_10104_7;

Selector_2 s10104_7(wires_2526_6[0], addr_2526_6, addr_positional[40419:40416], addr_10104_7);

wire[31:0] addr_10105_7;

Selector_2 s10105_7(wires_2526_6[1], addr_2526_6, addr_positional[40423:40420], addr_10105_7);

wire[31:0] addr_10106_7;

Selector_2 s10106_7(wires_2526_6[2], addr_2526_6, addr_positional[40427:40424], addr_10106_7);

wire[31:0] addr_10107_7;

Selector_2 s10107_7(wires_2526_6[3], addr_2526_6, addr_positional[40431:40428], addr_10107_7);

wire[31:0] addr_10108_7;

Selector_2 s10108_7(wires_2527_6[0], addr_2527_6, addr_positional[40435:40432], addr_10108_7);

wire[31:0] addr_10109_7;

Selector_2 s10109_7(wires_2527_6[1], addr_2527_6, addr_positional[40439:40436], addr_10109_7);

wire[31:0] addr_10110_7;

Selector_2 s10110_7(wires_2527_6[2], addr_2527_6, addr_positional[40443:40440], addr_10110_7);

wire[31:0] addr_10111_7;

Selector_2 s10111_7(wires_2527_6[3], addr_2527_6, addr_positional[40447:40444], addr_10111_7);

wire[31:0] addr_10112_7;

Selector_2 s10112_7(wires_2528_6[0], addr_2528_6, addr_positional[40451:40448], addr_10112_7);

wire[31:0] addr_10113_7;

Selector_2 s10113_7(wires_2528_6[1], addr_2528_6, addr_positional[40455:40452], addr_10113_7);

wire[31:0] addr_10114_7;

Selector_2 s10114_7(wires_2528_6[2], addr_2528_6, addr_positional[40459:40456], addr_10114_7);

wire[31:0] addr_10115_7;

Selector_2 s10115_7(wires_2528_6[3], addr_2528_6, addr_positional[40463:40460], addr_10115_7);

wire[31:0] addr_10116_7;

Selector_2 s10116_7(wires_2529_6[0], addr_2529_6, addr_positional[40467:40464], addr_10116_7);

wire[31:0] addr_10117_7;

Selector_2 s10117_7(wires_2529_6[1], addr_2529_6, addr_positional[40471:40468], addr_10117_7);

wire[31:0] addr_10118_7;

Selector_2 s10118_7(wires_2529_6[2], addr_2529_6, addr_positional[40475:40472], addr_10118_7);

wire[31:0] addr_10119_7;

Selector_2 s10119_7(wires_2529_6[3], addr_2529_6, addr_positional[40479:40476], addr_10119_7);

wire[31:0] addr_10120_7;

Selector_2 s10120_7(wires_2530_6[0], addr_2530_6, addr_positional[40483:40480], addr_10120_7);

wire[31:0] addr_10121_7;

Selector_2 s10121_7(wires_2530_6[1], addr_2530_6, addr_positional[40487:40484], addr_10121_7);

wire[31:0] addr_10122_7;

Selector_2 s10122_7(wires_2530_6[2], addr_2530_6, addr_positional[40491:40488], addr_10122_7);

wire[31:0] addr_10123_7;

Selector_2 s10123_7(wires_2530_6[3], addr_2530_6, addr_positional[40495:40492], addr_10123_7);

wire[31:0] addr_10124_7;

Selector_2 s10124_7(wires_2531_6[0], addr_2531_6, addr_positional[40499:40496], addr_10124_7);

wire[31:0] addr_10125_7;

Selector_2 s10125_7(wires_2531_6[1], addr_2531_6, addr_positional[40503:40500], addr_10125_7);

wire[31:0] addr_10126_7;

Selector_2 s10126_7(wires_2531_6[2], addr_2531_6, addr_positional[40507:40504], addr_10126_7);

wire[31:0] addr_10127_7;

Selector_2 s10127_7(wires_2531_6[3], addr_2531_6, addr_positional[40511:40508], addr_10127_7);

wire[31:0] addr_10128_7;

Selector_2 s10128_7(wires_2532_6[0], addr_2532_6, addr_positional[40515:40512], addr_10128_7);

wire[31:0] addr_10129_7;

Selector_2 s10129_7(wires_2532_6[1], addr_2532_6, addr_positional[40519:40516], addr_10129_7);

wire[31:0] addr_10130_7;

Selector_2 s10130_7(wires_2532_6[2], addr_2532_6, addr_positional[40523:40520], addr_10130_7);

wire[31:0] addr_10131_7;

Selector_2 s10131_7(wires_2532_6[3], addr_2532_6, addr_positional[40527:40524], addr_10131_7);

wire[31:0] addr_10132_7;

Selector_2 s10132_7(wires_2533_6[0], addr_2533_6, addr_positional[40531:40528], addr_10132_7);

wire[31:0] addr_10133_7;

Selector_2 s10133_7(wires_2533_6[1], addr_2533_6, addr_positional[40535:40532], addr_10133_7);

wire[31:0] addr_10134_7;

Selector_2 s10134_7(wires_2533_6[2], addr_2533_6, addr_positional[40539:40536], addr_10134_7);

wire[31:0] addr_10135_7;

Selector_2 s10135_7(wires_2533_6[3], addr_2533_6, addr_positional[40543:40540], addr_10135_7);

wire[31:0] addr_10136_7;

Selector_2 s10136_7(wires_2534_6[0], addr_2534_6, addr_positional[40547:40544], addr_10136_7);

wire[31:0] addr_10137_7;

Selector_2 s10137_7(wires_2534_6[1], addr_2534_6, addr_positional[40551:40548], addr_10137_7);

wire[31:0] addr_10138_7;

Selector_2 s10138_7(wires_2534_6[2], addr_2534_6, addr_positional[40555:40552], addr_10138_7);

wire[31:0] addr_10139_7;

Selector_2 s10139_7(wires_2534_6[3], addr_2534_6, addr_positional[40559:40556], addr_10139_7);

wire[31:0] addr_10140_7;

Selector_2 s10140_7(wires_2535_6[0], addr_2535_6, addr_positional[40563:40560], addr_10140_7);

wire[31:0] addr_10141_7;

Selector_2 s10141_7(wires_2535_6[1], addr_2535_6, addr_positional[40567:40564], addr_10141_7);

wire[31:0] addr_10142_7;

Selector_2 s10142_7(wires_2535_6[2], addr_2535_6, addr_positional[40571:40568], addr_10142_7);

wire[31:0] addr_10143_7;

Selector_2 s10143_7(wires_2535_6[3], addr_2535_6, addr_positional[40575:40572], addr_10143_7);

wire[31:0] addr_10144_7;

Selector_2 s10144_7(wires_2536_6[0], addr_2536_6, addr_positional[40579:40576], addr_10144_7);

wire[31:0] addr_10145_7;

Selector_2 s10145_7(wires_2536_6[1], addr_2536_6, addr_positional[40583:40580], addr_10145_7);

wire[31:0] addr_10146_7;

Selector_2 s10146_7(wires_2536_6[2], addr_2536_6, addr_positional[40587:40584], addr_10146_7);

wire[31:0] addr_10147_7;

Selector_2 s10147_7(wires_2536_6[3], addr_2536_6, addr_positional[40591:40588], addr_10147_7);

wire[31:0] addr_10148_7;

Selector_2 s10148_7(wires_2537_6[0], addr_2537_6, addr_positional[40595:40592], addr_10148_7);

wire[31:0] addr_10149_7;

Selector_2 s10149_7(wires_2537_6[1], addr_2537_6, addr_positional[40599:40596], addr_10149_7);

wire[31:0] addr_10150_7;

Selector_2 s10150_7(wires_2537_6[2], addr_2537_6, addr_positional[40603:40600], addr_10150_7);

wire[31:0] addr_10151_7;

Selector_2 s10151_7(wires_2537_6[3], addr_2537_6, addr_positional[40607:40604], addr_10151_7);

wire[31:0] addr_10152_7;

Selector_2 s10152_7(wires_2538_6[0], addr_2538_6, addr_positional[40611:40608], addr_10152_7);

wire[31:0] addr_10153_7;

Selector_2 s10153_7(wires_2538_6[1], addr_2538_6, addr_positional[40615:40612], addr_10153_7);

wire[31:0] addr_10154_7;

Selector_2 s10154_7(wires_2538_6[2], addr_2538_6, addr_positional[40619:40616], addr_10154_7);

wire[31:0] addr_10155_7;

Selector_2 s10155_7(wires_2538_6[3], addr_2538_6, addr_positional[40623:40620], addr_10155_7);

wire[31:0] addr_10156_7;

Selector_2 s10156_7(wires_2539_6[0], addr_2539_6, addr_positional[40627:40624], addr_10156_7);

wire[31:0] addr_10157_7;

Selector_2 s10157_7(wires_2539_6[1], addr_2539_6, addr_positional[40631:40628], addr_10157_7);

wire[31:0] addr_10158_7;

Selector_2 s10158_7(wires_2539_6[2], addr_2539_6, addr_positional[40635:40632], addr_10158_7);

wire[31:0] addr_10159_7;

Selector_2 s10159_7(wires_2539_6[3], addr_2539_6, addr_positional[40639:40636], addr_10159_7);

wire[31:0] addr_10160_7;

Selector_2 s10160_7(wires_2540_6[0], addr_2540_6, addr_positional[40643:40640], addr_10160_7);

wire[31:0] addr_10161_7;

Selector_2 s10161_7(wires_2540_6[1], addr_2540_6, addr_positional[40647:40644], addr_10161_7);

wire[31:0] addr_10162_7;

Selector_2 s10162_7(wires_2540_6[2], addr_2540_6, addr_positional[40651:40648], addr_10162_7);

wire[31:0] addr_10163_7;

Selector_2 s10163_7(wires_2540_6[3], addr_2540_6, addr_positional[40655:40652], addr_10163_7);

wire[31:0] addr_10164_7;

Selector_2 s10164_7(wires_2541_6[0], addr_2541_6, addr_positional[40659:40656], addr_10164_7);

wire[31:0] addr_10165_7;

Selector_2 s10165_7(wires_2541_6[1], addr_2541_6, addr_positional[40663:40660], addr_10165_7);

wire[31:0] addr_10166_7;

Selector_2 s10166_7(wires_2541_6[2], addr_2541_6, addr_positional[40667:40664], addr_10166_7);

wire[31:0] addr_10167_7;

Selector_2 s10167_7(wires_2541_6[3], addr_2541_6, addr_positional[40671:40668], addr_10167_7);

wire[31:0] addr_10168_7;

Selector_2 s10168_7(wires_2542_6[0], addr_2542_6, addr_positional[40675:40672], addr_10168_7);

wire[31:0] addr_10169_7;

Selector_2 s10169_7(wires_2542_6[1], addr_2542_6, addr_positional[40679:40676], addr_10169_7);

wire[31:0] addr_10170_7;

Selector_2 s10170_7(wires_2542_6[2], addr_2542_6, addr_positional[40683:40680], addr_10170_7);

wire[31:0] addr_10171_7;

Selector_2 s10171_7(wires_2542_6[3], addr_2542_6, addr_positional[40687:40684], addr_10171_7);

wire[31:0] addr_10172_7;

Selector_2 s10172_7(wires_2543_6[0], addr_2543_6, addr_positional[40691:40688], addr_10172_7);

wire[31:0] addr_10173_7;

Selector_2 s10173_7(wires_2543_6[1], addr_2543_6, addr_positional[40695:40692], addr_10173_7);

wire[31:0] addr_10174_7;

Selector_2 s10174_7(wires_2543_6[2], addr_2543_6, addr_positional[40699:40696], addr_10174_7);

wire[31:0] addr_10175_7;

Selector_2 s10175_7(wires_2543_6[3], addr_2543_6, addr_positional[40703:40700], addr_10175_7);

wire[31:0] addr_10176_7;

Selector_2 s10176_7(wires_2544_6[0], addr_2544_6, addr_positional[40707:40704], addr_10176_7);

wire[31:0] addr_10177_7;

Selector_2 s10177_7(wires_2544_6[1], addr_2544_6, addr_positional[40711:40708], addr_10177_7);

wire[31:0] addr_10178_7;

Selector_2 s10178_7(wires_2544_6[2], addr_2544_6, addr_positional[40715:40712], addr_10178_7);

wire[31:0] addr_10179_7;

Selector_2 s10179_7(wires_2544_6[3], addr_2544_6, addr_positional[40719:40716], addr_10179_7);

wire[31:0] addr_10180_7;

Selector_2 s10180_7(wires_2545_6[0], addr_2545_6, addr_positional[40723:40720], addr_10180_7);

wire[31:0] addr_10181_7;

Selector_2 s10181_7(wires_2545_6[1], addr_2545_6, addr_positional[40727:40724], addr_10181_7);

wire[31:0] addr_10182_7;

Selector_2 s10182_7(wires_2545_6[2], addr_2545_6, addr_positional[40731:40728], addr_10182_7);

wire[31:0] addr_10183_7;

Selector_2 s10183_7(wires_2545_6[3], addr_2545_6, addr_positional[40735:40732], addr_10183_7);

wire[31:0] addr_10184_7;

Selector_2 s10184_7(wires_2546_6[0], addr_2546_6, addr_positional[40739:40736], addr_10184_7);

wire[31:0] addr_10185_7;

Selector_2 s10185_7(wires_2546_6[1], addr_2546_6, addr_positional[40743:40740], addr_10185_7);

wire[31:0] addr_10186_7;

Selector_2 s10186_7(wires_2546_6[2], addr_2546_6, addr_positional[40747:40744], addr_10186_7);

wire[31:0] addr_10187_7;

Selector_2 s10187_7(wires_2546_6[3], addr_2546_6, addr_positional[40751:40748], addr_10187_7);

wire[31:0] addr_10188_7;

Selector_2 s10188_7(wires_2547_6[0], addr_2547_6, addr_positional[40755:40752], addr_10188_7);

wire[31:0] addr_10189_7;

Selector_2 s10189_7(wires_2547_6[1], addr_2547_6, addr_positional[40759:40756], addr_10189_7);

wire[31:0] addr_10190_7;

Selector_2 s10190_7(wires_2547_6[2], addr_2547_6, addr_positional[40763:40760], addr_10190_7);

wire[31:0] addr_10191_7;

Selector_2 s10191_7(wires_2547_6[3], addr_2547_6, addr_positional[40767:40764], addr_10191_7);

wire[31:0] addr_10192_7;

Selector_2 s10192_7(wires_2548_6[0], addr_2548_6, addr_positional[40771:40768], addr_10192_7);

wire[31:0] addr_10193_7;

Selector_2 s10193_7(wires_2548_6[1], addr_2548_6, addr_positional[40775:40772], addr_10193_7);

wire[31:0] addr_10194_7;

Selector_2 s10194_7(wires_2548_6[2], addr_2548_6, addr_positional[40779:40776], addr_10194_7);

wire[31:0] addr_10195_7;

Selector_2 s10195_7(wires_2548_6[3], addr_2548_6, addr_positional[40783:40780], addr_10195_7);

wire[31:0] addr_10196_7;

Selector_2 s10196_7(wires_2549_6[0], addr_2549_6, addr_positional[40787:40784], addr_10196_7);

wire[31:0] addr_10197_7;

Selector_2 s10197_7(wires_2549_6[1], addr_2549_6, addr_positional[40791:40788], addr_10197_7);

wire[31:0] addr_10198_7;

Selector_2 s10198_7(wires_2549_6[2], addr_2549_6, addr_positional[40795:40792], addr_10198_7);

wire[31:0] addr_10199_7;

Selector_2 s10199_7(wires_2549_6[3], addr_2549_6, addr_positional[40799:40796], addr_10199_7);

wire[31:0] addr_10200_7;

Selector_2 s10200_7(wires_2550_6[0], addr_2550_6, addr_positional[40803:40800], addr_10200_7);

wire[31:0] addr_10201_7;

Selector_2 s10201_7(wires_2550_6[1], addr_2550_6, addr_positional[40807:40804], addr_10201_7);

wire[31:0] addr_10202_7;

Selector_2 s10202_7(wires_2550_6[2], addr_2550_6, addr_positional[40811:40808], addr_10202_7);

wire[31:0] addr_10203_7;

Selector_2 s10203_7(wires_2550_6[3], addr_2550_6, addr_positional[40815:40812], addr_10203_7);

wire[31:0] addr_10204_7;

Selector_2 s10204_7(wires_2551_6[0], addr_2551_6, addr_positional[40819:40816], addr_10204_7);

wire[31:0] addr_10205_7;

Selector_2 s10205_7(wires_2551_6[1], addr_2551_6, addr_positional[40823:40820], addr_10205_7);

wire[31:0] addr_10206_7;

Selector_2 s10206_7(wires_2551_6[2], addr_2551_6, addr_positional[40827:40824], addr_10206_7);

wire[31:0] addr_10207_7;

Selector_2 s10207_7(wires_2551_6[3], addr_2551_6, addr_positional[40831:40828], addr_10207_7);

wire[31:0] addr_10208_7;

Selector_2 s10208_7(wires_2552_6[0], addr_2552_6, addr_positional[40835:40832], addr_10208_7);

wire[31:0] addr_10209_7;

Selector_2 s10209_7(wires_2552_6[1], addr_2552_6, addr_positional[40839:40836], addr_10209_7);

wire[31:0] addr_10210_7;

Selector_2 s10210_7(wires_2552_6[2], addr_2552_6, addr_positional[40843:40840], addr_10210_7);

wire[31:0] addr_10211_7;

Selector_2 s10211_7(wires_2552_6[3], addr_2552_6, addr_positional[40847:40844], addr_10211_7);

wire[31:0] addr_10212_7;

Selector_2 s10212_7(wires_2553_6[0], addr_2553_6, addr_positional[40851:40848], addr_10212_7);

wire[31:0] addr_10213_7;

Selector_2 s10213_7(wires_2553_6[1], addr_2553_6, addr_positional[40855:40852], addr_10213_7);

wire[31:0] addr_10214_7;

Selector_2 s10214_7(wires_2553_6[2], addr_2553_6, addr_positional[40859:40856], addr_10214_7);

wire[31:0] addr_10215_7;

Selector_2 s10215_7(wires_2553_6[3], addr_2553_6, addr_positional[40863:40860], addr_10215_7);

wire[31:0] addr_10216_7;

Selector_2 s10216_7(wires_2554_6[0], addr_2554_6, addr_positional[40867:40864], addr_10216_7);

wire[31:0] addr_10217_7;

Selector_2 s10217_7(wires_2554_6[1], addr_2554_6, addr_positional[40871:40868], addr_10217_7);

wire[31:0] addr_10218_7;

Selector_2 s10218_7(wires_2554_6[2], addr_2554_6, addr_positional[40875:40872], addr_10218_7);

wire[31:0] addr_10219_7;

Selector_2 s10219_7(wires_2554_6[3], addr_2554_6, addr_positional[40879:40876], addr_10219_7);

wire[31:0] addr_10220_7;

Selector_2 s10220_7(wires_2555_6[0], addr_2555_6, addr_positional[40883:40880], addr_10220_7);

wire[31:0] addr_10221_7;

Selector_2 s10221_7(wires_2555_6[1], addr_2555_6, addr_positional[40887:40884], addr_10221_7);

wire[31:0] addr_10222_7;

Selector_2 s10222_7(wires_2555_6[2], addr_2555_6, addr_positional[40891:40888], addr_10222_7);

wire[31:0] addr_10223_7;

Selector_2 s10223_7(wires_2555_6[3], addr_2555_6, addr_positional[40895:40892], addr_10223_7);

wire[31:0] addr_10224_7;

Selector_2 s10224_7(wires_2556_6[0], addr_2556_6, addr_positional[40899:40896], addr_10224_7);

wire[31:0] addr_10225_7;

Selector_2 s10225_7(wires_2556_6[1], addr_2556_6, addr_positional[40903:40900], addr_10225_7);

wire[31:0] addr_10226_7;

Selector_2 s10226_7(wires_2556_6[2], addr_2556_6, addr_positional[40907:40904], addr_10226_7);

wire[31:0] addr_10227_7;

Selector_2 s10227_7(wires_2556_6[3], addr_2556_6, addr_positional[40911:40908], addr_10227_7);

wire[31:0] addr_10228_7;

Selector_2 s10228_7(wires_2557_6[0], addr_2557_6, addr_positional[40915:40912], addr_10228_7);

wire[31:0] addr_10229_7;

Selector_2 s10229_7(wires_2557_6[1], addr_2557_6, addr_positional[40919:40916], addr_10229_7);

wire[31:0] addr_10230_7;

Selector_2 s10230_7(wires_2557_6[2], addr_2557_6, addr_positional[40923:40920], addr_10230_7);

wire[31:0] addr_10231_7;

Selector_2 s10231_7(wires_2557_6[3], addr_2557_6, addr_positional[40927:40924], addr_10231_7);

wire[31:0] addr_10232_7;

Selector_2 s10232_7(wires_2558_6[0], addr_2558_6, addr_positional[40931:40928], addr_10232_7);

wire[31:0] addr_10233_7;

Selector_2 s10233_7(wires_2558_6[1], addr_2558_6, addr_positional[40935:40932], addr_10233_7);

wire[31:0] addr_10234_7;

Selector_2 s10234_7(wires_2558_6[2], addr_2558_6, addr_positional[40939:40936], addr_10234_7);

wire[31:0] addr_10235_7;

Selector_2 s10235_7(wires_2558_6[3], addr_2558_6, addr_positional[40943:40940], addr_10235_7);

wire[31:0] addr_10236_7;

Selector_2 s10236_7(wires_2559_6[0], addr_2559_6, addr_positional[40947:40944], addr_10236_7);

wire[31:0] addr_10237_7;

Selector_2 s10237_7(wires_2559_6[1], addr_2559_6, addr_positional[40951:40948], addr_10237_7);

wire[31:0] addr_10238_7;

Selector_2 s10238_7(wires_2559_6[2], addr_2559_6, addr_positional[40955:40952], addr_10238_7);

wire[31:0] addr_10239_7;

Selector_2 s10239_7(wires_2559_6[3], addr_2559_6, addr_positional[40959:40956], addr_10239_7);

wire[31:0] addr_10240_7;

Selector_2 s10240_7(wires_2560_6[0], addr_2560_6, addr_positional[40963:40960], addr_10240_7);

wire[31:0] addr_10241_7;

Selector_2 s10241_7(wires_2560_6[1], addr_2560_6, addr_positional[40967:40964], addr_10241_7);

wire[31:0] addr_10242_7;

Selector_2 s10242_7(wires_2560_6[2], addr_2560_6, addr_positional[40971:40968], addr_10242_7);

wire[31:0] addr_10243_7;

Selector_2 s10243_7(wires_2560_6[3], addr_2560_6, addr_positional[40975:40972], addr_10243_7);

wire[31:0] addr_10244_7;

Selector_2 s10244_7(wires_2561_6[0], addr_2561_6, addr_positional[40979:40976], addr_10244_7);

wire[31:0] addr_10245_7;

Selector_2 s10245_7(wires_2561_6[1], addr_2561_6, addr_positional[40983:40980], addr_10245_7);

wire[31:0] addr_10246_7;

Selector_2 s10246_7(wires_2561_6[2], addr_2561_6, addr_positional[40987:40984], addr_10246_7);

wire[31:0] addr_10247_7;

Selector_2 s10247_7(wires_2561_6[3], addr_2561_6, addr_positional[40991:40988], addr_10247_7);

wire[31:0] addr_10248_7;

Selector_2 s10248_7(wires_2562_6[0], addr_2562_6, addr_positional[40995:40992], addr_10248_7);

wire[31:0] addr_10249_7;

Selector_2 s10249_7(wires_2562_6[1], addr_2562_6, addr_positional[40999:40996], addr_10249_7);

wire[31:0] addr_10250_7;

Selector_2 s10250_7(wires_2562_6[2], addr_2562_6, addr_positional[41003:41000], addr_10250_7);

wire[31:0] addr_10251_7;

Selector_2 s10251_7(wires_2562_6[3], addr_2562_6, addr_positional[41007:41004], addr_10251_7);

wire[31:0] addr_10252_7;

Selector_2 s10252_7(wires_2563_6[0], addr_2563_6, addr_positional[41011:41008], addr_10252_7);

wire[31:0] addr_10253_7;

Selector_2 s10253_7(wires_2563_6[1], addr_2563_6, addr_positional[41015:41012], addr_10253_7);

wire[31:0] addr_10254_7;

Selector_2 s10254_7(wires_2563_6[2], addr_2563_6, addr_positional[41019:41016], addr_10254_7);

wire[31:0] addr_10255_7;

Selector_2 s10255_7(wires_2563_6[3], addr_2563_6, addr_positional[41023:41020], addr_10255_7);

wire[31:0] addr_10256_7;

Selector_2 s10256_7(wires_2564_6[0], addr_2564_6, addr_positional[41027:41024], addr_10256_7);

wire[31:0] addr_10257_7;

Selector_2 s10257_7(wires_2564_6[1], addr_2564_6, addr_positional[41031:41028], addr_10257_7);

wire[31:0] addr_10258_7;

Selector_2 s10258_7(wires_2564_6[2], addr_2564_6, addr_positional[41035:41032], addr_10258_7);

wire[31:0] addr_10259_7;

Selector_2 s10259_7(wires_2564_6[3], addr_2564_6, addr_positional[41039:41036], addr_10259_7);

wire[31:0] addr_10260_7;

Selector_2 s10260_7(wires_2565_6[0], addr_2565_6, addr_positional[41043:41040], addr_10260_7);

wire[31:0] addr_10261_7;

Selector_2 s10261_7(wires_2565_6[1], addr_2565_6, addr_positional[41047:41044], addr_10261_7);

wire[31:0] addr_10262_7;

Selector_2 s10262_7(wires_2565_6[2], addr_2565_6, addr_positional[41051:41048], addr_10262_7);

wire[31:0] addr_10263_7;

Selector_2 s10263_7(wires_2565_6[3], addr_2565_6, addr_positional[41055:41052], addr_10263_7);

wire[31:0] addr_10264_7;

Selector_2 s10264_7(wires_2566_6[0], addr_2566_6, addr_positional[41059:41056], addr_10264_7);

wire[31:0] addr_10265_7;

Selector_2 s10265_7(wires_2566_6[1], addr_2566_6, addr_positional[41063:41060], addr_10265_7);

wire[31:0] addr_10266_7;

Selector_2 s10266_7(wires_2566_6[2], addr_2566_6, addr_positional[41067:41064], addr_10266_7);

wire[31:0] addr_10267_7;

Selector_2 s10267_7(wires_2566_6[3], addr_2566_6, addr_positional[41071:41068], addr_10267_7);

wire[31:0] addr_10268_7;

Selector_2 s10268_7(wires_2567_6[0], addr_2567_6, addr_positional[41075:41072], addr_10268_7);

wire[31:0] addr_10269_7;

Selector_2 s10269_7(wires_2567_6[1], addr_2567_6, addr_positional[41079:41076], addr_10269_7);

wire[31:0] addr_10270_7;

Selector_2 s10270_7(wires_2567_6[2], addr_2567_6, addr_positional[41083:41080], addr_10270_7);

wire[31:0] addr_10271_7;

Selector_2 s10271_7(wires_2567_6[3], addr_2567_6, addr_positional[41087:41084], addr_10271_7);

wire[31:0] addr_10272_7;

Selector_2 s10272_7(wires_2568_6[0], addr_2568_6, addr_positional[41091:41088], addr_10272_7);

wire[31:0] addr_10273_7;

Selector_2 s10273_7(wires_2568_6[1], addr_2568_6, addr_positional[41095:41092], addr_10273_7);

wire[31:0] addr_10274_7;

Selector_2 s10274_7(wires_2568_6[2], addr_2568_6, addr_positional[41099:41096], addr_10274_7);

wire[31:0] addr_10275_7;

Selector_2 s10275_7(wires_2568_6[3], addr_2568_6, addr_positional[41103:41100], addr_10275_7);

wire[31:0] addr_10276_7;

Selector_2 s10276_7(wires_2569_6[0], addr_2569_6, addr_positional[41107:41104], addr_10276_7);

wire[31:0] addr_10277_7;

Selector_2 s10277_7(wires_2569_6[1], addr_2569_6, addr_positional[41111:41108], addr_10277_7);

wire[31:0] addr_10278_7;

Selector_2 s10278_7(wires_2569_6[2], addr_2569_6, addr_positional[41115:41112], addr_10278_7);

wire[31:0] addr_10279_7;

Selector_2 s10279_7(wires_2569_6[3], addr_2569_6, addr_positional[41119:41116], addr_10279_7);

wire[31:0] addr_10280_7;

Selector_2 s10280_7(wires_2570_6[0], addr_2570_6, addr_positional[41123:41120], addr_10280_7);

wire[31:0] addr_10281_7;

Selector_2 s10281_7(wires_2570_6[1], addr_2570_6, addr_positional[41127:41124], addr_10281_7);

wire[31:0] addr_10282_7;

Selector_2 s10282_7(wires_2570_6[2], addr_2570_6, addr_positional[41131:41128], addr_10282_7);

wire[31:0] addr_10283_7;

Selector_2 s10283_7(wires_2570_6[3], addr_2570_6, addr_positional[41135:41132], addr_10283_7);

wire[31:0] addr_10284_7;

Selector_2 s10284_7(wires_2571_6[0], addr_2571_6, addr_positional[41139:41136], addr_10284_7);

wire[31:0] addr_10285_7;

Selector_2 s10285_7(wires_2571_6[1], addr_2571_6, addr_positional[41143:41140], addr_10285_7);

wire[31:0] addr_10286_7;

Selector_2 s10286_7(wires_2571_6[2], addr_2571_6, addr_positional[41147:41144], addr_10286_7);

wire[31:0] addr_10287_7;

Selector_2 s10287_7(wires_2571_6[3], addr_2571_6, addr_positional[41151:41148], addr_10287_7);

wire[31:0] addr_10288_7;

Selector_2 s10288_7(wires_2572_6[0], addr_2572_6, addr_positional[41155:41152], addr_10288_7);

wire[31:0] addr_10289_7;

Selector_2 s10289_7(wires_2572_6[1], addr_2572_6, addr_positional[41159:41156], addr_10289_7);

wire[31:0] addr_10290_7;

Selector_2 s10290_7(wires_2572_6[2], addr_2572_6, addr_positional[41163:41160], addr_10290_7);

wire[31:0] addr_10291_7;

Selector_2 s10291_7(wires_2572_6[3], addr_2572_6, addr_positional[41167:41164], addr_10291_7);

wire[31:0] addr_10292_7;

Selector_2 s10292_7(wires_2573_6[0], addr_2573_6, addr_positional[41171:41168], addr_10292_7);

wire[31:0] addr_10293_7;

Selector_2 s10293_7(wires_2573_6[1], addr_2573_6, addr_positional[41175:41172], addr_10293_7);

wire[31:0] addr_10294_7;

Selector_2 s10294_7(wires_2573_6[2], addr_2573_6, addr_positional[41179:41176], addr_10294_7);

wire[31:0] addr_10295_7;

Selector_2 s10295_7(wires_2573_6[3], addr_2573_6, addr_positional[41183:41180], addr_10295_7);

wire[31:0] addr_10296_7;

Selector_2 s10296_7(wires_2574_6[0], addr_2574_6, addr_positional[41187:41184], addr_10296_7);

wire[31:0] addr_10297_7;

Selector_2 s10297_7(wires_2574_6[1], addr_2574_6, addr_positional[41191:41188], addr_10297_7);

wire[31:0] addr_10298_7;

Selector_2 s10298_7(wires_2574_6[2], addr_2574_6, addr_positional[41195:41192], addr_10298_7);

wire[31:0] addr_10299_7;

Selector_2 s10299_7(wires_2574_6[3], addr_2574_6, addr_positional[41199:41196], addr_10299_7);

wire[31:0] addr_10300_7;

Selector_2 s10300_7(wires_2575_6[0], addr_2575_6, addr_positional[41203:41200], addr_10300_7);

wire[31:0] addr_10301_7;

Selector_2 s10301_7(wires_2575_6[1], addr_2575_6, addr_positional[41207:41204], addr_10301_7);

wire[31:0] addr_10302_7;

Selector_2 s10302_7(wires_2575_6[2], addr_2575_6, addr_positional[41211:41208], addr_10302_7);

wire[31:0] addr_10303_7;

Selector_2 s10303_7(wires_2575_6[3], addr_2575_6, addr_positional[41215:41212], addr_10303_7);

wire[31:0] addr_10304_7;

Selector_2 s10304_7(wires_2576_6[0], addr_2576_6, addr_positional[41219:41216], addr_10304_7);

wire[31:0] addr_10305_7;

Selector_2 s10305_7(wires_2576_6[1], addr_2576_6, addr_positional[41223:41220], addr_10305_7);

wire[31:0] addr_10306_7;

Selector_2 s10306_7(wires_2576_6[2], addr_2576_6, addr_positional[41227:41224], addr_10306_7);

wire[31:0] addr_10307_7;

Selector_2 s10307_7(wires_2576_6[3], addr_2576_6, addr_positional[41231:41228], addr_10307_7);

wire[31:0] addr_10308_7;

Selector_2 s10308_7(wires_2577_6[0], addr_2577_6, addr_positional[41235:41232], addr_10308_7);

wire[31:0] addr_10309_7;

Selector_2 s10309_7(wires_2577_6[1], addr_2577_6, addr_positional[41239:41236], addr_10309_7);

wire[31:0] addr_10310_7;

Selector_2 s10310_7(wires_2577_6[2], addr_2577_6, addr_positional[41243:41240], addr_10310_7);

wire[31:0] addr_10311_7;

Selector_2 s10311_7(wires_2577_6[3], addr_2577_6, addr_positional[41247:41244], addr_10311_7);

wire[31:0] addr_10312_7;

Selector_2 s10312_7(wires_2578_6[0], addr_2578_6, addr_positional[41251:41248], addr_10312_7);

wire[31:0] addr_10313_7;

Selector_2 s10313_7(wires_2578_6[1], addr_2578_6, addr_positional[41255:41252], addr_10313_7);

wire[31:0] addr_10314_7;

Selector_2 s10314_7(wires_2578_6[2], addr_2578_6, addr_positional[41259:41256], addr_10314_7);

wire[31:0] addr_10315_7;

Selector_2 s10315_7(wires_2578_6[3], addr_2578_6, addr_positional[41263:41260], addr_10315_7);

wire[31:0] addr_10316_7;

Selector_2 s10316_7(wires_2579_6[0], addr_2579_6, addr_positional[41267:41264], addr_10316_7);

wire[31:0] addr_10317_7;

Selector_2 s10317_7(wires_2579_6[1], addr_2579_6, addr_positional[41271:41268], addr_10317_7);

wire[31:0] addr_10318_7;

Selector_2 s10318_7(wires_2579_6[2], addr_2579_6, addr_positional[41275:41272], addr_10318_7);

wire[31:0] addr_10319_7;

Selector_2 s10319_7(wires_2579_6[3], addr_2579_6, addr_positional[41279:41276], addr_10319_7);

wire[31:0] addr_10320_7;

Selector_2 s10320_7(wires_2580_6[0], addr_2580_6, addr_positional[41283:41280], addr_10320_7);

wire[31:0] addr_10321_7;

Selector_2 s10321_7(wires_2580_6[1], addr_2580_6, addr_positional[41287:41284], addr_10321_7);

wire[31:0] addr_10322_7;

Selector_2 s10322_7(wires_2580_6[2], addr_2580_6, addr_positional[41291:41288], addr_10322_7);

wire[31:0] addr_10323_7;

Selector_2 s10323_7(wires_2580_6[3], addr_2580_6, addr_positional[41295:41292], addr_10323_7);

wire[31:0] addr_10324_7;

Selector_2 s10324_7(wires_2581_6[0], addr_2581_6, addr_positional[41299:41296], addr_10324_7);

wire[31:0] addr_10325_7;

Selector_2 s10325_7(wires_2581_6[1], addr_2581_6, addr_positional[41303:41300], addr_10325_7);

wire[31:0] addr_10326_7;

Selector_2 s10326_7(wires_2581_6[2], addr_2581_6, addr_positional[41307:41304], addr_10326_7);

wire[31:0] addr_10327_7;

Selector_2 s10327_7(wires_2581_6[3], addr_2581_6, addr_positional[41311:41308], addr_10327_7);

wire[31:0] addr_10328_7;

Selector_2 s10328_7(wires_2582_6[0], addr_2582_6, addr_positional[41315:41312], addr_10328_7);

wire[31:0] addr_10329_7;

Selector_2 s10329_7(wires_2582_6[1], addr_2582_6, addr_positional[41319:41316], addr_10329_7);

wire[31:0] addr_10330_7;

Selector_2 s10330_7(wires_2582_6[2], addr_2582_6, addr_positional[41323:41320], addr_10330_7);

wire[31:0] addr_10331_7;

Selector_2 s10331_7(wires_2582_6[3], addr_2582_6, addr_positional[41327:41324], addr_10331_7);

wire[31:0] addr_10332_7;

Selector_2 s10332_7(wires_2583_6[0], addr_2583_6, addr_positional[41331:41328], addr_10332_7);

wire[31:0] addr_10333_7;

Selector_2 s10333_7(wires_2583_6[1], addr_2583_6, addr_positional[41335:41332], addr_10333_7);

wire[31:0] addr_10334_7;

Selector_2 s10334_7(wires_2583_6[2], addr_2583_6, addr_positional[41339:41336], addr_10334_7);

wire[31:0] addr_10335_7;

Selector_2 s10335_7(wires_2583_6[3], addr_2583_6, addr_positional[41343:41340], addr_10335_7);

wire[31:0] addr_10336_7;

Selector_2 s10336_7(wires_2584_6[0], addr_2584_6, addr_positional[41347:41344], addr_10336_7);

wire[31:0] addr_10337_7;

Selector_2 s10337_7(wires_2584_6[1], addr_2584_6, addr_positional[41351:41348], addr_10337_7);

wire[31:0] addr_10338_7;

Selector_2 s10338_7(wires_2584_6[2], addr_2584_6, addr_positional[41355:41352], addr_10338_7);

wire[31:0] addr_10339_7;

Selector_2 s10339_7(wires_2584_6[3], addr_2584_6, addr_positional[41359:41356], addr_10339_7);

wire[31:0] addr_10340_7;

Selector_2 s10340_7(wires_2585_6[0], addr_2585_6, addr_positional[41363:41360], addr_10340_7);

wire[31:0] addr_10341_7;

Selector_2 s10341_7(wires_2585_6[1], addr_2585_6, addr_positional[41367:41364], addr_10341_7);

wire[31:0] addr_10342_7;

Selector_2 s10342_7(wires_2585_6[2], addr_2585_6, addr_positional[41371:41368], addr_10342_7);

wire[31:0] addr_10343_7;

Selector_2 s10343_7(wires_2585_6[3], addr_2585_6, addr_positional[41375:41372], addr_10343_7);

wire[31:0] addr_10344_7;

Selector_2 s10344_7(wires_2586_6[0], addr_2586_6, addr_positional[41379:41376], addr_10344_7);

wire[31:0] addr_10345_7;

Selector_2 s10345_7(wires_2586_6[1], addr_2586_6, addr_positional[41383:41380], addr_10345_7);

wire[31:0] addr_10346_7;

Selector_2 s10346_7(wires_2586_6[2], addr_2586_6, addr_positional[41387:41384], addr_10346_7);

wire[31:0] addr_10347_7;

Selector_2 s10347_7(wires_2586_6[3], addr_2586_6, addr_positional[41391:41388], addr_10347_7);

wire[31:0] addr_10348_7;

Selector_2 s10348_7(wires_2587_6[0], addr_2587_6, addr_positional[41395:41392], addr_10348_7);

wire[31:0] addr_10349_7;

Selector_2 s10349_7(wires_2587_6[1], addr_2587_6, addr_positional[41399:41396], addr_10349_7);

wire[31:0] addr_10350_7;

Selector_2 s10350_7(wires_2587_6[2], addr_2587_6, addr_positional[41403:41400], addr_10350_7);

wire[31:0] addr_10351_7;

Selector_2 s10351_7(wires_2587_6[3], addr_2587_6, addr_positional[41407:41404], addr_10351_7);

wire[31:0] addr_10352_7;

Selector_2 s10352_7(wires_2588_6[0], addr_2588_6, addr_positional[41411:41408], addr_10352_7);

wire[31:0] addr_10353_7;

Selector_2 s10353_7(wires_2588_6[1], addr_2588_6, addr_positional[41415:41412], addr_10353_7);

wire[31:0] addr_10354_7;

Selector_2 s10354_7(wires_2588_6[2], addr_2588_6, addr_positional[41419:41416], addr_10354_7);

wire[31:0] addr_10355_7;

Selector_2 s10355_7(wires_2588_6[3], addr_2588_6, addr_positional[41423:41420], addr_10355_7);

wire[31:0] addr_10356_7;

Selector_2 s10356_7(wires_2589_6[0], addr_2589_6, addr_positional[41427:41424], addr_10356_7);

wire[31:0] addr_10357_7;

Selector_2 s10357_7(wires_2589_6[1], addr_2589_6, addr_positional[41431:41428], addr_10357_7);

wire[31:0] addr_10358_7;

Selector_2 s10358_7(wires_2589_6[2], addr_2589_6, addr_positional[41435:41432], addr_10358_7);

wire[31:0] addr_10359_7;

Selector_2 s10359_7(wires_2589_6[3], addr_2589_6, addr_positional[41439:41436], addr_10359_7);

wire[31:0] addr_10360_7;

Selector_2 s10360_7(wires_2590_6[0], addr_2590_6, addr_positional[41443:41440], addr_10360_7);

wire[31:0] addr_10361_7;

Selector_2 s10361_7(wires_2590_6[1], addr_2590_6, addr_positional[41447:41444], addr_10361_7);

wire[31:0] addr_10362_7;

Selector_2 s10362_7(wires_2590_6[2], addr_2590_6, addr_positional[41451:41448], addr_10362_7);

wire[31:0] addr_10363_7;

Selector_2 s10363_7(wires_2590_6[3], addr_2590_6, addr_positional[41455:41452], addr_10363_7);

wire[31:0] addr_10364_7;

Selector_2 s10364_7(wires_2591_6[0], addr_2591_6, addr_positional[41459:41456], addr_10364_7);

wire[31:0] addr_10365_7;

Selector_2 s10365_7(wires_2591_6[1], addr_2591_6, addr_positional[41463:41460], addr_10365_7);

wire[31:0] addr_10366_7;

Selector_2 s10366_7(wires_2591_6[2], addr_2591_6, addr_positional[41467:41464], addr_10366_7);

wire[31:0] addr_10367_7;

Selector_2 s10367_7(wires_2591_6[3], addr_2591_6, addr_positional[41471:41468], addr_10367_7);

wire[31:0] addr_10368_7;

Selector_2 s10368_7(wires_2592_6[0], addr_2592_6, addr_positional[41475:41472], addr_10368_7);

wire[31:0] addr_10369_7;

Selector_2 s10369_7(wires_2592_6[1], addr_2592_6, addr_positional[41479:41476], addr_10369_7);

wire[31:0] addr_10370_7;

Selector_2 s10370_7(wires_2592_6[2], addr_2592_6, addr_positional[41483:41480], addr_10370_7);

wire[31:0] addr_10371_7;

Selector_2 s10371_7(wires_2592_6[3], addr_2592_6, addr_positional[41487:41484], addr_10371_7);

wire[31:0] addr_10372_7;

Selector_2 s10372_7(wires_2593_6[0], addr_2593_6, addr_positional[41491:41488], addr_10372_7);

wire[31:0] addr_10373_7;

Selector_2 s10373_7(wires_2593_6[1], addr_2593_6, addr_positional[41495:41492], addr_10373_7);

wire[31:0] addr_10374_7;

Selector_2 s10374_7(wires_2593_6[2], addr_2593_6, addr_positional[41499:41496], addr_10374_7);

wire[31:0] addr_10375_7;

Selector_2 s10375_7(wires_2593_6[3], addr_2593_6, addr_positional[41503:41500], addr_10375_7);

wire[31:0] addr_10376_7;

Selector_2 s10376_7(wires_2594_6[0], addr_2594_6, addr_positional[41507:41504], addr_10376_7);

wire[31:0] addr_10377_7;

Selector_2 s10377_7(wires_2594_6[1], addr_2594_6, addr_positional[41511:41508], addr_10377_7);

wire[31:0] addr_10378_7;

Selector_2 s10378_7(wires_2594_6[2], addr_2594_6, addr_positional[41515:41512], addr_10378_7);

wire[31:0] addr_10379_7;

Selector_2 s10379_7(wires_2594_6[3], addr_2594_6, addr_positional[41519:41516], addr_10379_7);

wire[31:0] addr_10380_7;

Selector_2 s10380_7(wires_2595_6[0], addr_2595_6, addr_positional[41523:41520], addr_10380_7);

wire[31:0] addr_10381_7;

Selector_2 s10381_7(wires_2595_6[1], addr_2595_6, addr_positional[41527:41524], addr_10381_7);

wire[31:0] addr_10382_7;

Selector_2 s10382_7(wires_2595_6[2], addr_2595_6, addr_positional[41531:41528], addr_10382_7);

wire[31:0] addr_10383_7;

Selector_2 s10383_7(wires_2595_6[3], addr_2595_6, addr_positional[41535:41532], addr_10383_7);

wire[31:0] addr_10384_7;

Selector_2 s10384_7(wires_2596_6[0], addr_2596_6, addr_positional[41539:41536], addr_10384_7);

wire[31:0] addr_10385_7;

Selector_2 s10385_7(wires_2596_6[1], addr_2596_6, addr_positional[41543:41540], addr_10385_7);

wire[31:0] addr_10386_7;

Selector_2 s10386_7(wires_2596_6[2], addr_2596_6, addr_positional[41547:41544], addr_10386_7);

wire[31:0] addr_10387_7;

Selector_2 s10387_7(wires_2596_6[3], addr_2596_6, addr_positional[41551:41548], addr_10387_7);

wire[31:0] addr_10388_7;

Selector_2 s10388_7(wires_2597_6[0], addr_2597_6, addr_positional[41555:41552], addr_10388_7);

wire[31:0] addr_10389_7;

Selector_2 s10389_7(wires_2597_6[1], addr_2597_6, addr_positional[41559:41556], addr_10389_7);

wire[31:0] addr_10390_7;

Selector_2 s10390_7(wires_2597_6[2], addr_2597_6, addr_positional[41563:41560], addr_10390_7);

wire[31:0] addr_10391_7;

Selector_2 s10391_7(wires_2597_6[3], addr_2597_6, addr_positional[41567:41564], addr_10391_7);

wire[31:0] addr_10392_7;

Selector_2 s10392_7(wires_2598_6[0], addr_2598_6, addr_positional[41571:41568], addr_10392_7);

wire[31:0] addr_10393_7;

Selector_2 s10393_7(wires_2598_6[1], addr_2598_6, addr_positional[41575:41572], addr_10393_7);

wire[31:0] addr_10394_7;

Selector_2 s10394_7(wires_2598_6[2], addr_2598_6, addr_positional[41579:41576], addr_10394_7);

wire[31:0] addr_10395_7;

Selector_2 s10395_7(wires_2598_6[3], addr_2598_6, addr_positional[41583:41580], addr_10395_7);

wire[31:0] addr_10396_7;

Selector_2 s10396_7(wires_2599_6[0], addr_2599_6, addr_positional[41587:41584], addr_10396_7);

wire[31:0] addr_10397_7;

Selector_2 s10397_7(wires_2599_6[1], addr_2599_6, addr_positional[41591:41588], addr_10397_7);

wire[31:0] addr_10398_7;

Selector_2 s10398_7(wires_2599_6[2], addr_2599_6, addr_positional[41595:41592], addr_10398_7);

wire[31:0] addr_10399_7;

Selector_2 s10399_7(wires_2599_6[3], addr_2599_6, addr_positional[41599:41596], addr_10399_7);

wire[31:0] addr_10400_7;

Selector_2 s10400_7(wires_2600_6[0], addr_2600_6, addr_positional[41603:41600], addr_10400_7);

wire[31:0] addr_10401_7;

Selector_2 s10401_7(wires_2600_6[1], addr_2600_6, addr_positional[41607:41604], addr_10401_7);

wire[31:0] addr_10402_7;

Selector_2 s10402_7(wires_2600_6[2], addr_2600_6, addr_positional[41611:41608], addr_10402_7);

wire[31:0] addr_10403_7;

Selector_2 s10403_7(wires_2600_6[3], addr_2600_6, addr_positional[41615:41612], addr_10403_7);

wire[31:0] addr_10404_7;

Selector_2 s10404_7(wires_2601_6[0], addr_2601_6, addr_positional[41619:41616], addr_10404_7);

wire[31:0] addr_10405_7;

Selector_2 s10405_7(wires_2601_6[1], addr_2601_6, addr_positional[41623:41620], addr_10405_7);

wire[31:0] addr_10406_7;

Selector_2 s10406_7(wires_2601_6[2], addr_2601_6, addr_positional[41627:41624], addr_10406_7);

wire[31:0] addr_10407_7;

Selector_2 s10407_7(wires_2601_6[3], addr_2601_6, addr_positional[41631:41628], addr_10407_7);

wire[31:0] addr_10408_7;

Selector_2 s10408_7(wires_2602_6[0], addr_2602_6, addr_positional[41635:41632], addr_10408_7);

wire[31:0] addr_10409_7;

Selector_2 s10409_7(wires_2602_6[1], addr_2602_6, addr_positional[41639:41636], addr_10409_7);

wire[31:0] addr_10410_7;

Selector_2 s10410_7(wires_2602_6[2], addr_2602_6, addr_positional[41643:41640], addr_10410_7);

wire[31:0] addr_10411_7;

Selector_2 s10411_7(wires_2602_6[3], addr_2602_6, addr_positional[41647:41644], addr_10411_7);

wire[31:0] addr_10412_7;

Selector_2 s10412_7(wires_2603_6[0], addr_2603_6, addr_positional[41651:41648], addr_10412_7);

wire[31:0] addr_10413_7;

Selector_2 s10413_7(wires_2603_6[1], addr_2603_6, addr_positional[41655:41652], addr_10413_7);

wire[31:0] addr_10414_7;

Selector_2 s10414_7(wires_2603_6[2], addr_2603_6, addr_positional[41659:41656], addr_10414_7);

wire[31:0] addr_10415_7;

Selector_2 s10415_7(wires_2603_6[3], addr_2603_6, addr_positional[41663:41660], addr_10415_7);

wire[31:0] addr_10416_7;

Selector_2 s10416_7(wires_2604_6[0], addr_2604_6, addr_positional[41667:41664], addr_10416_7);

wire[31:0] addr_10417_7;

Selector_2 s10417_7(wires_2604_6[1], addr_2604_6, addr_positional[41671:41668], addr_10417_7);

wire[31:0] addr_10418_7;

Selector_2 s10418_7(wires_2604_6[2], addr_2604_6, addr_positional[41675:41672], addr_10418_7);

wire[31:0] addr_10419_7;

Selector_2 s10419_7(wires_2604_6[3], addr_2604_6, addr_positional[41679:41676], addr_10419_7);

wire[31:0] addr_10420_7;

Selector_2 s10420_7(wires_2605_6[0], addr_2605_6, addr_positional[41683:41680], addr_10420_7);

wire[31:0] addr_10421_7;

Selector_2 s10421_7(wires_2605_6[1], addr_2605_6, addr_positional[41687:41684], addr_10421_7);

wire[31:0] addr_10422_7;

Selector_2 s10422_7(wires_2605_6[2], addr_2605_6, addr_positional[41691:41688], addr_10422_7);

wire[31:0] addr_10423_7;

Selector_2 s10423_7(wires_2605_6[3], addr_2605_6, addr_positional[41695:41692], addr_10423_7);

wire[31:0] addr_10424_7;

Selector_2 s10424_7(wires_2606_6[0], addr_2606_6, addr_positional[41699:41696], addr_10424_7);

wire[31:0] addr_10425_7;

Selector_2 s10425_7(wires_2606_6[1], addr_2606_6, addr_positional[41703:41700], addr_10425_7);

wire[31:0] addr_10426_7;

Selector_2 s10426_7(wires_2606_6[2], addr_2606_6, addr_positional[41707:41704], addr_10426_7);

wire[31:0] addr_10427_7;

Selector_2 s10427_7(wires_2606_6[3], addr_2606_6, addr_positional[41711:41708], addr_10427_7);

wire[31:0] addr_10428_7;

Selector_2 s10428_7(wires_2607_6[0], addr_2607_6, addr_positional[41715:41712], addr_10428_7);

wire[31:0] addr_10429_7;

Selector_2 s10429_7(wires_2607_6[1], addr_2607_6, addr_positional[41719:41716], addr_10429_7);

wire[31:0] addr_10430_7;

Selector_2 s10430_7(wires_2607_6[2], addr_2607_6, addr_positional[41723:41720], addr_10430_7);

wire[31:0] addr_10431_7;

Selector_2 s10431_7(wires_2607_6[3], addr_2607_6, addr_positional[41727:41724], addr_10431_7);

wire[31:0] addr_10432_7;

Selector_2 s10432_7(wires_2608_6[0], addr_2608_6, addr_positional[41731:41728], addr_10432_7);

wire[31:0] addr_10433_7;

Selector_2 s10433_7(wires_2608_6[1], addr_2608_6, addr_positional[41735:41732], addr_10433_7);

wire[31:0] addr_10434_7;

Selector_2 s10434_7(wires_2608_6[2], addr_2608_6, addr_positional[41739:41736], addr_10434_7);

wire[31:0] addr_10435_7;

Selector_2 s10435_7(wires_2608_6[3], addr_2608_6, addr_positional[41743:41740], addr_10435_7);

wire[31:0] addr_10436_7;

Selector_2 s10436_7(wires_2609_6[0], addr_2609_6, addr_positional[41747:41744], addr_10436_7);

wire[31:0] addr_10437_7;

Selector_2 s10437_7(wires_2609_6[1], addr_2609_6, addr_positional[41751:41748], addr_10437_7);

wire[31:0] addr_10438_7;

Selector_2 s10438_7(wires_2609_6[2], addr_2609_6, addr_positional[41755:41752], addr_10438_7);

wire[31:0] addr_10439_7;

Selector_2 s10439_7(wires_2609_6[3], addr_2609_6, addr_positional[41759:41756], addr_10439_7);

wire[31:0] addr_10440_7;

Selector_2 s10440_7(wires_2610_6[0], addr_2610_6, addr_positional[41763:41760], addr_10440_7);

wire[31:0] addr_10441_7;

Selector_2 s10441_7(wires_2610_6[1], addr_2610_6, addr_positional[41767:41764], addr_10441_7);

wire[31:0] addr_10442_7;

Selector_2 s10442_7(wires_2610_6[2], addr_2610_6, addr_positional[41771:41768], addr_10442_7);

wire[31:0] addr_10443_7;

Selector_2 s10443_7(wires_2610_6[3], addr_2610_6, addr_positional[41775:41772], addr_10443_7);

wire[31:0] addr_10444_7;

Selector_2 s10444_7(wires_2611_6[0], addr_2611_6, addr_positional[41779:41776], addr_10444_7);

wire[31:0] addr_10445_7;

Selector_2 s10445_7(wires_2611_6[1], addr_2611_6, addr_positional[41783:41780], addr_10445_7);

wire[31:0] addr_10446_7;

Selector_2 s10446_7(wires_2611_6[2], addr_2611_6, addr_positional[41787:41784], addr_10446_7);

wire[31:0] addr_10447_7;

Selector_2 s10447_7(wires_2611_6[3], addr_2611_6, addr_positional[41791:41788], addr_10447_7);

wire[31:0] addr_10448_7;

Selector_2 s10448_7(wires_2612_6[0], addr_2612_6, addr_positional[41795:41792], addr_10448_7);

wire[31:0] addr_10449_7;

Selector_2 s10449_7(wires_2612_6[1], addr_2612_6, addr_positional[41799:41796], addr_10449_7);

wire[31:0] addr_10450_7;

Selector_2 s10450_7(wires_2612_6[2], addr_2612_6, addr_positional[41803:41800], addr_10450_7);

wire[31:0] addr_10451_7;

Selector_2 s10451_7(wires_2612_6[3], addr_2612_6, addr_positional[41807:41804], addr_10451_7);

wire[31:0] addr_10452_7;

Selector_2 s10452_7(wires_2613_6[0], addr_2613_6, addr_positional[41811:41808], addr_10452_7);

wire[31:0] addr_10453_7;

Selector_2 s10453_7(wires_2613_6[1], addr_2613_6, addr_positional[41815:41812], addr_10453_7);

wire[31:0] addr_10454_7;

Selector_2 s10454_7(wires_2613_6[2], addr_2613_6, addr_positional[41819:41816], addr_10454_7);

wire[31:0] addr_10455_7;

Selector_2 s10455_7(wires_2613_6[3], addr_2613_6, addr_positional[41823:41820], addr_10455_7);

wire[31:0] addr_10456_7;

Selector_2 s10456_7(wires_2614_6[0], addr_2614_6, addr_positional[41827:41824], addr_10456_7);

wire[31:0] addr_10457_7;

Selector_2 s10457_7(wires_2614_6[1], addr_2614_6, addr_positional[41831:41828], addr_10457_7);

wire[31:0] addr_10458_7;

Selector_2 s10458_7(wires_2614_6[2], addr_2614_6, addr_positional[41835:41832], addr_10458_7);

wire[31:0] addr_10459_7;

Selector_2 s10459_7(wires_2614_6[3], addr_2614_6, addr_positional[41839:41836], addr_10459_7);

wire[31:0] addr_10460_7;

Selector_2 s10460_7(wires_2615_6[0], addr_2615_6, addr_positional[41843:41840], addr_10460_7);

wire[31:0] addr_10461_7;

Selector_2 s10461_7(wires_2615_6[1], addr_2615_6, addr_positional[41847:41844], addr_10461_7);

wire[31:0] addr_10462_7;

Selector_2 s10462_7(wires_2615_6[2], addr_2615_6, addr_positional[41851:41848], addr_10462_7);

wire[31:0] addr_10463_7;

Selector_2 s10463_7(wires_2615_6[3], addr_2615_6, addr_positional[41855:41852], addr_10463_7);

wire[31:0] addr_10464_7;

Selector_2 s10464_7(wires_2616_6[0], addr_2616_6, addr_positional[41859:41856], addr_10464_7);

wire[31:0] addr_10465_7;

Selector_2 s10465_7(wires_2616_6[1], addr_2616_6, addr_positional[41863:41860], addr_10465_7);

wire[31:0] addr_10466_7;

Selector_2 s10466_7(wires_2616_6[2], addr_2616_6, addr_positional[41867:41864], addr_10466_7);

wire[31:0] addr_10467_7;

Selector_2 s10467_7(wires_2616_6[3], addr_2616_6, addr_positional[41871:41868], addr_10467_7);

wire[31:0] addr_10468_7;

Selector_2 s10468_7(wires_2617_6[0], addr_2617_6, addr_positional[41875:41872], addr_10468_7);

wire[31:0] addr_10469_7;

Selector_2 s10469_7(wires_2617_6[1], addr_2617_6, addr_positional[41879:41876], addr_10469_7);

wire[31:0] addr_10470_7;

Selector_2 s10470_7(wires_2617_6[2], addr_2617_6, addr_positional[41883:41880], addr_10470_7);

wire[31:0] addr_10471_7;

Selector_2 s10471_7(wires_2617_6[3], addr_2617_6, addr_positional[41887:41884], addr_10471_7);

wire[31:0] addr_10472_7;

Selector_2 s10472_7(wires_2618_6[0], addr_2618_6, addr_positional[41891:41888], addr_10472_7);

wire[31:0] addr_10473_7;

Selector_2 s10473_7(wires_2618_6[1], addr_2618_6, addr_positional[41895:41892], addr_10473_7);

wire[31:0] addr_10474_7;

Selector_2 s10474_7(wires_2618_6[2], addr_2618_6, addr_positional[41899:41896], addr_10474_7);

wire[31:0] addr_10475_7;

Selector_2 s10475_7(wires_2618_6[3], addr_2618_6, addr_positional[41903:41900], addr_10475_7);

wire[31:0] addr_10476_7;

Selector_2 s10476_7(wires_2619_6[0], addr_2619_6, addr_positional[41907:41904], addr_10476_7);

wire[31:0] addr_10477_7;

Selector_2 s10477_7(wires_2619_6[1], addr_2619_6, addr_positional[41911:41908], addr_10477_7);

wire[31:0] addr_10478_7;

Selector_2 s10478_7(wires_2619_6[2], addr_2619_6, addr_positional[41915:41912], addr_10478_7);

wire[31:0] addr_10479_7;

Selector_2 s10479_7(wires_2619_6[3], addr_2619_6, addr_positional[41919:41916], addr_10479_7);

wire[31:0] addr_10480_7;

Selector_2 s10480_7(wires_2620_6[0], addr_2620_6, addr_positional[41923:41920], addr_10480_7);

wire[31:0] addr_10481_7;

Selector_2 s10481_7(wires_2620_6[1], addr_2620_6, addr_positional[41927:41924], addr_10481_7);

wire[31:0] addr_10482_7;

Selector_2 s10482_7(wires_2620_6[2], addr_2620_6, addr_positional[41931:41928], addr_10482_7);

wire[31:0] addr_10483_7;

Selector_2 s10483_7(wires_2620_6[3], addr_2620_6, addr_positional[41935:41932], addr_10483_7);

wire[31:0] addr_10484_7;

Selector_2 s10484_7(wires_2621_6[0], addr_2621_6, addr_positional[41939:41936], addr_10484_7);

wire[31:0] addr_10485_7;

Selector_2 s10485_7(wires_2621_6[1], addr_2621_6, addr_positional[41943:41940], addr_10485_7);

wire[31:0] addr_10486_7;

Selector_2 s10486_7(wires_2621_6[2], addr_2621_6, addr_positional[41947:41944], addr_10486_7);

wire[31:0] addr_10487_7;

Selector_2 s10487_7(wires_2621_6[3], addr_2621_6, addr_positional[41951:41948], addr_10487_7);

wire[31:0] addr_10488_7;

Selector_2 s10488_7(wires_2622_6[0], addr_2622_6, addr_positional[41955:41952], addr_10488_7);

wire[31:0] addr_10489_7;

Selector_2 s10489_7(wires_2622_6[1], addr_2622_6, addr_positional[41959:41956], addr_10489_7);

wire[31:0] addr_10490_7;

Selector_2 s10490_7(wires_2622_6[2], addr_2622_6, addr_positional[41963:41960], addr_10490_7);

wire[31:0] addr_10491_7;

Selector_2 s10491_7(wires_2622_6[3], addr_2622_6, addr_positional[41967:41964], addr_10491_7);

wire[31:0] addr_10492_7;

Selector_2 s10492_7(wires_2623_6[0], addr_2623_6, addr_positional[41971:41968], addr_10492_7);

wire[31:0] addr_10493_7;

Selector_2 s10493_7(wires_2623_6[1], addr_2623_6, addr_positional[41975:41972], addr_10493_7);

wire[31:0] addr_10494_7;

Selector_2 s10494_7(wires_2623_6[2], addr_2623_6, addr_positional[41979:41976], addr_10494_7);

wire[31:0] addr_10495_7;

Selector_2 s10495_7(wires_2623_6[3], addr_2623_6, addr_positional[41983:41980], addr_10495_7);

wire[31:0] addr_10496_7;

Selector_2 s10496_7(wires_2624_6[0], addr_2624_6, addr_positional[41987:41984], addr_10496_7);

wire[31:0] addr_10497_7;

Selector_2 s10497_7(wires_2624_6[1], addr_2624_6, addr_positional[41991:41988], addr_10497_7);

wire[31:0] addr_10498_7;

Selector_2 s10498_7(wires_2624_6[2], addr_2624_6, addr_positional[41995:41992], addr_10498_7);

wire[31:0] addr_10499_7;

Selector_2 s10499_7(wires_2624_6[3], addr_2624_6, addr_positional[41999:41996], addr_10499_7);

wire[31:0] addr_10500_7;

Selector_2 s10500_7(wires_2625_6[0], addr_2625_6, addr_positional[42003:42000], addr_10500_7);

wire[31:0] addr_10501_7;

Selector_2 s10501_7(wires_2625_6[1], addr_2625_6, addr_positional[42007:42004], addr_10501_7);

wire[31:0] addr_10502_7;

Selector_2 s10502_7(wires_2625_6[2], addr_2625_6, addr_positional[42011:42008], addr_10502_7);

wire[31:0] addr_10503_7;

Selector_2 s10503_7(wires_2625_6[3], addr_2625_6, addr_positional[42015:42012], addr_10503_7);

wire[31:0] addr_10504_7;

Selector_2 s10504_7(wires_2626_6[0], addr_2626_6, addr_positional[42019:42016], addr_10504_7);

wire[31:0] addr_10505_7;

Selector_2 s10505_7(wires_2626_6[1], addr_2626_6, addr_positional[42023:42020], addr_10505_7);

wire[31:0] addr_10506_7;

Selector_2 s10506_7(wires_2626_6[2], addr_2626_6, addr_positional[42027:42024], addr_10506_7);

wire[31:0] addr_10507_7;

Selector_2 s10507_7(wires_2626_6[3], addr_2626_6, addr_positional[42031:42028], addr_10507_7);

wire[31:0] addr_10508_7;

Selector_2 s10508_7(wires_2627_6[0], addr_2627_6, addr_positional[42035:42032], addr_10508_7);

wire[31:0] addr_10509_7;

Selector_2 s10509_7(wires_2627_6[1], addr_2627_6, addr_positional[42039:42036], addr_10509_7);

wire[31:0] addr_10510_7;

Selector_2 s10510_7(wires_2627_6[2], addr_2627_6, addr_positional[42043:42040], addr_10510_7);

wire[31:0] addr_10511_7;

Selector_2 s10511_7(wires_2627_6[3], addr_2627_6, addr_positional[42047:42044], addr_10511_7);

wire[31:0] addr_10512_7;

Selector_2 s10512_7(wires_2628_6[0], addr_2628_6, addr_positional[42051:42048], addr_10512_7);

wire[31:0] addr_10513_7;

Selector_2 s10513_7(wires_2628_6[1], addr_2628_6, addr_positional[42055:42052], addr_10513_7);

wire[31:0] addr_10514_7;

Selector_2 s10514_7(wires_2628_6[2], addr_2628_6, addr_positional[42059:42056], addr_10514_7);

wire[31:0] addr_10515_7;

Selector_2 s10515_7(wires_2628_6[3], addr_2628_6, addr_positional[42063:42060], addr_10515_7);

wire[31:0] addr_10516_7;

Selector_2 s10516_7(wires_2629_6[0], addr_2629_6, addr_positional[42067:42064], addr_10516_7);

wire[31:0] addr_10517_7;

Selector_2 s10517_7(wires_2629_6[1], addr_2629_6, addr_positional[42071:42068], addr_10517_7);

wire[31:0] addr_10518_7;

Selector_2 s10518_7(wires_2629_6[2], addr_2629_6, addr_positional[42075:42072], addr_10518_7);

wire[31:0] addr_10519_7;

Selector_2 s10519_7(wires_2629_6[3], addr_2629_6, addr_positional[42079:42076], addr_10519_7);

wire[31:0] addr_10520_7;

Selector_2 s10520_7(wires_2630_6[0], addr_2630_6, addr_positional[42083:42080], addr_10520_7);

wire[31:0] addr_10521_7;

Selector_2 s10521_7(wires_2630_6[1], addr_2630_6, addr_positional[42087:42084], addr_10521_7);

wire[31:0] addr_10522_7;

Selector_2 s10522_7(wires_2630_6[2], addr_2630_6, addr_positional[42091:42088], addr_10522_7);

wire[31:0] addr_10523_7;

Selector_2 s10523_7(wires_2630_6[3], addr_2630_6, addr_positional[42095:42092], addr_10523_7);

wire[31:0] addr_10524_7;

Selector_2 s10524_7(wires_2631_6[0], addr_2631_6, addr_positional[42099:42096], addr_10524_7);

wire[31:0] addr_10525_7;

Selector_2 s10525_7(wires_2631_6[1], addr_2631_6, addr_positional[42103:42100], addr_10525_7);

wire[31:0] addr_10526_7;

Selector_2 s10526_7(wires_2631_6[2], addr_2631_6, addr_positional[42107:42104], addr_10526_7);

wire[31:0] addr_10527_7;

Selector_2 s10527_7(wires_2631_6[3], addr_2631_6, addr_positional[42111:42108], addr_10527_7);

wire[31:0] addr_10528_7;

Selector_2 s10528_7(wires_2632_6[0], addr_2632_6, addr_positional[42115:42112], addr_10528_7);

wire[31:0] addr_10529_7;

Selector_2 s10529_7(wires_2632_6[1], addr_2632_6, addr_positional[42119:42116], addr_10529_7);

wire[31:0] addr_10530_7;

Selector_2 s10530_7(wires_2632_6[2], addr_2632_6, addr_positional[42123:42120], addr_10530_7);

wire[31:0] addr_10531_7;

Selector_2 s10531_7(wires_2632_6[3], addr_2632_6, addr_positional[42127:42124], addr_10531_7);

wire[31:0] addr_10532_7;

Selector_2 s10532_7(wires_2633_6[0], addr_2633_6, addr_positional[42131:42128], addr_10532_7);

wire[31:0] addr_10533_7;

Selector_2 s10533_7(wires_2633_6[1], addr_2633_6, addr_positional[42135:42132], addr_10533_7);

wire[31:0] addr_10534_7;

Selector_2 s10534_7(wires_2633_6[2], addr_2633_6, addr_positional[42139:42136], addr_10534_7);

wire[31:0] addr_10535_7;

Selector_2 s10535_7(wires_2633_6[3], addr_2633_6, addr_positional[42143:42140], addr_10535_7);

wire[31:0] addr_10536_7;

Selector_2 s10536_7(wires_2634_6[0], addr_2634_6, addr_positional[42147:42144], addr_10536_7);

wire[31:0] addr_10537_7;

Selector_2 s10537_7(wires_2634_6[1], addr_2634_6, addr_positional[42151:42148], addr_10537_7);

wire[31:0] addr_10538_7;

Selector_2 s10538_7(wires_2634_6[2], addr_2634_6, addr_positional[42155:42152], addr_10538_7);

wire[31:0] addr_10539_7;

Selector_2 s10539_7(wires_2634_6[3], addr_2634_6, addr_positional[42159:42156], addr_10539_7);

wire[31:0] addr_10540_7;

Selector_2 s10540_7(wires_2635_6[0], addr_2635_6, addr_positional[42163:42160], addr_10540_7);

wire[31:0] addr_10541_7;

Selector_2 s10541_7(wires_2635_6[1], addr_2635_6, addr_positional[42167:42164], addr_10541_7);

wire[31:0] addr_10542_7;

Selector_2 s10542_7(wires_2635_6[2], addr_2635_6, addr_positional[42171:42168], addr_10542_7);

wire[31:0] addr_10543_7;

Selector_2 s10543_7(wires_2635_6[3], addr_2635_6, addr_positional[42175:42172], addr_10543_7);

wire[31:0] addr_10544_7;

Selector_2 s10544_7(wires_2636_6[0], addr_2636_6, addr_positional[42179:42176], addr_10544_7);

wire[31:0] addr_10545_7;

Selector_2 s10545_7(wires_2636_6[1], addr_2636_6, addr_positional[42183:42180], addr_10545_7);

wire[31:0] addr_10546_7;

Selector_2 s10546_7(wires_2636_6[2], addr_2636_6, addr_positional[42187:42184], addr_10546_7);

wire[31:0] addr_10547_7;

Selector_2 s10547_7(wires_2636_6[3], addr_2636_6, addr_positional[42191:42188], addr_10547_7);

wire[31:0] addr_10548_7;

Selector_2 s10548_7(wires_2637_6[0], addr_2637_6, addr_positional[42195:42192], addr_10548_7);

wire[31:0] addr_10549_7;

Selector_2 s10549_7(wires_2637_6[1], addr_2637_6, addr_positional[42199:42196], addr_10549_7);

wire[31:0] addr_10550_7;

Selector_2 s10550_7(wires_2637_6[2], addr_2637_6, addr_positional[42203:42200], addr_10550_7);

wire[31:0] addr_10551_7;

Selector_2 s10551_7(wires_2637_6[3], addr_2637_6, addr_positional[42207:42204], addr_10551_7);

wire[31:0] addr_10552_7;

Selector_2 s10552_7(wires_2638_6[0], addr_2638_6, addr_positional[42211:42208], addr_10552_7);

wire[31:0] addr_10553_7;

Selector_2 s10553_7(wires_2638_6[1], addr_2638_6, addr_positional[42215:42212], addr_10553_7);

wire[31:0] addr_10554_7;

Selector_2 s10554_7(wires_2638_6[2], addr_2638_6, addr_positional[42219:42216], addr_10554_7);

wire[31:0] addr_10555_7;

Selector_2 s10555_7(wires_2638_6[3], addr_2638_6, addr_positional[42223:42220], addr_10555_7);

wire[31:0] addr_10556_7;

Selector_2 s10556_7(wires_2639_6[0], addr_2639_6, addr_positional[42227:42224], addr_10556_7);

wire[31:0] addr_10557_7;

Selector_2 s10557_7(wires_2639_6[1], addr_2639_6, addr_positional[42231:42228], addr_10557_7);

wire[31:0] addr_10558_7;

Selector_2 s10558_7(wires_2639_6[2], addr_2639_6, addr_positional[42235:42232], addr_10558_7);

wire[31:0] addr_10559_7;

Selector_2 s10559_7(wires_2639_6[3], addr_2639_6, addr_positional[42239:42236], addr_10559_7);

wire[31:0] addr_10560_7;

Selector_2 s10560_7(wires_2640_6[0], addr_2640_6, addr_positional[42243:42240], addr_10560_7);

wire[31:0] addr_10561_7;

Selector_2 s10561_7(wires_2640_6[1], addr_2640_6, addr_positional[42247:42244], addr_10561_7);

wire[31:0] addr_10562_7;

Selector_2 s10562_7(wires_2640_6[2], addr_2640_6, addr_positional[42251:42248], addr_10562_7);

wire[31:0] addr_10563_7;

Selector_2 s10563_7(wires_2640_6[3], addr_2640_6, addr_positional[42255:42252], addr_10563_7);

wire[31:0] addr_10564_7;

Selector_2 s10564_7(wires_2641_6[0], addr_2641_6, addr_positional[42259:42256], addr_10564_7);

wire[31:0] addr_10565_7;

Selector_2 s10565_7(wires_2641_6[1], addr_2641_6, addr_positional[42263:42260], addr_10565_7);

wire[31:0] addr_10566_7;

Selector_2 s10566_7(wires_2641_6[2], addr_2641_6, addr_positional[42267:42264], addr_10566_7);

wire[31:0] addr_10567_7;

Selector_2 s10567_7(wires_2641_6[3], addr_2641_6, addr_positional[42271:42268], addr_10567_7);

wire[31:0] addr_10568_7;

Selector_2 s10568_7(wires_2642_6[0], addr_2642_6, addr_positional[42275:42272], addr_10568_7);

wire[31:0] addr_10569_7;

Selector_2 s10569_7(wires_2642_6[1], addr_2642_6, addr_positional[42279:42276], addr_10569_7);

wire[31:0] addr_10570_7;

Selector_2 s10570_7(wires_2642_6[2], addr_2642_6, addr_positional[42283:42280], addr_10570_7);

wire[31:0] addr_10571_7;

Selector_2 s10571_7(wires_2642_6[3], addr_2642_6, addr_positional[42287:42284], addr_10571_7);

wire[31:0] addr_10572_7;

Selector_2 s10572_7(wires_2643_6[0], addr_2643_6, addr_positional[42291:42288], addr_10572_7);

wire[31:0] addr_10573_7;

Selector_2 s10573_7(wires_2643_6[1], addr_2643_6, addr_positional[42295:42292], addr_10573_7);

wire[31:0] addr_10574_7;

Selector_2 s10574_7(wires_2643_6[2], addr_2643_6, addr_positional[42299:42296], addr_10574_7);

wire[31:0] addr_10575_7;

Selector_2 s10575_7(wires_2643_6[3], addr_2643_6, addr_positional[42303:42300], addr_10575_7);

wire[31:0] addr_10576_7;

Selector_2 s10576_7(wires_2644_6[0], addr_2644_6, addr_positional[42307:42304], addr_10576_7);

wire[31:0] addr_10577_7;

Selector_2 s10577_7(wires_2644_6[1], addr_2644_6, addr_positional[42311:42308], addr_10577_7);

wire[31:0] addr_10578_7;

Selector_2 s10578_7(wires_2644_6[2], addr_2644_6, addr_positional[42315:42312], addr_10578_7);

wire[31:0] addr_10579_7;

Selector_2 s10579_7(wires_2644_6[3], addr_2644_6, addr_positional[42319:42316], addr_10579_7);

wire[31:0] addr_10580_7;

Selector_2 s10580_7(wires_2645_6[0], addr_2645_6, addr_positional[42323:42320], addr_10580_7);

wire[31:0] addr_10581_7;

Selector_2 s10581_7(wires_2645_6[1], addr_2645_6, addr_positional[42327:42324], addr_10581_7);

wire[31:0] addr_10582_7;

Selector_2 s10582_7(wires_2645_6[2], addr_2645_6, addr_positional[42331:42328], addr_10582_7);

wire[31:0] addr_10583_7;

Selector_2 s10583_7(wires_2645_6[3], addr_2645_6, addr_positional[42335:42332], addr_10583_7);

wire[31:0] addr_10584_7;

Selector_2 s10584_7(wires_2646_6[0], addr_2646_6, addr_positional[42339:42336], addr_10584_7);

wire[31:0] addr_10585_7;

Selector_2 s10585_7(wires_2646_6[1], addr_2646_6, addr_positional[42343:42340], addr_10585_7);

wire[31:0] addr_10586_7;

Selector_2 s10586_7(wires_2646_6[2], addr_2646_6, addr_positional[42347:42344], addr_10586_7);

wire[31:0] addr_10587_7;

Selector_2 s10587_7(wires_2646_6[3], addr_2646_6, addr_positional[42351:42348], addr_10587_7);

wire[31:0] addr_10588_7;

Selector_2 s10588_7(wires_2647_6[0], addr_2647_6, addr_positional[42355:42352], addr_10588_7);

wire[31:0] addr_10589_7;

Selector_2 s10589_7(wires_2647_6[1], addr_2647_6, addr_positional[42359:42356], addr_10589_7);

wire[31:0] addr_10590_7;

Selector_2 s10590_7(wires_2647_6[2], addr_2647_6, addr_positional[42363:42360], addr_10590_7);

wire[31:0] addr_10591_7;

Selector_2 s10591_7(wires_2647_6[3], addr_2647_6, addr_positional[42367:42364], addr_10591_7);

wire[31:0] addr_10592_7;

Selector_2 s10592_7(wires_2648_6[0], addr_2648_6, addr_positional[42371:42368], addr_10592_7);

wire[31:0] addr_10593_7;

Selector_2 s10593_7(wires_2648_6[1], addr_2648_6, addr_positional[42375:42372], addr_10593_7);

wire[31:0] addr_10594_7;

Selector_2 s10594_7(wires_2648_6[2], addr_2648_6, addr_positional[42379:42376], addr_10594_7);

wire[31:0] addr_10595_7;

Selector_2 s10595_7(wires_2648_6[3], addr_2648_6, addr_positional[42383:42380], addr_10595_7);

wire[31:0] addr_10596_7;

Selector_2 s10596_7(wires_2649_6[0], addr_2649_6, addr_positional[42387:42384], addr_10596_7);

wire[31:0] addr_10597_7;

Selector_2 s10597_7(wires_2649_6[1], addr_2649_6, addr_positional[42391:42388], addr_10597_7);

wire[31:0] addr_10598_7;

Selector_2 s10598_7(wires_2649_6[2], addr_2649_6, addr_positional[42395:42392], addr_10598_7);

wire[31:0] addr_10599_7;

Selector_2 s10599_7(wires_2649_6[3], addr_2649_6, addr_positional[42399:42396], addr_10599_7);

wire[31:0] addr_10600_7;

Selector_2 s10600_7(wires_2650_6[0], addr_2650_6, addr_positional[42403:42400], addr_10600_7);

wire[31:0] addr_10601_7;

Selector_2 s10601_7(wires_2650_6[1], addr_2650_6, addr_positional[42407:42404], addr_10601_7);

wire[31:0] addr_10602_7;

Selector_2 s10602_7(wires_2650_6[2], addr_2650_6, addr_positional[42411:42408], addr_10602_7);

wire[31:0] addr_10603_7;

Selector_2 s10603_7(wires_2650_6[3], addr_2650_6, addr_positional[42415:42412], addr_10603_7);

wire[31:0] addr_10604_7;

Selector_2 s10604_7(wires_2651_6[0], addr_2651_6, addr_positional[42419:42416], addr_10604_7);

wire[31:0] addr_10605_7;

Selector_2 s10605_7(wires_2651_6[1], addr_2651_6, addr_positional[42423:42420], addr_10605_7);

wire[31:0] addr_10606_7;

Selector_2 s10606_7(wires_2651_6[2], addr_2651_6, addr_positional[42427:42424], addr_10606_7);

wire[31:0] addr_10607_7;

Selector_2 s10607_7(wires_2651_6[3], addr_2651_6, addr_positional[42431:42428], addr_10607_7);

wire[31:0] addr_10608_7;

Selector_2 s10608_7(wires_2652_6[0], addr_2652_6, addr_positional[42435:42432], addr_10608_7);

wire[31:0] addr_10609_7;

Selector_2 s10609_7(wires_2652_6[1], addr_2652_6, addr_positional[42439:42436], addr_10609_7);

wire[31:0] addr_10610_7;

Selector_2 s10610_7(wires_2652_6[2], addr_2652_6, addr_positional[42443:42440], addr_10610_7);

wire[31:0] addr_10611_7;

Selector_2 s10611_7(wires_2652_6[3], addr_2652_6, addr_positional[42447:42444], addr_10611_7);

wire[31:0] addr_10612_7;

Selector_2 s10612_7(wires_2653_6[0], addr_2653_6, addr_positional[42451:42448], addr_10612_7);

wire[31:0] addr_10613_7;

Selector_2 s10613_7(wires_2653_6[1], addr_2653_6, addr_positional[42455:42452], addr_10613_7);

wire[31:0] addr_10614_7;

Selector_2 s10614_7(wires_2653_6[2], addr_2653_6, addr_positional[42459:42456], addr_10614_7);

wire[31:0] addr_10615_7;

Selector_2 s10615_7(wires_2653_6[3], addr_2653_6, addr_positional[42463:42460], addr_10615_7);

wire[31:0] addr_10616_7;

Selector_2 s10616_7(wires_2654_6[0], addr_2654_6, addr_positional[42467:42464], addr_10616_7);

wire[31:0] addr_10617_7;

Selector_2 s10617_7(wires_2654_6[1], addr_2654_6, addr_positional[42471:42468], addr_10617_7);

wire[31:0] addr_10618_7;

Selector_2 s10618_7(wires_2654_6[2], addr_2654_6, addr_positional[42475:42472], addr_10618_7);

wire[31:0] addr_10619_7;

Selector_2 s10619_7(wires_2654_6[3], addr_2654_6, addr_positional[42479:42476], addr_10619_7);

wire[31:0] addr_10620_7;

Selector_2 s10620_7(wires_2655_6[0], addr_2655_6, addr_positional[42483:42480], addr_10620_7);

wire[31:0] addr_10621_7;

Selector_2 s10621_7(wires_2655_6[1], addr_2655_6, addr_positional[42487:42484], addr_10621_7);

wire[31:0] addr_10622_7;

Selector_2 s10622_7(wires_2655_6[2], addr_2655_6, addr_positional[42491:42488], addr_10622_7);

wire[31:0] addr_10623_7;

Selector_2 s10623_7(wires_2655_6[3], addr_2655_6, addr_positional[42495:42492], addr_10623_7);

wire[31:0] addr_10624_7;

Selector_2 s10624_7(wires_2656_6[0], addr_2656_6, addr_positional[42499:42496], addr_10624_7);

wire[31:0] addr_10625_7;

Selector_2 s10625_7(wires_2656_6[1], addr_2656_6, addr_positional[42503:42500], addr_10625_7);

wire[31:0] addr_10626_7;

Selector_2 s10626_7(wires_2656_6[2], addr_2656_6, addr_positional[42507:42504], addr_10626_7);

wire[31:0] addr_10627_7;

Selector_2 s10627_7(wires_2656_6[3], addr_2656_6, addr_positional[42511:42508], addr_10627_7);

wire[31:0] addr_10628_7;

Selector_2 s10628_7(wires_2657_6[0], addr_2657_6, addr_positional[42515:42512], addr_10628_7);

wire[31:0] addr_10629_7;

Selector_2 s10629_7(wires_2657_6[1], addr_2657_6, addr_positional[42519:42516], addr_10629_7);

wire[31:0] addr_10630_7;

Selector_2 s10630_7(wires_2657_6[2], addr_2657_6, addr_positional[42523:42520], addr_10630_7);

wire[31:0] addr_10631_7;

Selector_2 s10631_7(wires_2657_6[3], addr_2657_6, addr_positional[42527:42524], addr_10631_7);

wire[31:0] addr_10632_7;

Selector_2 s10632_7(wires_2658_6[0], addr_2658_6, addr_positional[42531:42528], addr_10632_7);

wire[31:0] addr_10633_7;

Selector_2 s10633_7(wires_2658_6[1], addr_2658_6, addr_positional[42535:42532], addr_10633_7);

wire[31:0] addr_10634_7;

Selector_2 s10634_7(wires_2658_6[2], addr_2658_6, addr_positional[42539:42536], addr_10634_7);

wire[31:0] addr_10635_7;

Selector_2 s10635_7(wires_2658_6[3], addr_2658_6, addr_positional[42543:42540], addr_10635_7);

wire[31:0] addr_10636_7;

Selector_2 s10636_7(wires_2659_6[0], addr_2659_6, addr_positional[42547:42544], addr_10636_7);

wire[31:0] addr_10637_7;

Selector_2 s10637_7(wires_2659_6[1], addr_2659_6, addr_positional[42551:42548], addr_10637_7);

wire[31:0] addr_10638_7;

Selector_2 s10638_7(wires_2659_6[2], addr_2659_6, addr_positional[42555:42552], addr_10638_7);

wire[31:0] addr_10639_7;

Selector_2 s10639_7(wires_2659_6[3], addr_2659_6, addr_positional[42559:42556], addr_10639_7);

wire[31:0] addr_10640_7;

Selector_2 s10640_7(wires_2660_6[0], addr_2660_6, addr_positional[42563:42560], addr_10640_7);

wire[31:0] addr_10641_7;

Selector_2 s10641_7(wires_2660_6[1], addr_2660_6, addr_positional[42567:42564], addr_10641_7);

wire[31:0] addr_10642_7;

Selector_2 s10642_7(wires_2660_6[2], addr_2660_6, addr_positional[42571:42568], addr_10642_7);

wire[31:0] addr_10643_7;

Selector_2 s10643_7(wires_2660_6[3], addr_2660_6, addr_positional[42575:42572], addr_10643_7);

wire[31:0] addr_10644_7;

Selector_2 s10644_7(wires_2661_6[0], addr_2661_6, addr_positional[42579:42576], addr_10644_7);

wire[31:0] addr_10645_7;

Selector_2 s10645_7(wires_2661_6[1], addr_2661_6, addr_positional[42583:42580], addr_10645_7);

wire[31:0] addr_10646_7;

Selector_2 s10646_7(wires_2661_6[2], addr_2661_6, addr_positional[42587:42584], addr_10646_7);

wire[31:0] addr_10647_7;

Selector_2 s10647_7(wires_2661_6[3], addr_2661_6, addr_positional[42591:42588], addr_10647_7);

wire[31:0] addr_10648_7;

Selector_2 s10648_7(wires_2662_6[0], addr_2662_6, addr_positional[42595:42592], addr_10648_7);

wire[31:0] addr_10649_7;

Selector_2 s10649_7(wires_2662_6[1], addr_2662_6, addr_positional[42599:42596], addr_10649_7);

wire[31:0] addr_10650_7;

Selector_2 s10650_7(wires_2662_6[2], addr_2662_6, addr_positional[42603:42600], addr_10650_7);

wire[31:0] addr_10651_7;

Selector_2 s10651_7(wires_2662_6[3], addr_2662_6, addr_positional[42607:42604], addr_10651_7);

wire[31:0] addr_10652_7;

Selector_2 s10652_7(wires_2663_6[0], addr_2663_6, addr_positional[42611:42608], addr_10652_7);

wire[31:0] addr_10653_7;

Selector_2 s10653_7(wires_2663_6[1], addr_2663_6, addr_positional[42615:42612], addr_10653_7);

wire[31:0] addr_10654_7;

Selector_2 s10654_7(wires_2663_6[2], addr_2663_6, addr_positional[42619:42616], addr_10654_7);

wire[31:0] addr_10655_7;

Selector_2 s10655_7(wires_2663_6[3], addr_2663_6, addr_positional[42623:42620], addr_10655_7);

wire[31:0] addr_10656_7;

Selector_2 s10656_7(wires_2664_6[0], addr_2664_6, addr_positional[42627:42624], addr_10656_7);

wire[31:0] addr_10657_7;

Selector_2 s10657_7(wires_2664_6[1], addr_2664_6, addr_positional[42631:42628], addr_10657_7);

wire[31:0] addr_10658_7;

Selector_2 s10658_7(wires_2664_6[2], addr_2664_6, addr_positional[42635:42632], addr_10658_7);

wire[31:0] addr_10659_7;

Selector_2 s10659_7(wires_2664_6[3], addr_2664_6, addr_positional[42639:42636], addr_10659_7);

wire[31:0] addr_10660_7;

Selector_2 s10660_7(wires_2665_6[0], addr_2665_6, addr_positional[42643:42640], addr_10660_7);

wire[31:0] addr_10661_7;

Selector_2 s10661_7(wires_2665_6[1], addr_2665_6, addr_positional[42647:42644], addr_10661_7);

wire[31:0] addr_10662_7;

Selector_2 s10662_7(wires_2665_6[2], addr_2665_6, addr_positional[42651:42648], addr_10662_7);

wire[31:0] addr_10663_7;

Selector_2 s10663_7(wires_2665_6[3], addr_2665_6, addr_positional[42655:42652], addr_10663_7);

wire[31:0] addr_10664_7;

Selector_2 s10664_7(wires_2666_6[0], addr_2666_6, addr_positional[42659:42656], addr_10664_7);

wire[31:0] addr_10665_7;

Selector_2 s10665_7(wires_2666_6[1], addr_2666_6, addr_positional[42663:42660], addr_10665_7);

wire[31:0] addr_10666_7;

Selector_2 s10666_7(wires_2666_6[2], addr_2666_6, addr_positional[42667:42664], addr_10666_7);

wire[31:0] addr_10667_7;

Selector_2 s10667_7(wires_2666_6[3], addr_2666_6, addr_positional[42671:42668], addr_10667_7);

wire[31:0] addr_10668_7;

Selector_2 s10668_7(wires_2667_6[0], addr_2667_6, addr_positional[42675:42672], addr_10668_7);

wire[31:0] addr_10669_7;

Selector_2 s10669_7(wires_2667_6[1], addr_2667_6, addr_positional[42679:42676], addr_10669_7);

wire[31:0] addr_10670_7;

Selector_2 s10670_7(wires_2667_6[2], addr_2667_6, addr_positional[42683:42680], addr_10670_7);

wire[31:0] addr_10671_7;

Selector_2 s10671_7(wires_2667_6[3], addr_2667_6, addr_positional[42687:42684], addr_10671_7);

wire[31:0] addr_10672_7;

Selector_2 s10672_7(wires_2668_6[0], addr_2668_6, addr_positional[42691:42688], addr_10672_7);

wire[31:0] addr_10673_7;

Selector_2 s10673_7(wires_2668_6[1], addr_2668_6, addr_positional[42695:42692], addr_10673_7);

wire[31:0] addr_10674_7;

Selector_2 s10674_7(wires_2668_6[2], addr_2668_6, addr_positional[42699:42696], addr_10674_7);

wire[31:0] addr_10675_7;

Selector_2 s10675_7(wires_2668_6[3], addr_2668_6, addr_positional[42703:42700], addr_10675_7);

wire[31:0] addr_10676_7;

Selector_2 s10676_7(wires_2669_6[0], addr_2669_6, addr_positional[42707:42704], addr_10676_7);

wire[31:0] addr_10677_7;

Selector_2 s10677_7(wires_2669_6[1], addr_2669_6, addr_positional[42711:42708], addr_10677_7);

wire[31:0] addr_10678_7;

Selector_2 s10678_7(wires_2669_6[2], addr_2669_6, addr_positional[42715:42712], addr_10678_7);

wire[31:0] addr_10679_7;

Selector_2 s10679_7(wires_2669_6[3], addr_2669_6, addr_positional[42719:42716], addr_10679_7);

wire[31:0] addr_10680_7;

Selector_2 s10680_7(wires_2670_6[0], addr_2670_6, addr_positional[42723:42720], addr_10680_7);

wire[31:0] addr_10681_7;

Selector_2 s10681_7(wires_2670_6[1], addr_2670_6, addr_positional[42727:42724], addr_10681_7);

wire[31:0] addr_10682_7;

Selector_2 s10682_7(wires_2670_6[2], addr_2670_6, addr_positional[42731:42728], addr_10682_7);

wire[31:0] addr_10683_7;

Selector_2 s10683_7(wires_2670_6[3], addr_2670_6, addr_positional[42735:42732], addr_10683_7);

wire[31:0] addr_10684_7;

Selector_2 s10684_7(wires_2671_6[0], addr_2671_6, addr_positional[42739:42736], addr_10684_7);

wire[31:0] addr_10685_7;

Selector_2 s10685_7(wires_2671_6[1], addr_2671_6, addr_positional[42743:42740], addr_10685_7);

wire[31:0] addr_10686_7;

Selector_2 s10686_7(wires_2671_6[2], addr_2671_6, addr_positional[42747:42744], addr_10686_7);

wire[31:0] addr_10687_7;

Selector_2 s10687_7(wires_2671_6[3], addr_2671_6, addr_positional[42751:42748], addr_10687_7);

wire[31:0] addr_10688_7;

Selector_2 s10688_7(wires_2672_6[0], addr_2672_6, addr_positional[42755:42752], addr_10688_7);

wire[31:0] addr_10689_7;

Selector_2 s10689_7(wires_2672_6[1], addr_2672_6, addr_positional[42759:42756], addr_10689_7);

wire[31:0] addr_10690_7;

Selector_2 s10690_7(wires_2672_6[2], addr_2672_6, addr_positional[42763:42760], addr_10690_7);

wire[31:0] addr_10691_7;

Selector_2 s10691_7(wires_2672_6[3], addr_2672_6, addr_positional[42767:42764], addr_10691_7);

wire[31:0] addr_10692_7;

Selector_2 s10692_7(wires_2673_6[0], addr_2673_6, addr_positional[42771:42768], addr_10692_7);

wire[31:0] addr_10693_7;

Selector_2 s10693_7(wires_2673_6[1], addr_2673_6, addr_positional[42775:42772], addr_10693_7);

wire[31:0] addr_10694_7;

Selector_2 s10694_7(wires_2673_6[2], addr_2673_6, addr_positional[42779:42776], addr_10694_7);

wire[31:0] addr_10695_7;

Selector_2 s10695_7(wires_2673_6[3], addr_2673_6, addr_positional[42783:42780], addr_10695_7);

wire[31:0] addr_10696_7;

Selector_2 s10696_7(wires_2674_6[0], addr_2674_6, addr_positional[42787:42784], addr_10696_7);

wire[31:0] addr_10697_7;

Selector_2 s10697_7(wires_2674_6[1], addr_2674_6, addr_positional[42791:42788], addr_10697_7);

wire[31:0] addr_10698_7;

Selector_2 s10698_7(wires_2674_6[2], addr_2674_6, addr_positional[42795:42792], addr_10698_7);

wire[31:0] addr_10699_7;

Selector_2 s10699_7(wires_2674_6[3], addr_2674_6, addr_positional[42799:42796], addr_10699_7);

wire[31:0] addr_10700_7;

Selector_2 s10700_7(wires_2675_6[0], addr_2675_6, addr_positional[42803:42800], addr_10700_7);

wire[31:0] addr_10701_7;

Selector_2 s10701_7(wires_2675_6[1], addr_2675_6, addr_positional[42807:42804], addr_10701_7);

wire[31:0] addr_10702_7;

Selector_2 s10702_7(wires_2675_6[2], addr_2675_6, addr_positional[42811:42808], addr_10702_7);

wire[31:0] addr_10703_7;

Selector_2 s10703_7(wires_2675_6[3], addr_2675_6, addr_positional[42815:42812], addr_10703_7);

wire[31:0] addr_10704_7;

Selector_2 s10704_7(wires_2676_6[0], addr_2676_6, addr_positional[42819:42816], addr_10704_7);

wire[31:0] addr_10705_7;

Selector_2 s10705_7(wires_2676_6[1], addr_2676_6, addr_positional[42823:42820], addr_10705_7);

wire[31:0] addr_10706_7;

Selector_2 s10706_7(wires_2676_6[2], addr_2676_6, addr_positional[42827:42824], addr_10706_7);

wire[31:0] addr_10707_7;

Selector_2 s10707_7(wires_2676_6[3], addr_2676_6, addr_positional[42831:42828], addr_10707_7);

wire[31:0] addr_10708_7;

Selector_2 s10708_7(wires_2677_6[0], addr_2677_6, addr_positional[42835:42832], addr_10708_7);

wire[31:0] addr_10709_7;

Selector_2 s10709_7(wires_2677_6[1], addr_2677_6, addr_positional[42839:42836], addr_10709_7);

wire[31:0] addr_10710_7;

Selector_2 s10710_7(wires_2677_6[2], addr_2677_6, addr_positional[42843:42840], addr_10710_7);

wire[31:0] addr_10711_7;

Selector_2 s10711_7(wires_2677_6[3], addr_2677_6, addr_positional[42847:42844], addr_10711_7);

wire[31:0] addr_10712_7;

Selector_2 s10712_7(wires_2678_6[0], addr_2678_6, addr_positional[42851:42848], addr_10712_7);

wire[31:0] addr_10713_7;

Selector_2 s10713_7(wires_2678_6[1], addr_2678_6, addr_positional[42855:42852], addr_10713_7);

wire[31:0] addr_10714_7;

Selector_2 s10714_7(wires_2678_6[2], addr_2678_6, addr_positional[42859:42856], addr_10714_7);

wire[31:0] addr_10715_7;

Selector_2 s10715_7(wires_2678_6[3], addr_2678_6, addr_positional[42863:42860], addr_10715_7);

wire[31:0] addr_10716_7;

Selector_2 s10716_7(wires_2679_6[0], addr_2679_6, addr_positional[42867:42864], addr_10716_7);

wire[31:0] addr_10717_7;

Selector_2 s10717_7(wires_2679_6[1], addr_2679_6, addr_positional[42871:42868], addr_10717_7);

wire[31:0] addr_10718_7;

Selector_2 s10718_7(wires_2679_6[2], addr_2679_6, addr_positional[42875:42872], addr_10718_7);

wire[31:0] addr_10719_7;

Selector_2 s10719_7(wires_2679_6[3], addr_2679_6, addr_positional[42879:42876], addr_10719_7);

wire[31:0] addr_10720_7;

Selector_2 s10720_7(wires_2680_6[0], addr_2680_6, addr_positional[42883:42880], addr_10720_7);

wire[31:0] addr_10721_7;

Selector_2 s10721_7(wires_2680_6[1], addr_2680_6, addr_positional[42887:42884], addr_10721_7);

wire[31:0] addr_10722_7;

Selector_2 s10722_7(wires_2680_6[2], addr_2680_6, addr_positional[42891:42888], addr_10722_7);

wire[31:0] addr_10723_7;

Selector_2 s10723_7(wires_2680_6[3], addr_2680_6, addr_positional[42895:42892], addr_10723_7);

wire[31:0] addr_10724_7;

Selector_2 s10724_7(wires_2681_6[0], addr_2681_6, addr_positional[42899:42896], addr_10724_7);

wire[31:0] addr_10725_7;

Selector_2 s10725_7(wires_2681_6[1], addr_2681_6, addr_positional[42903:42900], addr_10725_7);

wire[31:0] addr_10726_7;

Selector_2 s10726_7(wires_2681_6[2], addr_2681_6, addr_positional[42907:42904], addr_10726_7);

wire[31:0] addr_10727_7;

Selector_2 s10727_7(wires_2681_6[3], addr_2681_6, addr_positional[42911:42908], addr_10727_7);

wire[31:0] addr_10728_7;

Selector_2 s10728_7(wires_2682_6[0], addr_2682_6, addr_positional[42915:42912], addr_10728_7);

wire[31:0] addr_10729_7;

Selector_2 s10729_7(wires_2682_6[1], addr_2682_6, addr_positional[42919:42916], addr_10729_7);

wire[31:0] addr_10730_7;

Selector_2 s10730_7(wires_2682_6[2], addr_2682_6, addr_positional[42923:42920], addr_10730_7);

wire[31:0] addr_10731_7;

Selector_2 s10731_7(wires_2682_6[3], addr_2682_6, addr_positional[42927:42924], addr_10731_7);

wire[31:0] addr_10732_7;

Selector_2 s10732_7(wires_2683_6[0], addr_2683_6, addr_positional[42931:42928], addr_10732_7);

wire[31:0] addr_10733_7;

Selector_2 s10733_7(wires_2683_6[1], addr_2683_6, addr_positional[42935:42932], addr_10733_7);

wire[31:0] addr_10734_7;

Selector_2 s10734_7(wires_2683_6[2], addr_2683_6, addr_positional[42939:42936], addr_10734_7);

wire[31:0] addr_10735_7;

Selector_2 s10735_7(wires_2683_6[3], addr_2683_6, addr_positional[42943:42940], addr_10735_7);

wire[31:0] addr_10736_7;

Selector_2 s10736_7(wires_2684_6[0], addr_2684_6, addr_positional[42947:42944], addr_10736_7);

wire[31:0] addr_10737_7;

Selector_2 s10737_7(wires_2684_6[1], addr_2684_6, addr_positional[42951:42948], addr_10737_7);

wire[31:0] addr_10738_7;

Selector_2 s10738_7(wires_2684_6[2], addr_2684_6, addr_positional[42955:42952], addr_10738_7);

wire[31:0] addr_10739_7;

Selector_2 s10739_7(wires_2684_6[3], addr_2684_6, addr_positional[42959:42956], addr_10739_7);

wire[31:0] addr_10740_7;

Selector_2 s10740_7(wires_2685_6[0], addr_2685_6, addr_positional[42963:42960], addr_10740_7);

wire[31:0] addr_10741_7;

Selector_2 s10741_7(wires_2685_6[1], addr_2685_6, addr_positional[42967:42964], addr_10741_7);

wire[31:0] addr_10742_7;

Selector_2 s10742_7(wires_2685_6[2], addr_2685_6, addr_positional[42971:42968], addr_10742_7);

wire[31:0] addr_10743_7;

Selector_2 s10743_7(wires_2685_6[3], addr_2685_6, addr_positional[42975:42972], addr_10743_7);

wire[31:0] addr_10744_7;

Selector_2 s10744_7(wires_2686_6[0], addr_2686_6, addr_positional[42979:42976], addr_10744_7);

wire[31:0] addr_10745_7;

Selector_2 s10745_7(wires_2686_6[1], addr_2686_6, addr_positional[42983:42980], addr_10745_7);

wire[31:0] addr_10746_7;

Selector_2 s10746_7(wires_2686_6[2], addr_2686_6, addr_positional[42987:42984], addr_10746_7);

wire[31:0] addr_10747_7;

Selector_2 s10747_7(wires_2686_6[3], addr_2686_6, addr_positional[42991:42988], addr_10747_7);

wire[31:0] addr_10748_7;

Selector_2 s10748_7(wires_2687_6[0], addr_2687_6, addr_positional[42995:42992], addr_10748_7);

wire[31:0] addr_10749_7;

Selector_2 s10749_7(wires_2687_6[1], addr_2687_6, addr_positional[42999:42996], addr_10749_7);

wire[31:0] addr_10750_7;

Selector_2 s10750_7(wires_2687_6[2], addr_2687_6, addr_positional[43003:43000], addr_10750_7);

wire[31:0] addr_10751_7;

Selector_2 s10751_7(wires_2687_6[3], addr_2687_6, addr_positional[43007:43004], addr_10751_7);

wire[31:0] addr_10752_7;

Selector_2 s10752_7(wires_2688_6[0], addr_2688_6, addr_positional[43011:43008], addr_10752_7);

wire[31:0] addr_10753_7;

Selector_2 s10753_7(wires_2688_6[1], addr_2688_6, addr_positional[43015:43012], addr_10753_7);

wire[31:0] addr_10754_7;

Selector_2 s10754_7(wires_2688_6[2], addr_2688_6, addr_positional[43019:43016], addr_10754_7);

wire[31:0] addr_10755_7;

Selector_2 s10755_7(wires_2688_6[3], addr_2688_6, addr_positional[43023:43020], addr_10755_7);

wire[31:0] addr_10756_7;

Selector_2 s10756_7(wires_2689_6[0], addr_2689_6, addr_positional[43027:43024], addr_10756_7);

wire[31:0] addr_10757_7;

Selector_2 s10757_7(wires_2689_6[1], addr_2689_6, addr_positional[43031:43028], addr_10757_7);

wire[31:0] addr_10758_7;

Selector_2 s10758_7(wires_2689_6[2], addr_2689_6, addr_positional[43035:43032], addr_10758_7);

wire[31:0] addr_10759_7;

Selector_2 s10759_7(wires_2689_6[3], addr_2689_6, addr_positional[43039:43036], addr_10759_7);

wire[31:0] addr_10760_7;

Selector_2 s10760_7(wires_2690_6[0], addr_2690_6, addr_positional[43043:43040], addr_10760_7);

wire[31:0] addr_10761_7;

Selector_2 s10761_7(wires_2690_6[1], addr_2690_6, addr_positional[43047:43044], addr_10761_7);

wire[31:0] addr_10762_7;

Selector_2 s10762_7(wires_2690_6[2], addr_2690_6, addr_positional[43051:43048], addr_10762_7);

wire[31:0] addr_10763_7;

Selector_2 s10763_7(wires_2690_6[3], addr_2690_6, addr_positional[43055:43052], addr_10763_7);

wire[31:0] addr_10764_7;

Selector_2 s10764_7(wires_2691_6[0], addr_2691_6, addr_positional[43059:43056], addr_10764_7);

wire[31:0] addr_10765_7;

Selector_2 s10765_7(wires_2691_6[1], addr_2691_6, addr_positional[43063:43060], addr_10765_7);

wire[31:0] addr_10766_7;

Selector_2 s10766_7(wires_2691_6[2], addr_2691_6, addr_positional[43067:43064], addr_10766_7);

wire[31:0] addr_10767_7;

Selector_2 s10767_7(wires_2691_6[3], addr_2691_6, addr_positional[43071:43068], addr_10767_7);

wire[31:0] addr_10768_7;

Selector_2 s10768_7(wires_2692_6[0], addr_2692_6, addr_positional[43075:43072], addr_10768_7);

wire[31:0] addr_10769_7;

Selector_2 s10769_7(wires_2692_6[1], addr_2692_6, addr_positional[43079:43076], addr_10769_7);

wire[31:0] addr_10770_7;

Selector_2 s10770_7(wires_2692_6[2], addr_2692_6, addr_positional[43083:43080], addr_10770_7);

wire[31:0] addr_10771_7;

Selector_2 s10771_7(wires_2692_6[3], addr_2692_6, addr_positional[43087:43084], addr_10771_7);

wire[31:0] addr_10772_7;

Selector_2 s10772_7(wires_2693_6[0], addr_2693_6, addr_positional[43091:43088], addr_10772_7);

wire[31:0] addr_10773_7;

Selector_2 s10773_7(wires_2693_6[1], addr_2693_6, addr_positional[43095:43092], addr_10773_7);

wire[31:0] addr_10774_7;

Selector_2 s10774_7(wires_2693_6[2], addr_2693_6, addr_positional[43099:43096], addr_10774_7);

wire[31:0] addr_10775_7;

Selector_2 s10775_7(wires_2693_6[3], addr_2693_6, addr_positional[43103:43100], addr_10775_7);

wire[31:0] addr_10776_7;

Selector_2 s10776_7(wires_2694_6[0], addr_2694_6, addr_positional[43107:43104], addr_10776_7);

wire[31:0] addr_10777_7;

Selector_2 s10777_7(wires_2694_6[1], addr_2694_6, addr_positional[43111:43108], addr_10777_7);

wire[31:0] addr_10778_7;

Selector_2 s10778_7(wires_2694_6[2], addr_2694_6, addr_positional[43115:43112], addr_10778_7);

wire[31:0] addr_10779_7;

Selector_2 s10779_7(wires_2694_6[3], addr_2694_6, addr_positional[43119:43116], addr_10779_7);

wire[31:0] addr_10780_7;

Selector_2 s10780_7(wires_2695_6[0], addr_2695_6, addr_positional[43123:43120], addr_10780_7);

wire[31:0] addr_10781_7;

Selector_2 s10781_7(wires_2695_6[1], addr_2695_6, addr_positional[43127:43124], addr_10781_7);

wire[31:0] addr_10782_7;

Selector_2 s10782_7(wires_2695_6[2], addr_2695_6, addr_positional[43131:43128], addr_10782_7);

wire[31:0] addr_10783_7;

Selector_2 s10783_7(wires_2695_6[3], addr_2695_6, addr_positional[43135:43132], addr_10783_7);

wire[31:0] addr_10784_7;

Selector_2 s10784_7(wires_2696_6[0], addr_2696_6, addr_positional[43139:43136], addr_10784_7);

wire[31:0] addr_10785_7;

Selector_2 s10785_7(wires_2696_6[1], addr_2696_6, addr_positional[43143:43140], addr_10785_7);

wire[31:0] addr_10786_7;

Selector_2 s10786_7(wires_2696_6[2], addr_2696_6, addr_positional[43147:43144], addr_10786_7);

wire[31:0] addr_10787_7;

Selector_2 s10787_7(wires_2696_6[3], addr_2696_6, addr_positional[43151:43148], addr_10787_7);

wire[31:0] addr_10788_7;

Selector_2 s10788_7(wires_2697_6[0], addr_2697_6, addr_positional[43155:43152], addr_10788_7);

wire[31:0] addr_10789_7;

Selector_2 s10789_7(wires_2697_6[1], addr_2697_6, addr_positional[43159:43156], addr_10789_7);

wire[31:0] addr_10790_7;

Selector_2 s10790_7(wires_2697_6[2], addr_2697_6, addr_positional[43163:43160], addr_10790_7);

wire[31:0] addr_10791_7;

Selector_2 s10791_7(wires_2697_6[3], addr_2697_6, addr_positional[43167:43164], addr_10791_7);

wire[31:0] addr_10792_7;

Selector_2 s10792_7(wires_2698_6[0], addr_2698_6, addr_positional[43171:43168], addr_10792_7);

wire[31:0] addr_10793_7;

Selector_2 s10793_7(wires_2698_6[1], addr_2698_6, addr_positional[43175:43172], addr_10793_7);

wire[31:0] addr_10794_7;

Selector_2 s10794_7(wires_2698_6[2], addr_2698_6, addr_positional[43179:43176], addr_10794_7);

wire[31:0] addr_10795_7;

Selector_2 s10795_7(wires_2698_6[3], addr_2698_6, addr_positional[43183:43180], addr_10795_7);

wire[31:0] addr_10796_7;

Selector_2 s10796_7(wires_2699_6[0], addr_2699_6, addr_positional[43187:43184], addr_10796_7);

wire[31:0] addr_10797_7;

Selector_2 s10797_7(wires_2699_6[1], addr_2699_6, addr_positional[43191:43188], addr_10797_7);

wire[31:0] addr_10798_7;

Selector_2 s10798_7(wires_2699_6[2], addr_2699_6, addr_positional[43195:43192], addr_10798_7);

wire[31:0] addr_10799_7;

Selector_2 s10799_7(wires_2699_6[3], addr_2699_6, addr_positional[43199:43196], addr_10799_7);

wire[31:0] addr_10800_7;

Selector_2 s10800_7(wires_2700_6[0], addr_2700_6, addr_positional[43203:43200], addr_10800_7);

wire[31:0] addr_10801_7;

Selector_2 s10801_7(wires_2700_6[1], addr_2700_6, addr_positional[43207:43204], addr_10801_7);

wire[31:0] addr_10802_7;

Selector_2 s10802_7(wires_2700_6[2], addr_2700_6, addr_positional[43211:43208], addr_10802_7);

wire[31:0] addr_10803_7;

Selector_2 s10803_7(wires_2700_6[3], addr_2700_6, addr_positional[43215:43212], addr_10803_7);

wire[31:0] addr_10804_7;

Selector_2 s10804_7(wires_2701_6[0], addr_2701_6, addr_positional[43219:43216], addr_10804_7);

wire[31:0] addr_10805_7;

Selector_2 s10805_7(wires_2701_6[1], addr_2701_6, addr_positional[43223:43220], addr_10805_7);

wire[31:0] addr_10806_7;

Selector_2 s10806_7(wires_2701_6[2], addr_2701_6, addr_positional[43227:43224], addr_10806_7);

wire[31:0] addr_10807_7;

Selector_2 s10807_7(wires_2701_6[3], addr_2701_6, addr_positional[43231:43228], addr_10807_7);

wire[31:0] addr_10808_7;

Selector_2 s10808_7(wires_2702_6[0], addr_2702_6, addr_positional[43235:43232], addr_10808_7);

wire[31:0] addr_10809_7;

Selector_2 s10809_7(wires_2702_6[1], addr_2702_6, addr_positional[43239:43236], addr_10809_7);

wire[31:0] addr_10810_7;

Selector_2 s10810_7(wires_2702_6[2], addr_2702_6, addr_positional[43243:43240], addr_10810_7);

wire[31:0] addr_10811_7;

Selector_2 s10811_7(wires_2702_6[3], addr_2702_6, addr_positional[43247:43244], addr_10811_7);

wire[31:0] addr_10812_7;

Selector_2 s10812_7(wires_2703_6[0], addr_2703_6, addr_positional[43251:43248], addr_10812_7);

wire[31:0] addr_10813_7;

Selector_2 s10813_7(wires_2703_6[1], addr_2703_6, addr_positional[43255:43252], addr_10813_7);

wire[31:0] addr_10814_7;

Selector_2 s10814_7(wires_2703_6[2], addr_2703_6, addr_positional[43259:43256], addr_10814_7);

wire[31:0] addr_10815_7;

Selector_2 s10815_7(wires_2703_6[3], addr_2703_6, addr_positional[43263:43260], addr_10815_7);

wire[31:0] addr_10816_7;

Selector_2 s10816_7(wires_2704_6[0], addr_2704_6, addr_positional[43267:43264], addr_10816_7);

wire[31:0] addr_10817_7;

Selector_2 s10817_7(wires_2704_6[1], addr_2704_6, addr_positional[43271:43268], addr_10817_7);

wire[31:0] addr_10818_7;

Selector_2 s10818_7(wires_2704_6[2], addr_2704_6, addr_positional[43275:43272], addr_10818_7);

wire[31:0] addr_10819_7;

Selector_2 s10819_7(wires_2704_6[3], addr_2704_6, addr_positional[43279:43276], addr_10819_7);

wire[31:0] addr_10820_7;

Selector_2 s10820_7(wires_2705_6[0], addr_2705_6, addr_positional[43283:43280], addr_10820_7);

wire[31:0] addr_10821_7;

Selector_2 s10821_7(wires_2705_6[1], addr_2705_6, addr_positional[43287:43284], addr_10821_7);

wire[31:0] addr_10822_7;

Selector_2 s10822_7(wires_2705_6[2], addr_2705_6, addr_positional[43291:43288], addr_10822_7);

wire[31:0] addr_10823_7;

Selector_2 s10823_7(wires_2705_6[3], addr_2705_6, addr_positional[43295:43292], addr_10823_7);

wire[31:0] addr_10824_7;

Selector_2 s10824_7(wires_2706_6[0], addr_2706_6, addr_positional[43299:43296], addr_10824_7);

wire[31:0] addr_10825_7;

Selector_2 s10825_7(wires_2706_6[1], addr_2706_6, addr_positional[43303:43300], addr_10825_7);

wire[31:0] addr_10826_7;

Selector_2 s10826_7(wires_2706_6[2], addr_2706_6, addr_positional[43307:43304], addr_10826_7);

wire[31:0] addr_10827_7;

Selector_2 s10827_7(wires_2706_6[3], addr_2706_6, addr_positional[43311:43308], addr_10827_7);

wire[31:0] addr_10828_7;

Selector_2 s10828_7(wires_2707_6[0], addr_2707_6, addr_positional[43315:43312], addr_10828_7);

wire[31:0] addr_10829_7;

Selector_2 s10829_7(wires_2707_6[1], addr_2707_6, addr_positional[43319:43316], addr_10829_7);

wire[31:0] addr_10830_7;

Selector_2 s10830_7(wires_2707_6[2], addr_2707_6, addr_positional[43323:43320], addr_10830_7);

wire[31:0] addr_10831_7;

Selector_2 s10831_7(wires_2707_6[3], addr_2707_6, addr_positional[43327:43324], addr_10831_7);

wire[31:0] addr_10832_7;

Selector_2 s10832_7(wires_2708_6[0], addr_2708_6, addr_positional[43331:43328], addr_10832_7);

wire[31:0] addr_10833_7;

Selector_2 s10833_7(wires_2708_6[1], addr_2708_6, addr_positional[43335:43332], addr_10833_7);

wire[31:0] addr_10834_7;

Selector_2 s10834_7(wires_2708_6[2], addr_2708_6, addr_positional[43339:43336], addr_10834_7);

wire[31:0] addr_10835_7;

Selector_2 s10835_7(wires_2708_6[3], addr_2708_6, addr_positional[43343:43340], addr_10835_7);

wire[31:0] addr_10836_7;

Selector_2 s10836_7(wires_2709_6[0], addr_2709_6, addr_positional[43347:43344], addr_10836_7);

wire[31:0] addr_10837_7;

Selector_2 s10837_7(wires_2709_6[1], addr_2709_6, addr_positional[43351:43348], addr_10837_7);

wire[31:0] addr_10838_7;

Selector_2 s10838_7(wires_2709_6[2], addr_2709_6, addr_positional[43355:43352], addr_10838_7);

wire[31:0] addr_10839_7;

Selector_2 s10839_7(wires_2709_6[3], addr_2709_6, addr_positional[43359:43356], addr_10839_7);

wire[31:0] addr_10840_7;

Selector_2 s10840_7(wires_2710_6[0], addr_2710_6, addr_positional[43363:43360], addr_10840_7);

wire[31:0] addr_10841_7;

Selector_2 s10841_7(wires_2710_6[1], addr_2710_6, addr_positional[43367:43364], addr_10841_7);

wire[31:0] addr_10842_7;

Selector_2 s10842_7(wires_2710_6[2], addr_2710_6, addr_positional[43371:43368], addr_10842_7);

wire[31:0] addr_10843_7;

Selector_2 s10843_7(wires_2710_6[3], addr_2710_6, addr_positional[43375:43372], addr_10843_7);

wire[31:0] addr_10844_7;

Selector_2 s10844_7(wires_2711_6[0], addr_2711_6, addr_positional[43379:43376], addr_10844_7);

wire[31:0] addr_10845_7;

Selector_2 s10845_7(wires_2711_6[1], addr_2711_6, addr_positional[43383:43380], addr_10845_7);

wire[31:0] addr_10846_7;

Selector_2 s10846_7(wires_2711_6[2], addr_2711_6, addr_positional[43387:43384], addr_10846_7);

wire[31:0] addr_10847_7;

Selector_2 s10847_7(wires_2711_6[3], addr_2711_6, addr_positional[43391:43388], addr_10847_7);

wire[31:0] addr_10848_7;

Selector_2 s10848_7(wires_2712_6[0], addr_2712_6, addr_positional[43395:43392], addr_10848_7);

wire[31:0] addr_10849_7;

Selector_2 s10849_7(wires_2712_6[1], addr_2712_6, addr_positional[43399:43396], addr_10849_7);

wire[31:0] addr_10850_7;

Selector_2 s10850_7(wires_2712_6[2], addr_2712_6, addr_positional[43403:43400], addr_10850_7);

wire[31:0] addr_10851_7;

Selector_2 s10851_7(wires_2712_6[3], addr_2712_6, addr_positional[43407:43404], addr_10851_7);

wire[31:0] addr_10852_7;

Selector_2 s10852_7(wires_2713_6[0], addr_2713_6, addr_positional[43411:43408], addr_10852_7);

wire[31:0] addr_10853_7;

Selector_2 s10853_7(wires_2713_6[1], addr_2713_6, addr_positional[43415:43412], addr_10853_7);

wire[31:0] addr_10854_7;

Selector_2 s10854_7(wires_2713_6[2], addr_2713_6, addr_positional[43419:43416], addr_10854_7);

wire[31:0] addr_10855_7;

Selector_2 s10855_7(wires_2713_6[3], addr_2713_6, addr_positional[43423:43420], addr_10855_7);

wire[31:0] addr_10856_7;

Selector_2 s10856_7(wires_2714_6[0], addr_2714_6, addr_positional[43427:43424], addr_10856_7);

wire[31:0] addr_10857_7;

Selector_2 s10857_7(wires_2714_6[1], addr_2714_6, addr_positional[43431:43428], addr_10857_7);

wire[31:0] addr_10858_7;

Selector_2 s10858_7(wires_2714_6[2], addr_2714_6, addr_positional[43435:43432], addr_10858_7);

wire[31:0] addr_10859_7;

Selector_2 s10859_7(wires_2714_6[3], addr_2714_6, addr_positional[43439:43436], addr_10859_7);

wire[31:0] addr_10860_7;

Selector_2 s10860_7(wires_2715_6[0], addr_2715_6, addr_positional[43443:43440], addr_10860_7);

wire[31:0] addr_10861_7;

Selector_2 s10861_7(wires_2715_6[1], addr_2715_6, addr_positional[43447:43444], addr_10861_7);

wire[31:0] addr_10862_7;

Selector_2 s10862_7(wires_2715_6[2], addr_2715_6, addr_positional[43451:43448], addr_10862_7);

wire[31:0] addr_10863_7;

Selector_2 s10863_7(wires_2715_6[3], addr_2715_6, addr_positional[43455:43452], addr_10863_7);

wire[31:0] addr_10864_7;

Selector_2 s10864_7(wires_2716_6[0], addr_2716_6, addr_positional[43459:43456], addr_10864_7);

wire[31:0] addr_10865_7;

Selector_2 s10865_7(wires_2716_6[1], addr_2716_6, addr_positional[43463:43460], addr_10865_7);

wire[31:0] addr_10866_7;

Selector_2 s10866_7(wires_2716_6[2], addr_2716_6, addr_positional[43467:43464], addr_10866_7);

wire[31:0] addr_10867_7;

Selector_2 s10867_7(wires_2716_6[3], addr_2716_6, addr_positional[43471:43468], addr_10867_7);

wire[31:0] addr_10868_7;

Selector_2 s10868_7(wires_2717_6[0], addr_2717_6, addr_positional[43475:43472], addr_10868_7);

wire[31:0] addr_10869_7;

Selector_2 s10869_7(wires_2717_6[1], addr_2717_6, addr_positional[43479:43476], addr_10869_7);

wire[31:0] addr_10870_7;

Selector_2 s10870_7(wires_2717_6[2], addr_2717_6, addr_positional[43483:43480], addr_10870_7);

wire[31:0] addr_10871_7;

Selector_2 s10871_7(wires_2717_6[3], addr_2717_6, addr_positional[43487:43484], addr_10871_7);

wire[31:0] addr_10872_7;

Selector_2 s10872_7(wires_2718_6[0], addr_2718_6, addr_positional[43491:43488], addr_10872_7);

wire[31:0] addr_10873_7;

Selector_2 s10873_7(wires_2718_6[1], addr_2718_6, addr_positional[43495:43492], addr_10873_7);

wire[31:0] addr_10874_7;

Selector_2 s10874_7(wires_2718_6[2], addr_2718_6, addr_positional[43499:43496], addr_10874_7);

wire[31:0] addr_10875_7;

Selector_2 s10875_7(wires_2718_6[3], addr_2718_6, addr_positional[43503:43500], addr_10875_7);

wire[31:0] addr_10876_7;

Selector_2 s10876_7(wires_2719_6[0], addr_2719_6, addr_positional[43507:43504], addr_10876_7);

wire[31:0] addr_10877_7;

Selector_2 s10877_7(wires_2719_6[1], addr_2719_6, addr_positional[43511:43508], addr_10877_7);

wire[31:0] addr_10878_7;

Selector_2 s10878_7(wires_2719_6[2], addr_2719_6, addr_positional[43515:43512], addr_10878_7);

wire[31:0] addr_10879_7;

Selector_2 s10879_7(wires_2719_6[3], addr_2719_6, addr_positional[43519:43516], addr_10879_7);

wire[31:0] addr_10880_7;

Selector_2 s10880_7(wires_2720_6[0], addr_2720_6, addr_positional[43523:43520], addr_10880_7);

wire[31:0] addr_10881_7;

Selector_2 s10881_7(wires_2720_6[1], addr_2720_6, addr_positional[43527:43524], addr_10881_7);

wire[31:0] addr_10882_7;

Selector_2 s10882_7(wires_2720_6[2], addr_2720_6, addr_positional[43531:43528], addr_10882_7);

wire[31:0] addr_10883_7;

Selector_2 s10883_7(wires_2720_6[3], addr_2720_6, addr_positional[43535:43532], addr_10883_7);

wire[31:0] addr_10884_7;

Selector_2 s10884_7(wires_2721_6[0], addr_2721_6, addr_positional[43539:43536], addr_10884_7);

wire[31:0] addr_10885_7;

Selector_2 s10885_7(wires_2721_6[1], addr_2721_6, addr_positional[43543:43540], addr_10885_7);

wire[31:0] addr_10886_7;

Selector_2 s10886_7(wires_2721_6[2], addr_2721_6, addr_positional[43547:43544], addr_10886_7);

wire[31:0] addr_10887_7;

Selector_2 s10887_7(wires_2721_6[3], addr_2721_6, addr_positional[43551:43548], addr_10887_7);

wire[31:0] addr_10888_7;

Selector_2 s10888_7(wires_2722_6[0], addr_2722_6, addr_positional[43555:43552], addr_10888_7);

wire[31:0] addr_10889_7;

Selector_2 s10889_7(wires_2722_6[1], addr_2722_6, addr_positional[43559:43556], addr_10889_7);

wire[31:0] addr_10890_7;

Selector_2 s10890_7(wires_2722_6[2], addr_2722_6, addr_positional[43563:43560], addr_10890_7);

wire[31:0] addr_10891_7;

Selector_2 s10891_7(wires_2722_6[3], addr_2722_6, addr_positional[43567:43564], addr_10891_7);

wire[31:0] addr_10892_7;

Selector_2 s10892_7(wires_2723_6[0], addr_2723_6, addr_positional[43571:43568], addr_10892_7);

wire[31:0] addr_10893_7;

Selector_2 s10893_7(wires_2723_6[1], addr_2723_6, addr_positional[43575:43572], addr_10893_7);

wire[31:0] addr_10894_7;

Selector_2 s10894_7(wires_2723_6[2], addr_2723_6, addr_positional[43579:43576], addr_10894_7);

wire[31:0] addr_10895_7;

Selector_2 s10895_7(wires_2723_6[3], addr_2723_6, addr_positional[43583:43580], addr_10895_7);

wire[31:0] addr_10896_7;

Selector_2 s10896_7(wires_2724_6[0], addr_2724_6, addr_positional[43587:43584], addr_10896_7);

wire[31:0] addr_10897_7;

Selector_2 s10897_7(wires_2724_6[1], addr_2724_6, addr_positional[43591:43588], addr_10897_7);

wire[31:0] addr_10898_7;

Selector_2 s10898_7(wires_2724_6[2], addr_2724_6, addr_positional[43595:43592], addr_10898_7);

wire[31:0] addr_10899_7;

Selector_2 s10899_7(wires_2724_6[3], addr_2724_6, addr_positional[43599:43596], addr_10899_7);

wire[31:0] addr_10900_7;

Selector_2 s10900_7(wires_2725_6[0], addr_2725_6, addr_positional[43603:43600], addr_10900_7);

wire[31:0] addr_10901_7;

Selector_2 s10901_7(wires_2725_6[1], addr_2725_6, addr_positional[43607:43604], addr_10901_7);

wire[31:0] addr_10902_7;

Selector_2 s10902_7(wires_2725_6[2], addr_2725_6, addr_positional[43611:43608], addr_10902_7);

wire[31:0] addr_10903_7;

Selector_2 s10903_7(wires_2725_6[3], addr_2725_6, addr_positional[43615:43612], addr_10903_7);

wire[31:0] addr_10904_7;

Selector_2 s10904_7(wires_2726_6[0], addr_2726_6, addr_positional[43619:43616], addr_10904_7);

wire[31:0] addr_10905_7;

Selector_2 s10905_7(wires_2726_6[1], addr_2726_6, addr_positional[43623:43620], addr_10905_7);

wire[31:0] addr_10906_7;

Selector_2 s10906_7(wires_2726_6[2], addr_2726_6, addr_positional[43627:43624], addr_10906_7);

wire[31:0] addr_10907_7;

Selector_2 s10907_7(wires_2726_6[3], addr_2726_6, addr_positional[43631:43628], addr_10907_7);

wire[31:0] addr_10908_7;

Selector_2 s10908_7(wires_2727_6[0], addr_2727_6, addr_positional[43635:43632], addr_10908_7);

wire[31:0] addr_10909_7;

Selector_2 s10909_7(wires_2727_6[1], addr_2727_6, addr_positional[43639:43636], addr_10909_7);

wire[31:0] addr_10910_7;

Selector_2 s10910_7(wires_2727_6[2], addr_2727_6, addr_positional[43643:43640], addr_10910_7);

wire[31:0] addr_10911_7;

Selector_2 s10911_7(wires_2727_6[3], addr_2727_6, addr_positional[43647:43644], addr_10911_7);

wire[31:0] addr_10912_7;

Selector_2 s10912_7(wires_2728_6[0], addr_2728_6, addr_positional[43651:43648], addr_10912_7);

wire[31:0] addr_10913_7;

Selector_2 s10913_7(wires_2728_6[1], addr_2728_6, addr_positional[43655:43652], addr_10913_7);

wire[31:0] addr_10914_7;

Selector_2 s10914_7(wires_2728_6[2], addr_2728_6, addr_positional[43659:43656], addr_10914_7);

wire[31:0] addr_10915_7;

Selector_2 s10915_7(wires_2728_6[3], addr_2728_6, addr_positional[43663:43660], addr_10915_7);

wire[31:0] addr_10916_7;

Selector_2 s10916_7(wires_2729_6[0], addr_2729_6, addr_positional[43667:43664], addr_10916_7);

wire[31:0] addr_10917_7;

Selector_2 s10917_7(wires_2729_6[1], addr_2729_6, addr_positional[43671:43668], addr_10917_7);

wire[31:0] addr_10918_7;

Selector_2 s10918_7(wires_2729_6[2], addr_2729_6, addr_positional[43675:43672], addr_10918_7);

wire[31:0] addr_10919_7;

Selector_2 s10919_7(wires_2729_6[3], addr_2729_6, addr_positional[43679:43676], addr_10919_7);

wire[31:0] addr_10920_7;

Selector_2 s10920_7(wires_2730_6[0], addr_2730_6, addr_positional[43683:43680], addr_10920_7);

wire[31:0] addr_10921_7;

Selector_2 s10921_7(wires_2730_6[1], addr_2730_6, addr_positional[43687:43684], addr_10921_7);

wire[31:0] addr_10922_7;

Selector_2 s10922_7(wires_2730_6[2], addr_2730_6, addr_positional[43691:43688], addr_10922_7);

wire[31:0] addr_10923_7;

Selector_2 s10923_7(wires_2730_6[3], addr_2730_6, addr_positional[43695:43692], addr_10923_7);

wire[31:0] addr_10924_7;

Selector_2 s10924_7(wires_2731_6[0], addr_2731_6, addr_positional[43699:43696], addr_10924_7);

wire[31:0] addr_10925_7;

Selector_2 s10925_7(wires_2731_6[1], addr_2731_6, addr_positional[43703:43700], addr_10925_7);

wire[31:0] addr_10926_7;

Selector_2 s10926_7(wires_2731_6[2], addr_2731_6, addr_positional[43707:43704], addr_10926_7);

wire[31:0] addr_10927_7;

Selector_2 s10927_7(wires_2731_6[3], addr_2731_6, addr_positional[43711:43708], addr_10927_7);

wire[31:0] addr_10928_7;

Selector_2 s10928_7(wires_2732_6[0], addr_2732_6, addr_positional[43715:43712], addr_10928_7);

wire[31:0] addr_10929_7;

Selector_2 s10929_7(wires_2732_6[1], addr_2732_6, addr_positional[43719:43716], addr_10929_7);

wire[31:0] addr_10930_7;

Selector_2 s10930_7(wires_2732_6[2], addr_2732_6, addr_positional[43723:43720], addr_10930_7);

wire[31:0] addr_10931_7;

Selector_2 s10931_7(wires_2732_6[3], addr_2732_6, addr_positional[43727:43724], addr_10931_7);

wire[31:0] addr_10932_7;

Selector_2 s10932_7(wires_2733_6[0], addr_2733_6, addr_positional[43731:43728], addr_10932_7);

wire[31:0] addr_10933_7;

Selector_2 s10933_7(wires_2733_6[1], addr_2733_6, addr_positional[43735:43732], addr_10933_7);

wire[31:0] addr_10934_7;

Selector_2 s10934_7(wires_2733_6[2], addr_2733_6, addr_positional[43739:43736], addr_10934_7);

wire[31:0] addr_10935_7;

Selector_2 s10935_7(wires_2733_6[3], addr_2733_6, addr_positional[43743:43740], addr_10935_7);

wire[31:0] addr_10936_7;

Selector_2 s10936_7(wires_2734_6[0], addr_2734_6, addr_positional[43747:43744], addr_10936_7);

wire[31:0] addr_10937_7;

Selector_2 s10937_7(wires_2734_6[1], addr_2734_6, addr_positional[43751:43748], addr_10937_7);

wire[31:0] addr_10938_7;

Selector_2 s10938_7(wires_2734_6[2], addr_2734_6, addr_positional[43755:43752], addr_10938_7);

wire[31:0] addr_10939_7;

Selector_2 s10939_7(wires_2734_6[3], addr_2734_6, addr_positional[43759:43756], addr_10939_7);

wire[31:0] addr_10940_7;

Selector_2 s10940_7(wires_2735_6[0], addr_2735_6, addr_positional[43763:43760], addr_10940_7);

wire[31:0] addr_10941_7;

Selector_2 s10941_7(wires_2735_6[1], addr_2735_6, addr_positional[43767:43764], addr_10941_7);

wire[31:0] addr_10942_7;

Selector_2 s10942_7(wires_2735_6[2], addr_2735_6, addr_positional[43771:43768], addr_10942_7);

wire[31:0] addr_10943_7;

Selector_2 s10943_7(wires_2735_6[3], addr_2735_6, addr_positional[43775:43772], addr_10943_7);

wire[31:0] addr_10944_7;

Selector_2 s10944_7(wires_2736_6[0], addr_2736_6, addr_positional[43779:43776], addr_10944_7);

wire[31:0] addr_10945_7;

Selector_2 s10945_7(wires_2736_6[1], addr_2736_6, addr_positional[43783:43780], addr_10945_7);

wire[31:0] addr_10946_7;

Selector_2 s10946_7(wires_2736_6[2], addr_2736_6, addr_positional[43787:43784], addr_10946_7);

wire[31:0] addr_10947_7;

Selector_2 s10947_7(wires_2736_6[3], addr_2736_6, addr_positional[43791:43788], addr_10947_7);

wire[31:0] addr_10948_7;

Selector_2 s10948_7(wires_2737_6[0], addr_2737_6, addr_positional[43795:43792], addr_10948_7);

wire[31:0] addr_10949_7;

Selector_2 s10949_7(wires_2737_6[1], addr_2737_6, addr_positional[43799:43796], addr_10949_7);

wire[31:0] addr_10950_7;

Selector_2 s10950_7(wires_2737_6[2], addr_2737_6, addr_positional[43803:43800], addr_10950_7);

wire[31:0] addr_10951_7;

Selector_2 s10951_7(wires_2737_6[3], addr_2737_6, addr_positional[43807:43804], addr_10951_7);

wire[31:0] addr_10952_7;

Selector_2 s10952_7(wires_2738_6[0], addr_2738_6, addr_positional[43811:43808], addr_10952_7);

wire[31:0] addr_10953_7;

Selector_2 s10953_7(wires_2738_6[1], addr_2738_6, addr_positional[43815:43812], addr_10953_7);

wire[31:0] addr_10954_7;

Selector_2 s10954_7(wires_2738_6[2], addr_2738_6, addr_positional[43819:43816], addr_10954_7);

wire[31:0] addr_10955_7;

Selector_2 s10955_7(wires_2738_6[3], addr_2738_6, addr_positional[43823:43820], addr_10955_7);

wire[31:0] addr_10956_7;

Selector_2 s10956_7(wires_2739_6[0], addr_2739_6, addr_positional[43827:43824], addr_10956_7);

wire[31:0] addr_10957_7;

Selector_2 s10957_7(wires_2739_6[1], addr_2739_6, addr_positional[43831:43828], addr_10957_7);

wire[31:0] addr_10958_7;

Selector_2 s10958_7(wires_2739_6[2], addr_2739_6, addr_positional[43835:43832], addr_10958_7);

wire[31:0] addr_10959_7;

Selector_2 s10959_7(wires_2739_6[3], addr_2739_6, addr_positional[43839:43836], addr_10959_7);

wire[31:0] addr_10960_7;

Selector_2 s10960_7(wires_2740_6[0], addr_2740_6, addr_positional[43843:43840], addr_10960_7);

wire[31:0] addr_10961_7;

Selector_2 s10961_7(wires_2740_6[1], addr_2740_6, addr_positional[43847:43844], addr_10961_7);

wire[31:0] addr_10962_7;

Selector_2 s10962_7(wires_2740_6[2], addr_2740_6, addr_positional[43851:43848], addr_10962_7);

wire[31:0] addr_10963_7;

Selector_2 s10963_7(wires_2740_6[3], addr_2740_6, addr_positional[43855:43852], addr_10963_7);

wire[31:0] addr_10964_7;

Selector_2 s10964_7(wires_2741_6[0], addr_2741_6, addr_positional[43859:43856], addr_10964_7);

wire[31:0] addr_10965_7;

Selector_2 s10965_7(wires_2741_6[1], addr_2741_6, addr_positional[43863:43860], addr_10965_7);

wire[31:0] addr_10966_7;

Selector_2 s10966_7(wires_2741_6[2], addr_2741_6, addr_positional[43867:43864], addr_10966_7);

wire[31:0] addr_10967_7;

Selector_2 s10967_7(wires_2741_6[3], addr_2741_6, addr_positional[43871:43868], addr_10967_7);

wire[31:0] addr_10968_7;

Selector_2 s10968_7(wires_2742_6[0], addr_2742_6, addr_positional[43875:43872], addr_10968_7);

wire[31:0] addr_10969_7;

Selector_2 s10969_7(wires_2742_6[1], addr_2742_6, addr_positional[43879:43876], addr_10969_7);

wire[31:0] addr_10970_7;

Selector_2 s10970_7(wires_2742_6[2], addr_2742_6, addr_positional[43883:43880], addr_10970_7);

wire[31:0] addr_10971_7;

Selector_2 s10971_7(wires_2742_6[3], addr_2742_6, addr_positional[43887:43884], addr_10971_7);

wire[31:0] addr_10972_7;

Selector_2 s10972_7(wires_2743_6[0], addr_2743_6, addr_positional[43891:43888], addr_10972_7);

wire[31:0] addr_10973_7;

Selector_2 s10973_7(wires_2743_6[1], addr_2743_6, addr_positional[43895:43892], addr_10973_7);

wire[31:0] addr_10974_7;

Selector_2 s10974_7(wires_2743_6[2], addr_2743_6, addr_positional[43899:43896], addr_10974_7);

wire[31:0] addr_10975_7;

Selector_2 s10975_7(wires_2743_6[3], addr_2743_6, addr_positional[43903:43900], addr_10975_7);

wire[31:0] addr_10976_7;

Selector_2 s10976_7(wires_2744_6[0], addr_2744_6, addr_positional[43907:43904], addr_10976_7);

wire[31:0] addr_10977_7;

Selector_2 s10977_7(wires_2744_6[1], addr_2744_6, addr_positional[43911:43908], addr_10977_7);

wire[31:0] addr_10978_7;

Selector_2 s10978_7(wires_2744_6[2], addr_2744_6, addr_positional[43915:43912], addr_10978_7);

wire[31:0] addr_10979_7;

Selector_2 s10979_7(wires_2744_6[3], addr_2744_6, addr_positional[43919:43916], addr_10979_7);

wire[31:0] addr_10980_7;

Selector_2 s10980_7(wires_2745_6[0], addr_2745_6, addr_positional[43923:43920], addr_10980_7);

wire[31:0] addr_10981_7;

Selector_2 s10981_7(wires_2745_6[1], addr_2745_6, addr_positional[43927:43924], addr_10981_7);

wire[31:0] addr_10982_7;

Selector_2 s10982_7(wires_2745_6[2], addr_2745_6, addr_positional[43931:43928], addr_10982_7);

wire[31:0] addr_10983_7;

Selector_2 s10983_7(wires_2745_6[3], addr_2745_6, addr_positional[43935:43932], addr_10983_7);

wire[31:0] addr_10984_7;

Selector_2 s10984_7(wires_2746_6[0], addr_2746_6, addr_positional[43939:43936], addr_10984_7);

wire[31:0] addr_10985_7;

Selector_2 s10985_7(wires_2746_6[1], addr_2746_6, addr_positional[43943:43940], addr_10985_7);

wire[31:0] addr_10986_7;

Selector_2 s10986_7(wires_2746_6[2], addr_2746_6, addr_positional[43947:43944], addr_10986_7);

wire[31:0] addr_10987_7;

Selector_2 s10987_7(wires_2746_6[3], addr_2746_6, addr_positional[43951:43948], addr_10987_7);

wire[31:0] addr_10988_7;

Selector_2 s10988_7(wires_2747_6[0], addr_2747_6, addr_positional[43955:43952], addr_10988_7);

wire[31:0] addr_10989_7;

Selector_2 s10989_7(wires_2747_6[1], addr_2747_6, addr_positional[43959:43956], addr_10989_7);

wire[31:0] addr_10990_7;

Selector_2 s10990_7(wires_2747_6[2], addr_2747_6, addr_positional[43963:43960], addr_10990_7);

wire[31:0] addr_10991_7;

Selector_2 s10991_7(wires_2747_6[3], addr_2747_6, addr_positional[43967:43964], addr_10991_7);

wire[31:0] addr_10992_7;

Selector_2 s10992_7(wires_2748_6[0], addr_2748_6, addr_positional[43971:43968], addr_10992_7);

wire[31:0] addr_10993_7;

Selector_2 s10993_7(wires_2748_6[1], addr_2748_6, addr_positional[43975:43972], addr_10993_7);

wire[31:0] addr_10994_7;

Selector_2 s10994_7(wires_2748_6[2], addr_2748_6, addr_positional[43979:43976], addr_10994_7);

wire[31:0] addr_10995_7;

Selector_2 s10995_7(wires_2748_6[3], addr_2748_6, addr_positional[43983:43980], addr_10995_7);

wire[31:0] addr_10996_7;

Selector_2 s10996_7(wires_2749_6[0], addr_2749_6, addr_positional[43987:43984], addr_10996_7);

wire[31:0] addr_10997_7;

Selector_2 s10997_7(wires_2749_6[1], addr_2749_6, addr_positional[43991:43988], addr_10997_7);

wire[31:0] addr_10998_7;

Selector_2 s10998_7(wires_2749_6[2], addr_2749_6, addr_positional[43995:43992], addr_10998_7);

wire[31:0] addr_10999_7;

Selector_2 s10999_7(wires_2749_6[3], addr_2749_6, addr_positional[43999:43996], addr_10999_7);

wire[31:0] addr_11000_7;

Selector_2 s11000_7(wires_2750_6[0], addr_2750_6, addr_positional[44003:44000], addr_11000_7);

wire[31:0] addr_11001_7;

Selector_2 s11001_7(wires_2750_6[1], addr_2750_6, addr_positional[44007:44004], addr_11001_7);

wire[31:0] addr_11002_7;

Selector_2 s11002_7(wires_2750_6[2], addr_2750_6, addr_positional[44011:44008], addr_11002_7);

wire[31:0] addr_11003_7;

Selector_2 s11003_7(wires_2750_6[3], addr_2750_6, addr_positional[44015:44012], addr_11003_7);

wire[31:0] addr_11004_7;

Selector_2 s11004_7(wires_2751_6[0], addr_2751_6, addr_positional[44019:44016], addr_11004_7);

wire[31:0] addr_11005_7;

Selector_2 s11005_7(wires_2751_6[1], addr_2751_6, addr_positional[44023:44020], addr_11005_7);

wire[31:0] addr_11006_7;

Selector_2 s11006_7(wires_2751_6[2], addr_2751_6, addr_positional[44027:44024], addr_11006_7);

wire[31:0] addr_11007_7;

Selector_2 s11007_7(wires_2751_6[3], addr_2751_6, addr_positional[44031:44028], addr_11007_7);

wire[31:0] addr_11008_7;

Selector_2 s11008_7(wires_2752_6[0], addr_2752_6, addr_positional[44035:44032], addr_11008_7);

wire[31:0] addr_11009_7;

Selector_2 s11009_7(wires_2752_6[1], addr_2752_6, addr_positional[44039:44036], addr_11009_7);

wire[31:0] addr_11010_7;

Selector_2 s11010_7(wires_2752_6[2], addr_2752_6, addr_positional[44043:44040], addr_11010_7);

wire[31:0] addr_11011_7;

Selector_2 s11011_7(wires_2752_6[3], addr_2752_6, addr_positional[44047:44044], addr_11011_7);

wire[31:0] addr_11012_7;

Selector_2 s11012_7(wires_2753_6[0], addr_2753_6, addr_positional[44051:44048], addr_11012_7);

wire[31:0] addr_11013_7;

Selector_2 s11013_7(wires_2753_6[1], addr_2753_6, addr_positional[44055:44052], addr_11013_7);

wire[31:0] addr_11014_7;

Selector_2 s11014_7(wires_2753_6[2], addr_2753_6, addr_positional[44059:44056], addr_11014_7);

wire[31:0] addr_11015_7;

Selector_2 s11015_7(wires_2753_6[3], addr_2753_6, addr_positional[44063:44060], addr_11015_7);

wire[31:0] addr_11016_7;

Selector_2 s11016_7(wires_2754_6[0], addr_2754_6, addr_positional[44067:44064], addr_11016_7);

wire[31:0] addr_11017_7;

Selector_2 s11017_7(wires_2754_6[1], addr_2754_6, addr_positional[44071:44068], addr_11017_7);

wire[31:0] addr_11018_7;

Selector_2 s11018_7(wires_2754_6[2], addr_2754_6, addr_positional[44075:44072], addr_11018_7);

wire[31:0] addr_11019_7;

Selector_2 s11019_7(wires_2754_6[3], addr_2754_6, addr_positional[44079:44076], addr_11019_7);

wire[31:0] addr_11020_7;

Selector_2 s11020_7(wires_2755_6[0], addr_2755_6, addr_positional[44083:44080], addr_11020_7);

wire[31:0] addr_11021_7;

Selector_2 s11021_7(wires_2755_6[1], addr_2755_6, addr_positional[44087:44084], addr_11021_7);

wire[31:0] addr_11022_7;

Selector_2 s11022_7(wires_2755_6[2], addr_2755_6, addr_positional[44091:44088], addr_11022_7);

wire[31:0] addr_11023_7;

Selector_2 s11023_7(wires_2755_6[3], addr_2755_6, addr_positional[44095:44092], addr_11023_7);

wire[31:0] addr_11024_7;

Selector_2 s11024_7(wires_2756_6[0], addr_2756_6, addr_positional[44099:44096], addr_11024_7);

wire[31:0] addr_11025_7;

Selector_2 s11025_7(wires_2756_6[1], addr_2756_6, addr_positional[44103:44100], addr_11025_7);

wire[31:0] addr_11026_7;

Selector_2 s11026_7(wires_2756_6[2], addr_2756_6, addr_positional[44107:44104], addr_11026_7);

wire[31:0] addr_11027_7;

Selector_2 s11027_7(wires_2756_6[3], addr_2756_6, addr_positional[44111:44108], addr_11027_7);

wire[31:0] addr_11028_7;

Selector_2 s11028_7(wires_2757_6[0], addr_2757_6, addr_positional[44115:44112], addr_11028_7);

wire[31:0] addr_11029_7;

Selector_2 s11029_7(wires_2757_6[1], addr_2757_6, addr_positional[44119:44116], addr_11029_7);

wire[31:0] addr_11030_7;

Selector_2 s11030_7(wires_2757_6[2], addr_2757_6, addr_positional[44123:44120], addr_11030_7);

wire[31:0] addr_11031_7;

Selector_2 s11031_7(wires_2757_6[3], addr_2757_6, addr_positional[44127:44124], addr_11031_7);

wire[31:0] addr_11032_7;

Selector_2 s11032_7(wires_2758_6[0], addr_2758_6, addr_positional[44131:44128], addr_11032_7);

wire[31:0] addr_11033_7;

Selector_2 s11033_7(wires_2758_6[1], addr_2758_6, addr_positional[44135:44132], addr_11033_7);

wire[31:0] addr_11034_7;

Selector_2 s11034_7(wires_2758_6[2], addr_2758_6, addr_positional[44139:44136], addr_11034_7);

wire[31:0] addr_11035_7;

Selector_2 s11035_7(wires_2758_6[3], addr_2758_6, addr_positional[44143:44140], addr_11035_7);

wire[31:0] addr_11036_7;

Selector_2 s11036_7(wires_2759_6[0], addr_2759_6, addr_positional[44147:44144], addr_11036_7);

wire[31:0] addr_11037_7;

Selector_2 s11037_7(wires_2759_6[1], addr_2759_6, addr_positional[44151:44148], addr_11037_7);

wire[31:0] addr_11038_7;

Selector_2 s11038_7(wires_2759_6[2], addr_2759_6, addr_positional[44155:44152], addr_11038_7);

wire[31:0] addr_11039_7;

Selector_2 s11039_7(wires_2759_6[3], addr_2759_6, addr_positional[44159:44156], addr_11039_7);

wire[31:0] addr_11040_7;

Selector_2 s11040_7(wires_2760_6[0], addr_2760_6, addr_positional[44163:44160], addr_11040_7);

wire[31:0] addr_11041_7;

Selector_2 s11041_7(wires_2760_6[1], addr_2760_6, addr_positional[44167:44164], addr_11041_7);

wire[31:0] addr_11042_7;

Selector_2 s11042_7(wires_2760_6[2], addr_2760_6, addr_positional[44171:44168], addr_11042_7);

wire[31:0] addr_11043_7;

Selector_2 s11043_7(wires_2760_6[3], addr_2760_6, addr_positional[44175:44172], addr_11043_7);

wire[31:0] addr_11044_7;

Selector_2 s11044_7(wires_2761_6[0], addr_2761_6, addr_positional[44179:44176], addr_11044_7);

wire[31:0] addr_11045_7;

Selector_2 s11045_7(wires_2761_6[1], addr_2761_6, addr_positional[44183:44180], addr_11045_7);

wire[31:0] addr_11046_7;

Selector_2 s11046_7(wires_2761_6[2], addr_2761_6, addr_positional[44187:44184], addr_11046_7);

wire[31:0] addr_11047_7;

Selector_2 s11047_7(wires_2761_6[3], addr_2761_6, addr_positional[44191:44188], addr_11047_7);

wire[31:0] addr_11048_7;

Selector_2 s11048_7(wires_2762_6[0], addr_2762_6, addr_positional[44195:44192], addr_11048_7);

wire[31:0] addr_11049_7;

Selector_2 s11049_7(wires_2762_6[1], addr_2762_6, addr_positional[44199:44196], addr_11049_7);

wire[31:0] addr_11050_7;

Selector_2 s11050_7(wires_2762_6[2], addr_2762_6, addr_positional[44203:44200], addr_11050_7);

wire[31:0] addr_11051_7;

Selector_2 s11051_7(wires_2762_6[3], addr_2762_6, addr_positional[44207:44204], addr_11051_7);

wire[31:0] addr_11052_7;

Selector_2 s11052_7(wires_2763_6[0], addr_2763_6, addr_positional[44211:44208], addr_11052_7);

wire[31:0] addr_11053_7;

Selector_2 s11053_7(wires_2763_6[1], addr_2763_6, addr_positional[44215:44212], addr_11053_7);

wire[31:0] addr_11054_7;

Selector_2 s11054_7(wires_2763_6[2], addr_2763_6, addr_positional[44219:44216], addr_11054_7);

wire[31:0] addr_11055_7;

Selector_2 s11055_7(wires_2763_6[3], addr_2763_6, addr_positional[44223:44220], addr_11055_7);

wire[31:0] addr_11056_7;

Selector_2 s11056_7(wires_2764_6[0], addr_2764_6, addr_positional[44227:44224], addr_11056_7);

wire[31:0] addr_11057_7;

Selector_2 s11057_7(wires_2764_6[1], addr_2764_6, addr_positional[44231:44228], addr_11057_7);

wire[31:0] addr_11058_7;

Selector_2 s11058_7(wires_2764_6[2], addr_2764_6, addr_positional[44235:44232], addr_11058_7);

wire[31:0] addr_11059_7;

Selector_2 s11059_7(wires_2764_6[3], addr_2764_6, addr_positional[44239:44236], addr_11059_7);

wire[31:0] addr_11060_7;

Selector_2 s11060_7(wires_2765_6[0], addr_2765_6, addr_positional[44243:44240], addr_11060_7);

wire[31:0] addr_11061_7;

Selector_2 s11061_7(wires_2765_6[1], addr_2765_6, addr_positional[44247:44244], addr_11061_7);

wire[31:0] addr_11062_7;

Selector_2 s11062_7(wires_2765_6[2], addr_2765_6, addr_positional[44251:44248], addr_11062_7);

wire[31:0] addr_11063_7;

Selector_2 s11063_7(wires_2765_6[3], addr_2765_6, addr_positional[44255:44252], addr_11063_7);

wire[31:0] addr_11064_7;

Selector_2 s11064_7(wires_2766_6[0], addr_2766_6, addr_positional[44259:44256], addr_11064_7);

wire[31:0] addr_11065_7;

Selector_2 s11065_7(wires_2766_6[1], addr_2766_6, addr_positional[44263:44260], addr_11065_7);

wire[31:0] addr_11066_7;

Selector_2 s11066_7(wires_2766_6[2], addr_2766_6, addr_positional[44267:44264], addr_11066_7);

wire[31:0] addr_11067_7;

Selector_2 s11067_7(wires_2766_6[3], addr_2766_6, addr_positional[44271:44268], addr_11067_7);

wire[31:0] addr_11068_7;

Selector_2 s11068_7(wires_2767_6[0], addr_2767_6, addr_positional[44275:44272], addr_11068_7);

wire[31:0] addr_11069_7;

Selector_2 s11069_7(wires_2767_6[1], addr_2767_6, addr_positional[44279:44276], addr_11069_7);

wire[31:0] addr_11070_7;

Selector_2 s11070_7(wires_2767_6[2], addr_2767_6, addr_positional[44283:44280], addr_11070_7);

wire[31:0] addr_11071_7;

Selector_2 s11071_7(wires_2767_6[3], addr_2767_6, addr_positional[44287:44284], addr_11071_7);

wire[31:0] addr_11072_7;

Selector_2 s11072_7(wires_2768_6[0], addr_2768_6, addr_positional[44291:44288], addr_11072_7);

wire[31:0] addr_11073_7;

Selector_2 s11073_7(wires_2768_6[1], addr_2768_6, addr_positional[44295:44292], addr_11073_7);

wire[31:0] addr_11074_7;

Selector_2 s11074_7(wires_2768_6[2], addr_2768_6, addr_positional[44299:44296], addr_11074_7);

wire[31:0] addr_11075_7;

Selector_2 s11075_7(wires_2768_6[3], addr_2768_6, addr_positional[44303:44300], addr_11075_7);

wire[31:0] addr_11076_7;

Selector_2 s11076_7(wires_2769_6[0], addr_2769_6, addr_positional[44307:44304], addr_11076_7);

wire[31:0] addr_11077_7;

Selector_2 s11077_7(wires_2769_6[1], addr_2769_6, addr_positional[44311:44308], addr_11077_7);

wire[31:0] addr_11078_7;

Selector_2 s11078_7(wires_2769_6[2], addr_2769_6, addr_positional[44315:44312], addr_11078_7);

wire[31:0] addr_11079_7;

Selector_2 s11079_7(wires_2769_6[3], addr_2769_6, addr_positional[44319:44316], addr_11079_7);

wire[31:0] addr_11080_7;

Selector_2 s11080_7(wires_2770_6[0], addr_2770_6, addr_positional[44323:44320], addr_11080_7);

wire[31:0] addr_11081_7;

Selector_2 s11081_7(wires_2770_6[1], addr_2770_6, addr_positional[44327:44324], addr_11081_7);

wire[31:0] addr_11082_7;

Selector_2 s11082_7(wires_2770_6[2], addr_2770_6, addr_positional[44331:44328], addr_11082_7);

wire[31:0] addr_11083_7;

Selector_2 s11083_7(wires_2770_6[3], addr_2770_6, addr_positional[44335:44332], addr_11083_7);

wire[31:0] addr_11084_7;

Selector_2 s11084_7(wires_2771_6[0], addr_2771_6, addr_positional[44339:44336], addr_11084_7);

wire[31:0] addr_11085_7;

Selector_2 s11085_7(wires_2771_6[1], addr_2771_6, addr_positional[44343:44340], addr_11085_7);

wire[31:0] addr_11086_7;

Selector_2 s11086_7(wires_2771_6[2], addr_2771_6, addr_positional[44347:44344], addr_11086_7);

wire[31:0] addr_11087_7;

Selector_2 s11087_7(wires_2771_6[3], addr_2771_6, addr_positional[44351:44348], addr_11087_7);

wire[31:0] addr_11088_7;

Selector_2 s11088_7(wires_2772_6[0], addr_2772_6, addr_positional[44355:44352], addr_11088_7);

wire[31:0] addr_11089_7;

Selector_2 s11089_7(wires_2772_6[1], addr_2772_6, addr_positional[44359:44356], addr_11089_7);

wire[31:0] addr_11090_7;

Selector_2 s11090_7(wires_2772_6[2], addr_2772_6, addr_positional[44363:44360], addr_11090_7);

wire[31:0] addr_11091_7;

Selector_2 s11091_7(wires_2772_6[3], addr_2772_6, addr_positional[44367:44364], addr_11091_7);

wire[31:0] addr_11092_7;

Selector_2 s11092_7(wires_2773_6[0], addr_2773_6, addr_positional[44371:44368], addr_11092_7);

wire[31:0] addr_11093_7;

Selector_2 s11093_7(wires_2773_6[1], addr_2773_6, addr_positional[44375:44372], addr_11093_7);

wire[31:0] addr_11094_7;

Selector_2 s11094_7(wires_2773_6[2], addr_2773_6, addr_positional[44379:44376], addr_11094_7);

wire[31:0] addr_11095_7;

Selector_2 s11095_7(wires_2773_6[3], addr_2773_6, addr_positional[44383:44380], addr_11095_7);

wire[31:0] addr_11096_7;

Selector_2 s11096_7(wires_2774_6[0], addr_2774_6, addr_positional[44387:44384], addr_11096_7);

wire[31:0] addr_11097_7;

Selector_2 s11097_7(wires_2774_6[1], addr_2774_6, addr_positional[44391:44388], addr_11097_7);

wire[31:0] addr_11098_7;

Selector_2 s11098_7(wires_2774_6[2], addr_2774_6, addr_positional[44395:44392], addr_11098_7);

wire[31:0] addr_11099_7;

Selector_2 s11099_7(wires_2774_6[3], addr_2774_6, addr_positional[44399:44396], addr_11099_7);

wire[31:0] addr_11100_7;

Selector_2 s11100_7(wires_2775_6[0], addr_2775_6, addr_positional[44403:44400], addr_11100_7);

wire[31:0] addr_11101_7;

Selector_2 s11101_7(wires_2775_6[1], addr_2775_6, addr_positional[44407:44404], addr_11101_7);

wire[31:0] addr_11102_7;

Selector_2 s11102_7(wires_2775_6[2], addr_2775_6, addr_positional[44411:44408], addr_11102_7);

wire[31:0] addr_11103_7;

Selector_2 s11103_7(wires_2775_6[3], addr_2775_6, addr_positional[44415:44412], addr_11103_7);

wire[31:0] addr_11104_7;

Selector_2 s11104_7(wires_2776_6[0], addr_2776_6, addr_positional[44419:44416], addr_11104_7);

wire[31:0] addr_11105_7;

Selector_2 s11105_7(wires_2776_6[1], addr_2776_6, addr_positional[44423:44420], addr_11105_7);

wire[31:0] addr_11106_7;

Selector_2 s11106_7(wires_2776_6[2], addr_2776_6, addr_positional[44427:44424], addr_11106_7);

wire[31:0] addr_11107_7;

Selector_2 s11107_7(wires_2776_6[3], addr_2776_6, addr_positional[44431:44428], addr_11107_7);

wire[31:0] addr_11108_7;

Selector_2 s11108_7(wires_2777_6[0], addr_2777_6, addr_positional[44435:44432], addr_11108_7);

wire[31:0] addr_11109_7;

Selector_2 s11109_7(wires_2777_6[1], addr_2777_6, addr_positional[44439:44436], addr_11109_7);

wire[31:0] addr_11110_7;

Selector_2 s11110_7(wires_2777_6[2], addr_2777_6, addr_positional[44443:44440], addr_11110_7);

wire[31:0] addr_11111_7;

Selector_2 s11111_7(wires_2777_6[3], addr_2777_6, addr_positional[44447:44444], addr_11111_7);

wire[31:0] addr_11112_7;

Selector_2 s11112_7(wires_2778_6[0], addr_2778_6, addr_positional[44451:44448], addr_11112_7);

wire[31:0] addr_11113_7;

Selector_2 s11113_7(wires_2778_6[1], addr_2778_6, addr_positional[44455:44452], addr_11113_7);

wire[31:0] addr_11114_7;

Selector_2 s11114_7(wires_2778_6[2], addr_2778_6, addr_positional[44459:44456], addr_11114_7);

wire[31:0] addr_11115_7;

Selector_2 s11115_7(wires_2778_6[3], addr_2778_6, addr_positional[44463:44460], addr_11115_7);

wire[31:0] addr_11116_7;

Selector_2 s11116_7(wires_2779_6[0], addr_2779_6, addr_positional[44467:44464], addr_11116_7);

wire[31:0] addr_11117_7;

Selector_2 s11117_7(wires_2779_6[1], addr_2779_6, addr_positional[44471:44468], addr_11117_7);

wire[31:0] addr_11118_7;

Selector_2 s11118_7(wires_2779_6[2], addr_2779_6, addr_positional[44475:44472], addr_11118_7);

wire[31:0] addr_11119_7;

Selector_2 s11119_7(wires_2779_6[3], addr_2779_6, addr_positional[44479:44476], addr_11119_7);

wire[31:0] addr_11120_7;

Selector_2 s11120_7(wires_2780_6[0], addr_2780_6, addr_positional[44483:44480], addr_11120_7);

wire[31:0] addr_11121_7;

Selector_2 s11121_7(wires_2780_6[1], addr_2780_6, addr_positional[44487:44484], addr_11121_7);

wire[31:0] addr_11122_7;

Selector_2 s11122_7(wires_2780_6[2], addr_2780_6, addr_positional[44491:44488], addr_11122_7);

wire[31:0] addr_11123_7;

Selector_2 s11123_7(wires_2780_6[3], addr_2780_6, addr_positional[44495:44492], addr_11123_7);

wire[31:0] addr_11124_7;

Selector_2 s11124_7(wires_2781_6[0], addr_2781_6, addr_positional[44499:44496], addr_11124_7);

wire[31:0] addr_11125_7;

Selector_2 s11125_7(wires_2781_6[1], addr_2781_6, addr_positional[44503:44500], addr_11125_7);

wire[31:0] addr_11126_7;

Selector_2 s11126_7(wires_2781_6[2], addr_2781_6, addr_positional[44507:44504], addr_11126_7);

wire[31:0] addr_11127_7;

Selector_2 s11127_7(wires_2781_6[3], addr_2781_6, addr_positional[44511:44508], addr_11127_7);

wire[31:0] addr_11128_7;

Selector_2 s11128_7(wires_2782_6[0], addr_2782_6, addr_positional[44515:44512], addr_11128_7);

wire[31:0] addr_11129_7;

Selector_2 s11129_7(wires_2782_6[1], addr_2782_6, addr_positional[44519:44516], addr_11129_7);

wire[31:0] addr_11130_7;

Selector_2 s11130_7(wires_2782_6[2], addr_2782_6, addr_positional[44523:44520], addr_11130_7);

wire[31:0] addr_11131_7;

Selector_2 s11131_7(wires_2782_6[3], addr_2782_6, addr_positional[44527:44524], addr_11131_7);

wire[31:0] addr_11132_7;

Selector_2 s11132_7(wires_2783_6[0], addr_2783_6, addr_positional[44531:44528], addr_11132_7);

wire[31:0] addr_11133_7;

Selector_2 s11133_7(wires_2783_6[1], addr_2783_6, addr_positional[44535:44532], addr_11133_7);

wire[31:0] addr_11134_7;

Selector_2 s11134_7(wires_2783_6[2], addr_2783_6, addr_positional[44539:44536], addr_11134_7);

wire[31:0] addr_11135_7;

Selector_2 s11135_7(wires_2783_6[3], addr_2783_6, addr_positional[44543:44540], addr_11135_7);

wire[31:0] addr_11136_7;

Selector_2 s11136_7(wires_2784_6[0], addr_2784_6, addr_positional[44547:44544], addr_11136_7);

wire[31:0] addr_11137_7;

Selector_2 s11137_7(wires_2784_6[1], addr_2784_6, addr_positional[44551:44548], addr_11137_7);

wire[31:0] addr_11138_7;

Selector_2 s11138_7(wires_2784_6[2], addr_2784_6, addr_positional[44555:44552], addr_11138_7);

wire[31:0] addr_11139_7;

Selector_2 s11139_7(wires_2784_6[3], addr_2784_6, addr_positional[44559:44556], addr_11139_7);

wire[31:0] addr_11140_7;

Selector_2 s11140_7(wires_2785_6[0], addr_2785_6, addr_positional[44563:44560], addr_11140_7);

wire[31:0] addr_11141_7;

Selector_2 s11141_7(wires_2785_6[1], addr_2785_6, addr_positional[44567:44564], addr_11141_7);

wire[31:0] addr_11142_7;

Selector_2 s11142_7(wires_2785_6[2], addr_2785_6, addr_positional[44571:44568], addr_11142_7);

wire[31:0] addr_11143_7;

Selector_2 s11143_7(wires_2785_6[3], addr_2785_6, addr_positional[44575:44572], addr_11143_7);

wire[31:0] addr_11144_7;

Selector_2 s11144_7(wires_2786_6[0], addr_2786_6, addr_positional[44579:44576], addr_11144_7);

wire[31:0] addr_11145_7;

Selector_2 s11145_7(wires_2786_6[1], addr_2786_6, addr_positional[44583:44580], addr_11145_7);

wire[31:0] addr_11146_7;

Selector_2 s11146_7(wires_2786_6[2], addr_2786_6, addr_positional[44587:44584], addr_11146_7);

wire[31:0] addr_11147_7;

Selector_2 s11147_7(wires_2786_6[3], addr_2786_6, addr_positional[44591:44588], addr_11147_7);

wire[31:0] addr_11148_7;

Selector_2 s11148_7(wires_2787_6[0], addr_2787_6, addr_positional[44595:44592], addr_11148_7);

wire[31:0] addr_11149_7;

Selector_2 s11149_7(wires_2787_6[1], addr_2787_6, addr_positional[44599:44596], addr_11149_7);

wire[31:0] addr_11150_7;

Selector_2 s11150_7(wires_2787_6[2], addr_2787_6, addr_positional[44603:44600], addr_11150_7);

wire[31:0] addr_11151_7;

Selector_2 s11151_7(wires_2787_6[3], addr_2787_6, addr_positional[44607:44604], addr_11151_7);

wire[31:0] addr_11152_7;

Selector_2 s11152_7(wires_2788_6[0], addr_2788_6, addr_positional[44611:44608], addr_11152_7);

wire[31:0] addr_11153_7;

Selector_2 s11153_7(wires_2788_6[1], addr_2788_6, addr_positional[44615:44612], addr_11153_7);

wire[31:0] addr_11154_7;

Selector_2 s11154_7(wires_2788_6[2], addr_2788_6, addr_positional[44619:44616], addr_11154_7);

wire[31:0] addr_11155_7;

Selector_2 s11155_7(wires_2788_6[3], addr_2788_6, addr_positional[44623:44620], addr_11155_7);

wire[31:0] addr_11156_7;

Selector_2 s11156_7(wires_2789_6[0], addr_2789_6, addr_positional[44627:44624], addr_11156_7);

wire[31:0] addr_11157_7;

Selector_2 s11157_7(wires_2789_6[1], addr_2789_6, addr_positional[44631:44628], addr_11157_7);

wire[31:0] addr_11158_7;

Selector_2 s11158_7(wires_2789_6[2], addr_2789_6, addr_positional[44635:44632], addr_11158_7);

wire[31:0] addr_11159_7;

Selector_2 s11159_7(wires_2789_6[3], addr_2789_6, addr_positional[44639:44636], addr_11159_7);

wire[31:0] addr_11160_7;

Selector_2 s11160_7(wires_2790_6[0], addr_2790_6, addr_positional[44643:44640], addr_11160_7);

wire[31:0] addr_11161_7;

Selector_2 s11161_7(wires_2790_6[1], addr_2790_6, addr_positional[44647:44644], addr_11161_7);

wire[31:0] addr_11162_7;

Selector_2 s11162_7(wires_2790_6[2], addr_2790_6, addr_positional[44651:44648], addr_11162_7);

wire[31:0] addr_11163_7;

Selector_2 s11163_7(wires_2790_6[3], addr_2790_6, addr_positional[44655:44652], addr_11163_7);

wire[31:0] addr_11164_7;

Selector_2 s11164_7(wires_2791_6[0], addr_2791_6, addr_positional[44659:44656], addr_11164_7);

wire[31:0] addr_11165_7;

Selector_2 s11165_7(wires_2791_6[1], addr_2791_6, addr_positional[44663:44660], addr_11165_7);

wire[31:0] addr_11166_7;

Selector_2 s11166_7(wires_2791_6[2], addr_2791_6, addr_positional[44667:44664], addr_11166_7);

wire[31:0] addr_11167_7;

Selector_2 s11167_7(wires_2791_6[3], addr_2791_6, addr_positional[44671:44668], addr_11167_7);

wire[31:0] addr_11168_7;

Selector_2 s11168_7(wires_2792_6[0], addr_2792_6, addr_positional[44675:44672], addr_11168_7);

wire[31:0] addr_11169_7;

Selector_2 s11169_7(wires_2792_6[1], addr_2792_6, addr_positional[44679:44676], addr_11169_7);

wire[31:0] addr_11170_7;

Selector_2 s11170_7(wires_2792_6[2], addr_2792_6, addr_positional[44683:44680], addr_11170_7);

wire[31:0] addr_11171_7;

Selector_2 s11171_7(wires_2792_6[3], addr_2792_6, addr_positional[44687:44684], addr_11171_7);

wire[31:0] addr_11172_7;

Selector_2 s11172_7(wires_2793_6[0], addr_2793_6, addr_positional[44691:44688], addr_11172_7);

wire[31:0] addr_11173_7;

Selector_2 s11173_7(wires_2793_6[1], addr_2793_6, addr_positional[44695:44692], addr_11173_7);

wire[31:0] addr_11174_7;

Selector_2 s11174_7(wires_2793_6[2], addr_2793_6, addr_positional[44699:44696], addr_11174_7);

wire[31:0] addr_11175_7;

Selector_2 s11175_7(wires_2793_6[3], addr_2793_6, addr_positional[44703:44700], addr_11175_7);

wire[31:0] addr_11176_7;

Selector_2 s11176_7(wires_2794_6[0], addr_2794_6, addr_positional[44707:44704], addr_11176_7);

wire[31:0] addr_11177_7;

Selector_2 s11177_7(wires_2794_6[1], addr_2794_6, addr_positional[44711:44708], addr_11177_7);

wire[31:0] addr_11178_7;

Selector_2 s11178_7(wires_2794_6[2], addr_2794_6, addr_positional[44715:44712], addr_11178_7);

wire[31:0] addr_11179_7;

Selector_2 s11179_7(wires_2794_6[3], addr_2794_6, addr_positional[44719:44716], addr_11179_7);

wire[31:0] addr_11180_7;

Selector_2 s11180_7(wires_2795_6[0], addr_2795_6, addr_positional[44723:44720], addr_11180_7);

wire[31:0] addr_11181_7;

Selector_2 s11181_7(wires_2795_6[1], addr_2795_6, addr_positional[44727:44724], addr_11181_7);

wire[31:0] addr_11182_7;

Selector_2 s11182_7(wires_2795_6[2], addr_2795_6, addr_positional[44731:44728], addr_11182_7);

wire[31:0] addr_11183_7;

Selector_2 s11183_7(wires_2795_6[3], addr_2795_6, addr_positional[44735:44732], addr_11183_7);

wire[31:0] addr_11184_7;

Selector_2 s11184_7(wires_2796_6[0], addr_2796_6, addr_positional[44739:44736], addr_11184_7);

wire[31:0] addr_11185_7;

Selector_2 s11185_7(wires_2796_6[1], addr_2796_6, addr_positional[44743:44740], addr_11185_7);

wire[31:0] addr_11186_7;

Selector_2 s11186_7(wires_2796_6[2], addr_2796_6, addr_positional[44747:44744], addr_11186_7);

wire[31:0] addr_11187_7;

Selector_2 s11187_7(wires_2796_6[3], addr_2796_6, addr_positional[44751:44748], addr_11187_7);

wire[31:0] addr_11188_7;

Selector_2 s11188_7(wires_2797_6[0], addr_2797_6, addr_positional[44755:44752], addr_11188_7);

wire[31:0] addr_11189_7;

Selector_2 s11189_7(wires_2797_6[1], addr_2797_6, addr_positional[44759:44756], addr_11189_7);

wire[31:0] addr_11190_7;

Selector_2 s11190_7(wires_2797_6[2], addr_2797_6, addr_positional[44763:44760], addr_11190_7);

wire[31:0] addr_11191_7;

Selector_2 s11191_7(wires_2797_6[3], addr_2797_6, addr_positional[44767:44764], addr_11191_7);

wire[31:0] addr_11192_7;

Selector_2 s11192_7(wires_2798_6[0], addr_2798_6, addr_positional[44771:44768], addr_11192_7);

wire[31:0] addr_11193_7;

Selector_2 s11193_7(wires_2798_6[1], addr_2798_6, addr_positional[44775:44772], addr_11193_7);

wire[31:0] addr_11194_7;

Selector_2 s11194_7(wires_2798_6[2], addr_2798_6, addr_positional[44779:44776], addr_11194_7);

wire[31:0] addr_11195_7;

Selector_2 s11195_7(wires_2798_6[3], addr_2798_6, addr_positional[44783:44780], addr_11195_7);

wire[31:0] addr_11196_7;

Selector_2 s11196_7(wires_2799_6[0], addr_2799_6, addr_positional[44787:44784], addr_11196_7);

wire[31:0] addr_11197_7;

Selector_2 s11197_7(wires_2799_6[1], addr_2799_6, addr_positional[44791:44788], addr_11197_7);

wire[31:0] addr_11198_7;

Selector_2 s11198_7(wires_2799_6[2], addr_2799_6, addr_positional[44795:44792], addr_11198_7);

wire[31:0] addr_11199_7;

Selector_2 s11199_7(wires_2799_6[3], addr_2799_6, addr_positional[44799:44796], addr_11199_7);

wire[31:0] addr_11200_7;

Selector_2 s11200_7(wires_2800_6[0], addr_2800_6, addr_positional[44803:44800], addr_11200_7);

wire[31:0] addr_11201_7;

Selector_2 s11201_7(wires_2800_6[1], addr_2800_6, addr_positional[44807:44804], addr_11201_7);

wire[31:0] addr_11202_7;

Selector_2 s11202_7(wires_2800_6[2], addr_2800_6, addr_positional[44811:44808], addr_11202_7);

wire[31:0] addr_11203_7;

Selector_2 s11203_7(wires_2800_6[3], addr_2800_6, addr_positional[44815:44812], addr_11203_7);

wire[31:0] addr_11204_7;

Selector_2 s11204_7(wires_2801_6[0], addr_2801_6, addr_positional[44819:44816], addr_11204_7);

wire[31:0] addr_11205_7;

Selector_2 s11205_7(wires_2801_6[1], addr_2801_6, addr_positional[44823:44820], addr_11205_7);

wire[31:0] addr_11206_7;

Selector_2 s11206_7(wires_2801_6[2], addr_2801_6, addr_positional[44827:44824], addr_11206_7);

wire[31:0] addr_11207_7;

Selector_2 s11207_7(wires_2801_6[3], addr_2801_6, addr_positional[44831:44828], addr_11207_7);

wire[31:0] addr_11208_7;

Selector_2 s11208_7(wires_2802_6[0], addr_2802_6, addr_positional[44835:44832], addr_11208_7);

wire[31:0] addr_11209_7;

Selector_2 s11209_7(wires_2802_6[1], addr_2802_6, addr_positional[44839:44836], addr_11209_7);

wire[31:0] addr_11210_7;

Selector_2 s11210_7(wires_2802_6[2], addr_2802_6, addr_positional[44843:44840], addr_11210_7);

wire[31:0] addr_11211_7;

Selector_2 s11211_7(wires_2802_6[3], addr_2802_6, addr_positional[44847:44844], addr_11211_7);

wire[31:0] addr_11212_7;

Selector_2 s11212_7(wires_2803_6[0], addr_2803_6, addr_positional[44851:44848], addr_11212_7);

wire[31:0] addr_11213_7;

Selector_2 s11213_7(wires_2803_6[1], addr_2803_6, addr_positional[44855:44852], addr_11213_7);

wire[31:0] addr_11214_7;

Selector_2 s11214_7(wires_2803_6[2], addr_2803_6, addr_positional[44859:44856], addr_11214_7);

wire[31:0] addr_11215_7;

Selector_2 s11215_7(wires_2803_6[3], addr_2803_6, addr_positional[44863:44860], addr_11215_7);

wire[31:0] addr_11216_7;

Selector_2 s11216_7(wires_2804_6[0], addr_2804_6, addr_positional[44867:44864], addr_11216_7);

wire[31:0] addr_11217_7;

Selector_2 s11217_7(wires_2804_6[1], addr_2804_6, addr_positional[44871:44868], addr_11217_7);

wire[31:0] addr_11218_7;

Selector_2 s11218_7(wires_2804_6[2], addr_2804_6, addr_positional[44875:44872], addr_11218_7);

wire[31:0] addr_11219_7;

Selector_2 s11219_7(wires_2804_6[3], addr_2804_6, addr_positional[44879:44876], addr_11219_7);

wire[31:0] addr_11220_7;

Selector_2 s11220_7(wires_2805_6[0], addr_2805_6, addr_positional[44883:44880], addr_11220_7);

wire[31:0] addr_11221_7;

Selector_2 s11221_7(wires_2805_6[1], addr_2805_6, addr_positional[44887:44884], addr_11221_7);

wire[31:0] addr_11222_7;

Selector_2 s11222_7(wires_2805_6[2], addr_2805_6, addr_positional[44891:44888], addr_11222_7);

wire[31:0] addr_11223_7;

Selector_2 s11223_7(wires_2805_6[3], addr_2805_6, addr_positional[44895:44892], addr_11223_7);

wire[31:0] addr_11224_7;

Selector_2 s11224_7(wires_2806_6[0], addr_2806_6, addr_positional[44899:44896], addr_11224_7);

wire[31:0] addr_11225_7;

Selector_2 s11225_7(wires_2806_6[1], addr_2806_6, addr_positional[44903:44900], addr_11225_7);

wire[31:0] addr_11226_7;

Selector_2 s11226_7(wires_2806_6[2], addr_2806_6, addr_positional[44907:44904], addr_11226_7);

wire[31:0] addr_11227_7;

Selector_2 s11227_7(wires_2806_6[3], addr_2806_6, addr_positional[44911:44908], addr_11227_7);

wire[31:0] addr_11228_7;

Selector_2 s11228_7(wires_2807_6[0], addr_2807_6, addr_positional[44915:44912], addr_11228_7);

wire[31:0] addr_11229_7;

Selector_2 s11229_7(wires_2807_6[1], addr_2807_6, addr_positional[44919:44916], addr_11229_7);

wire[31:0] addr_11230_7;

Selector_2 s11230_7(wires_2807_6[2], addr_2807_6, addr_positional[44923:44920], addr_11230_7);

wire[31:0] addr_11231_7;

Selector_2 s11231_7(wires_2807_6[3], addr_2807_6, addr_positional[44927:44924], addr_11231_7);

wire[31:0] addr_11232_7;

Selector_2 s11232_7(wires_2808_6[0], addr_2808_6, addr_positional[44931:44928], addr_11232_7);

wire[31:0] addr_11233_7;

Selector_2 s11233_7(wires_2808_6[1], addr_2808_6, addr_positional[44935:44932], addr_11233_7);

wire[31:0] addr_11234_7;

Selector_2 s11234_7(wires_2808_6[2], addr_2808_6, addr_positional[44939:44936], addr_11234_7);

wire[31:0] addr_11235_7;

Selector_2 s11235_7(wires_2808_6[3], addr_2808_6, addr_positional[44943:44940], addr_11235_7);

wire[31:0] addr_11236_7;

Selector_2 s11236_7(wires_2809_6[0], addr_2809_6, addr_positional[44947:44944], addr_11236_7);

wire[31:0] addr_11237_7;

Selector_2 s11237_7(wires_2809_6[1], addr_2809_6, addr_positional[44951:44948], addr_11237_7);

wire[31:0] addr_11238_7;

Selector_2 s11238_7(wires_2809_6[2], addr_2809_6, addr_positional[44955:44952], addr_11238_7);

wire[31:0] addr_11239_7;

Selector_2 s11239_7(wires_2809_6[3], addr_2809_6, addr_positional[44959:44956], addr_11239_7);

wire[31:0] addr_11240_7;

Selector_2 s11240_7(wires_2810_6[0], addr_2810_6, addr_positional[44963:44960], addr_11240_7);

wire[31:0] addr_11241_7;

Selector_2 s11241_7(wires_2810_6[1], addr_2810_6, addr_positional[44967:44964], addr_11241_7);

wire[31:0] addr_11242_7;

Selector_2 s11242_7(wires_2810_6[2], addr_2810_6, addr_positional[44971:44968], addr_11242_7);

wire[31:0] addr_11243_7;

Selector_2 s11243_7(wires_2810_6[3], addr_2810_6, addr_positional[44975:44972], addr_11243_7);

wire[31:0] addr_11244_7;

Selector_2 s11244_7(wires_2811_6[0], addr_2811_6, addr_positional[44979:44976], addr_11244_7);

wire[31:0] addr_11245_7;

Selector_2 s11245_7(wires_2811_6[1], addr_2811_6, addr_positional[44983:44980], addr_11245_7);

wire[31:0] addr_11246_7;

Selector_2 s11246_7(wires_2811_6[2], addr_2811_6, addr_positional[44987:44984], addr_11246_7);

wire[31:0] addr_11247_7;

Selector_2 s11247_7(wires_2811_6[3], addr_2811_6, addr_positional[44991:44988], addr_11247_7);

wire[31:0] addr_11248_7;

Selector_2 s11248_7(wires_2812_6[0], addr_2812_6, addr_positional[44995:44992], addr_11248_7);

wire[31:0] addr_11249_7;

Selector_2 s11249_7(wires_2812_6[1], addr_2812_6, addr_positional[44999:44996], addr_11249_7);

wire[31:0] addr_11250_7;

Selector_2 s11250_7(wires_2812_6[2], addr_2812_6, addr_positional[45003:45000], addr_11250_7);

wire[31:0] addr_11251_7;

Selector_2 s11251_7(wires_2812_6[3], addr_2812_6, addr_positional[45007:45004], addr_11251_7);

wire[31:0] addr_11252_7;

Selector_2 s11252_7(wires_2813_6[0], addr_2813_6, addr_positional[45011:45008], addr_11252_7);

wire[31:0] addr_11253_7;

Selector_2 s11253_7(wires_2813_6[1], addr_2813_6, addr_positional[45015:45012], addr_11253_7);

wire[31:0] addr_11254_7;

Selector_2 s11254_7(wires_2813_6[2], addr_2813_6, addr_positional[45019:45016], addr_11254_7);

wire[31:0] addr_11255_7;

Selector_2 s11255_7(wires_2813_6[3], addr_2813_6, addr_positional[45023:45020], addr_11255_7);

wire[31:0] addr_11256_7;

Selector_2 s11256_7(wires_2814_6[0], addr_2814_6, addr_positional[45027:45024], addr_11256_7);

wire[31:0] addr_11257_7;

Selector_2 s11257_7(wires_2814_6[1], addr_2814_6, addr_positional[45031:45028], addr_11257_7);

wire[31:0] addr_11258_7;

Selector_2 s11258_7(wires_2814_6[2], addr_2814_6, addr_positional[45035:45032], addr_11258_7);

wire[31:0] addr_11259_7;

Selector_2 s11259_7(wires_2814_6[3], addr_2814_6, addr_positional[45039:45036], addr_11259_7);

wire[31:0] addr_11260_7;

Selector_2 s11260_7(wires_2815_6[0], addr_2815_6, addr_positional[45043:45040], addr_11260_7);

wire[31:0] addr_11261_7;

Selector_2 s11261_7(wires_2815_6[1], addr_2815_6, addr_positional[45047:45044], addr_11261_7);

wire[31:0] addr_11262_7;

Selector_2 s11262_7(wires_2815_6[2], addr_2815_6, addr_positional[45051:45048], addr_11262_7);

wire[31:0] addr_11263_7;

Selector_2 s11263_7(wires_2815_6[3], addr_2815_6, addr_positional[45055:45052], addr_11263_7);

wire[31:0] addr_11264_7;

Selector_2 s11264_7(wires_2816_6[0], addr_2816_6, addr_positional[45059:45056], addr_11264_7);

wire[31:0] addr_11265_7;

Selector_2 s11265_7(wires_2816_6[1], addr_2816_6, addr_positional[45063:45060], addr_11265_7);

wire[31:0] addr_11266_7;

Selector_2 s11266_7(wires_2816_6[2], addr_2816_6, addr_positional[45067:45064], addr_11266_7);

wire[31:0] addr_11267_7;

Selector_2 s11267_7(wires_2816_6[3], addr_2816_6, addr_positional[45071:45068], addr_11267_7);

wire[31:0] addr_11268_7;

Selector_2 s11268_7(wires_2817_6[0], addr_2817_6, addr_positional[45075:45072], addr_11268_7);

wire[31:0] addr_11269_7;

Selector_2 s11269_7(wires_2817_6[1], addr_2817_6, addr_positional[45079:45076], addr_11269_7);

wire[31:0] addr_11270_7;

Selector_2 s11270_7(wires_2817_6[2], addr_2817_6, addr_positional[45083:45080], addr_11270_7);

wire[31:0] addr_11271_7;

Selector_2 s11271_7(wires_2817_6[3], addr_2817_6, addr_positional[45087:45084], addr_11271_7);

wire[31:0] addr_11272_7;

Selector_2 s11272_7(wires_2818_6[0], addr_2818_6, addr_positional[45091:45088], addr_11272_7);

wire[31:0] addr_11273_7;

Selector_2 s11273_7(wires_2818_6[1], addr_2818_6, addr_positional[45095:45092], addr_11273_7);

wire[31:0] addr_11274_7;

Selector_2 s11274_7(wires_2818_6[2], addr_2818_6, addr_positional[45099:45096], addr_11274_7);

wire[31:0] addr_11275_7;

Selector_2 s11275_7(wires_2818_6[3], addr_2818_6, addr_positional[45103:45100], addr_11275_7);

wire[31:0] addr_11276_7;

Selector_2 s11276_7(wires_2819_6[0], addr_2819_6, addr_positional[45107:45104], addr_11276_7);

wire[31:0] addr_11277_7;

Selector_2 s11277_7(wires_2819_6[1], addr_2819_6, addr_positional[45111:45108], addr_11277_7);

wire[31:0] addr_11278_7;

Selector_2 s11278_7(wires_2819_6[2], addr_2819_6, addr_positional[45115:45112], addr_11278_7);

wire[31:0] addr_11279_7;

Selector_2 s11279_7(wires_2819_6[3], addr_2819_6, addr_positional[45119:45116], addr_11279_7);

wire[31:0] addr_11280_7;

Selector_2 s11280_7(wires_2820_6[0], addr_2820_6, addr_positional[45123:45120], addr_11280_7);

wire[31:0] addr_11281_7;

Selector_2 s11281_7(wires_2820_6[1], addr_2820_6, addr_positional[45127:45124], addr_11281_7);

wire[31:0] addr_11282_7;

Selector_2 s11282_7(wires_2820_6[2], addr_2820_6, addr_positional[45131:45128], addr_11282_7);

wire[31:0] addr_11283_7;

Selector_2 s11283_7(wires_2820_6[3], addr_2820_6, addr_positional[45135:45132], addr_11283_7);

wire[31:0] addr_11284_7;

Selector_2 s11284_7(wires_2821_6[0], addr_2821_6, addr_positional[45139:45136], addr_11284_7);

wire[31:0] addr_11285_7;

Selector_2 s11285_7(wires_2821_6[1], addr_2821_6, addr_positional[45143:45140], addr_11285_7);

wire[31:0] addr_11286_7;

Selector_2 s11286_7(wires_2821_6[2], addr_2821_6, addr_positional[45147:45144], addr_11286_7);

wire[31:0] addr_11287_7;

Selector_2 s11287_7(wires_2821_6[3], addr_2821_6, addr_positional[45151:45148], addr_11287_7);

wire[31:0] addr_11288_7;

Selector_2 s11288_7(wires_2822_6[0], addr_2822_6, addr_positional[45155:45152], addr_11288_7);

wire[31:0] addr_11289_7;

Selector_2 s11289_7(wires_2822_6[1], addr_2822_6, addr_positional[45159:45156], addr_11289_7);

wire[31:0] addr_11290_7;

Selector_2 s11290_7(wires_2822_6[2], addr_2822_6, addr_positional[45163:45160], addr_11290_7);

wire[31:0] addr_11291_7;

Selector_2 s11291_7(wires_2822_6[3], addr_2822_6, addr_positional[45167:45164], addr_11291_7);

wire[31:0] addr_11292_7;

Selector_2 s11292_7(wires_2823_6[0], addr_2823_6, addr_positional[45171:45168], addr_11292_7);

wire[31:0] addr_11293_7;

Selector_2 s11293_7(wires_2823_6[1], addr_2823_6, addr_positional[45175:45172], addr_11293_7);

wire[31:0] addr_11294_7;

Selector_2 s11294_7(wires_2823_6[2], addr_2823_6, addr_positional[45179:45176], addr_11294_7);

wire[31:0] addr_11295_7;

Selector_2 s11295_7(wires_2823_6[3], addr_2823_6, addr_positional[45183:45180], addr_11295_7);

wire[31:0] addr_11296_7;

Selector_2 s11296_7(wires_2824_6[0], addr_2824_6, addr_positional[45187:45184], addr_11296_7);

wire[31:0] addr_11297_7;

Selector_2 s11297_7(wires_2824_6[1], addr_2824_6, addr_positional[45191:45188], addr_11297_7);

wire[31:0] addr_11298_7;

Selector_2 s11298_7(wires_2824_6[2], addr_2824_6, addr_positional[45195:45192], addr_11298_7);

wire[31:0] addr_11299_7;

Selector_2 s11299_7(wires_2824_6[3], addr_2824_6, addr_positional[45199:45196], addr_11299_7);

wire[31:0] addr_11300_7;

Selector_2 s11300_7(wires_2825_6[0], addr_2825_6, addr_positional[45203:45200], addr_11300_7);

wire[31:0] addr_11301_7;

Selector_2 s11301_7(wires_2825_6[1], addr_2825_6, addr_positional[45207:45204], addr_11301_7);

wire[31:0] addr_11302_7;

Selector_2 s11302_7(wires_2825_6[2], addr_2825_6, addr_positional[45211:45208], addr_11302_7);

wire[31:0] addr_11303_7;

Selector_2 s11303_7(wires_2825_6[3], addr_2825_6, addr_positional[45215:45212], addr_11303_7);

wire[31:0] addr_11304_7;

Selector_2 s11304_7(wires_2826_6[0], addr_2826_6, addr_positional[45219:45216], addr_11304_7);

wire[31:0] addr_11305_7;

Selector_2 s11305_7(wires_2826_6[1], addr_2826_6, addr_positional[45223:45220], addr_11305_7);

wire[31:0] addr_11306_7;

Selector_2 s11306_7(wires_2826_6[2], addr_2826_6, addr_positional[45227:45224], addr_11306_7);

wire[31:0] addr_11307_7;

Selector_2 s11307_7(wires_2826_6[3], addr_2826_6, addr_positional[45231:45228], addr_11307_7);

wire[31:0] addr_11308_7;

Selector_2 s11308_7(wires_2827_6[0], addr_2827_6, addr_positional[45235:45232], addr_11308_7);

wire[31:0] addr_11309_7;

Selector_2 s11309_7(wires_2827_6[1], addr_2827_6, addr_positional[45239:45236], addr_11309_7);

wire[31:0] addr_11310_7;

Selector_2 s11310_7(wires_2827_6[2], addr_2827_6, addr_positional[45243:45240], addr_11310_7);

wire[31:0] addr_11311_7;

Selector_2 s11311_7(wires_2827_6[3], addr_2827_6, addr_positional[45247:45244], addr_11311_7);

wire[31:0] addr_11312_7;

Selector_2 s11312_7(wires_2828_6[0], addr_2828_6, addr_positional[45251:45248], addr_11312_7);

wire[31:0] addr_11313_7;

Selector_2 s11313_7(wires_2828_6[1], addr_2828_6, addr_positional[45255:45252], addr_11313_7);

wire[31:0] addr_11314_7;

Selector_2 s11314_7(wires_2828_6[2], addr_2828_6, addr_positional[45259:45256], addr_11314_7);

wire[31:0] addr_11315_7;

Selector_2 s11315_7(wires_2828_6[3], addr_2828_6, addr_positional[45263:45260], addr_11315_7);

wire[31:0] addr_11316_7;

Selector_2 s11316_7(wires_2829_6[0], addr_2829_6, addr_positional[45267:45264], addr_11316_7);

wire[31:0] addr_11317_7;

Selector_2 s11317_7(wires_2829_6[1], addr_2829_6, addr_positional[45271:45268], addr_11317_7);

wire[31:0] addr_11318_7;

Selector_2 s11318_7(wires_2829_6[2], addr_2829_6, addr_positional[45275:45272], addr_11318_7);

wire[31:0] addr_11319_7;

Selector_2 s11319_7(wires_2829_6[3], addr_2829_6, addr_positional[45279:45276], addr_11319_7);

wire[31:0] addr_11320_7;

Selector_2 s11320_7(wires_2830_6[0], addr_2830_6, addr_positional[45283:45280], addr_11320_7);

wire[31:0] addr_11321_7;

Selector_2 s11321_7(wires_2830_6[1], addr_2830_6, addr_positional[45287:45284], addr_11321_7);

wire[31:0] addr_11322_7;

Selector_2 s11322_7(wires_2830_6[2], addr_2830_6, addr_positional[45291:45288], addr_11322_7);

wire[31:0] addr_11323_7;

Selector_2 s11323_7(wires_2830_6[3], addr_2830_6, addr_positional[45295:45292], addr_11323_7);

wire[31:0] addr_11324_7;

Selector_2 s11324_7(wires_2831_6[0], addr_2831_6, addr_positional[45299:45296], addr_11324_7);

wire[31:0] addr_11325_7;

Selector_2 s11325_7(wires_2831_6[1], addr_2831_6, addr_positional[45303:45300], addr_11325_7);

wire[31:0] addr_11326_7;

Selector_2 s11326_7(wires_2831_6[2], addr_2831_6, addr_positional[45307:45304], addr_11326_7);

wire[31:0] addr_11327_7;

Selector_2 s11327_7(wires_2831_6[3], addr_2831_6, addr_positional[45311:45308], addr_11327_7);

wire[31:0] addr_11328_7;

Selector_2 s11328_7(wires_2832_6[0], addr_2832_6, addr_positional[45315:45312], addr_11328_7);

wire[31:0] addr_11329_7;

Selector_2 s11329_7(wires_2832_6[1], addr_2832_6, addr_positional[45319:45316], addr_11329_7);

wire[31:0] addr_11330_7;

Selector_2 s11330_7(wires_2832_6[2], addr_2832_6, addr_positional[45323:45320], addr_11330_7);

wire[31:0] addr_11331_7;

Selector_2 s11331_7(wires_2832_6[3], addr_2832_6, addr_positional[45327:45324], addr_11331_7);

wire[31:0] addr_11332_7;

Selector_2 s11332_7(wires_2833_6[0], addr_2833_6, addr_positional[45331:45328], addr_11332_7);

wire[31:0] addr_11333_7;

Selector_2 s11333_7(wires_2833_6[1], addr_2833_6, addr_positional[45335:45332], addr_11333_7);

wire[31:0] addr_11334_7;

Selector_2 s11334_7(wires_2833_6[2], addr_2833_6, addr_positional[45339:45336], addr_11334_7);

wire[31:0] addr_11335_7;

Selector_2 s11335_7(wires_2833_6[3], addr_2833_6, addr_positional[45343:45340], addr_11335_7);

wire[31:0] addr_11336_7;

Selector_2 s11336_7(wires_2834_6[0], addr_2834_6, addr_positional[45347:45344], addr_11336_7);

wire[31:0] addr_11337_7;

Selector_2 s11337_7(wires_2834_6[1], addr_2834_6, addr_positional[45351:45348], addr_11337_7);

wire[31:0] addr_11338_7;

Selector_2 s11338_7(wires_2834_6[2], addr_2834_6, addr_positional[45355:45352], addr_11338_7);

wire[31:0] addr_11339_7;

Selector_2 s11339_7(wires_2834_6[3], addr_2834_6, addr_positional[45359:45356], addr_11339_7);

wire[31:0] addr_11340_7;

Selector_2 s11340_7(wires_2835_6[0], addr_2835_6, addr_positional[45363:45360], addr_11340_7);

wire[31:0] addr_11341_7;

Selector_2 s11341_7(wires_2835_6[1], addr_2835_6, addr_positional[45367:45364], addr_11341_7);

wire[31:0] addr_11342_7;

Selector_2 s11342_7(wires_2835_6[2], addr_2835_6, addr_positional[45371:45368], addr_11342_7);

wire[31:0] addr_11343_7;

Selector_2 s11343_7(wires_2835_6[3], addr_2835_6, addr_positional[45375:45372], addr_11343_7);

wire[31:0] addr_11344_7;

Selector_2 s11344_7(wires_2836_6[0], addr_2836_6, addr_positional[45379:45376], addr_11344_7);

wire[31:0] addr_11345_7;

Selector_2 s11345_7(wires_2836_6[1], addr_2836_6, addr_positional[45383:45380], addr_11345_7);

wire[31:0] addr_11346_7;

Selector_2 s11346_7(wires_2836_6[2], addr_2836_6, addr_positional[45387:45384], addr_11346_7);

wire[31:0] addr_11347_7;

Selector_2 s11347_7(wires_2836_6[3], addr_2836_6, addr_positional[45391:45388], addr_11347_7);

wire[31:0] addr_11348_7;

Selector_2 s11348_7(wires_2837_6[0], addr_2837_6, addr_positional[45395:45392], addr_11348_7);

wire[31:0] addr_11349_7;

Selector_2 s11349_7(wires_2837_6[1], addr_2837_6, addr_positional[45399:45396], addr_11349_7);

wire[31:0] addr_11350_7;

Selector_2 s11350_7(wires_2837_6[2], addr_2837_6, addr_positional[45403:45400], addr_11350_7);

wire[31:0] addr_11351_7;

Selector_2 s11351_7(wires_2837_6[3], addr_2837_6, addr_positional[45407:45404], addr_11351_7);

wire[31:0] addr_11352_7;

Selector_2 s11352_7(wires_2838_6[0], addr_2838_6, addr_positional[45411:45408], addr_11352_7);

wire[31:0] addr_11353_7;

Selector_2 s11353_7(wires_2838_6[1], addr_2838_6, addr_positional[45415:45412], addr_11353_7);

wire[31:0] addr_11354_7;

Selector_2 s11354_7(wires_2838_6[2], addr_2838_6, addr_positional[45419:45416], addr_11354_7);

wire[31:0] addr_11355_7;

Selector_2 s11355_7(wires_2838_6[3], addr_2838_6, addr_positional[45423:45420], addr_11355_7);

wire[31:0] addr_11356_7;

Selector_2 s11356_7(wires_2839_6[0], addr_2839_6, addr_positional[45427:45424], addr_11356_7);

wire[31:0] addr_11357_7;

Selector_2 s11357_7(wires_2839_6[1], addr_2839_6, addr_positional[45431:45428], addr_11357_7);

wire[31:0] addr_11358_7;

Selector_2 s11358_7(wires_2839_6[2], addr_2839_6, addr_positional[45435:45432], addr_11358_7);

wire[31:0] addr_11359_7;

Selector_2 s11359_7(wires_2839_6[3], addr_2839_6, addr_positional[45439:45436], addr_11359_7);

wire[31:0] addr_11360_7;

Selector_2 s11360_7(wires_2840_6[0], addr_2840_6, addr_positional[45443:45440], addr_11360_7);

wire[31:0] addr_11361_7;

Selector_2 s11361_7(wires_2840_6[1], addr_2840_6, addr_positional[45447:45444], addr_11361_7);

wire[31:0] addr_11362_7;

Selector_2 s11362_7(wires_2840_6[2], addr_2840_6, addr_positional[45451:45448], addr_11362_7);

wire[31:0] addr_11363_7;

Selector_2 s11363_7(wires_2840_6[3], addr_2840_6, addr_positional[45455:45452], addr_11363_7);

wire[31:0] addr_11364_7;

Selector_2 s11364_7(wires_2841_6[0], addr_2841_6, addr_positional[45459:45456], addr_11364_7);

wire[31:0] addr_11365_7;

Selector_2 s11365_7(wires_2841_6[1], addr_2841_6, addr_positional[45463:45460], addr_11365_7);

wire[31:0] addr_11366_7;

Selector_2 s11366_7(wires_2841_6[2], addr_2841_6, addr_positional[45467:45464], addr_11366_7);

wire[31:0] addr_11367_7;

Selector_2 s11367_7(wires_2841_6[3], addr_2841_6, addr_positional[45471:45468], addr_11367_7);

wire[31:0] addr_11368_7;

Selector_2 s11368_7(wires_2842_6[0], addr_2842_6, addr_positional[45475:45472], addr_11368_7);

wire[31:0] addr_11369_7;

Selector_2 s11369_7(wires_2842_6[1], addr_2842_6, addr_positional[45479:45476], addr_11369_7);

wire[31:0] addr_11370_7;

Selector_2 s11370_7(wires_2842_6[2], addr_2842_6, addr_positional[45483:45480], addr_11370_7);

wire[31:0] addr_11371_7;

Selector_2 s11371_7(wires_2842_6[3], addr_2842_6, addr_positional[45487:45484], addr_11371_7);

wire[31:0] addr_11372_7;

Selector_2 s11372_7(wires_2843_6[0], addr_2843_6, addr_positional[45491:45488], addr_11372_7);

wire[31:0] addr_11373_7;

Selector_2 s11373_7(wires_2843_6[1], addr_2843_6, addr_positional[45495:45492], addr_11373_7);

wire[31:0] addr_11374_7;

Selector_2 s11374_7(wires_2843_6[2], addr_2843_6, addr_positional[45499:45496], addr_11374_7);

wire[31:0] addr_11375_7;

Selector_2 s11375_7(wires_2843_6[3], addr_2843_6, addr_positional[45503:45500], addr_11375_7);

wire[31:0] addr_11376_7;

Selector_2 s11376_7(wires_2844_6[0], addr_2844_6, addr_positional[45507:45504], addr_11376_7);

wire[31:0] addr_11377_7;

Selector_2 s11377_7(wires_2844_6[1], addr_2844_6, addr_positional[45511:45508], addr_11377_7);

wire[31:0] addr_11378_7;

Selector_2 s11378_7(wires_2844_6[2], addr_2844_6, addr_positional[45515:45512], addr_11378_7);

wire[31:0] addr_11379_7;

Selector_2 s11379_7(wires_2844_6[3], addr_2844_6, addr_positional[45519:45516], addr_11379_7);

wire[31:0] addr_11380_7;

Selector_2 s11380_7(wires_2845_6[0], addr_2845_6, addr_positional[45523:45520], addr_11380_7);

wire[31:0] addr_11381_7;

Selector_2 s11381_7(wires_2845_6[1], addr_2845_6, addr_positional[45527:45524], addr_11381_7);

wire[31:0] addr_11382_7;

Selector_2 s11382_7(wires_2845_6[2], addr_2845_6, addr_positional[45531:45528], addr_11382_7);

wire[31:0] addr_11383_7;

Selector_2 s11383_7(wires_2845_6[3], addr_2845_6, addr_positional[45535:45532], addr_11383_7);

wire[31:0] addr_11384_7;

Selector_2 s11384_7(wires_2846_6[0], addr_2846_6, addr_positional[45539:45536], addr_11384_7);

wire[31:0] addr_11385_7;

Selector_2 s11385_7(wires_2846_6[1], addr_2846_6, addr_positional[45543:45540], addr_11385_7);

wire[31:0] addr_11386_7;

Selector_2 s11386_7(wires_2846_6[2], addr_2846_6, addr_positional[45547:45544], addr_11386_7);

wire[31:0] addr_11387_7;

Selector_2 s11387_7(wires_2846_6[3], addr_2846_6, addr_positional[45551:45548], addr_11387_7);

wire[31:0] addr_11388_7;

Selector_2 s11388_7(wires_2847_6[0], addr_2847_6, addr_positional[45555:45552], addr_11388_7);

wire[31:0] addr_11389_7;

Selector_2 s11389_7(wires_2847_6[1], addr_2847_6, addr_positional[45559:45556], addr_11389_7);

wire[31:0] addr_11390_7;

Selector_2 s11390_7(wires_2847_6[2], addr_2847_6, addr_positional[45563:45560], addr_11390_7);

wire[31:0] addr_11391_7;

Selector_2 s11391_7(wires_2847_6[3], addr_2847_6, addr_positional[45567:45564], addr_11391_7);

wire[31:0] addr_11392_7;

Selector_2 s11392_7(wires_2848_6[0], addr_2848_6, addr_positional[45571:45568], addr_11392_7);

wire[31:0] addr_11393_7;

Selector_2 s11393_7(wires_2848_6[1], addr_2848_6, addr_positional[45575:45572], addr_11393_7);

wire[31:0] addr_11394_7;

Selector_2 s11394_7(wires_2848_6[2], addr_2848_6, addr_positional[45579:45576], addr_11394_7);

wire[31:0] addr_11395_7;

Selector_2 s11395_7(wires_2848_6[3], addr_2848_6, addr_positional[45583:45580], addr_11395_7);

wire[31:0] addr_11396_7;

Selector_2 s11396_7(wires_2849_6[0], addr_2849_6, addr_positional[45587:45584], addr_11396_7);

wire[31:0] addr_11397_7;

Selector_2 s11397_7(wires_2849_6[1], addr_2849_6, addr_positional[45591:45588], addr_11397_7);

wire[31:0] addr_11398_7;

Selector_2 s11398_7(wires_2849_6[2], addr_2849_6, addr_positional[45595:45592], addr_11398_7);

wire[31:0] addr_11399_7;

Selector_2 s11399_7(wires_2849_6[3], addr_2849_6, addr_positional[45599:45596], addr_11399_7);

wire[31:0] addr_11400_7;

Selector_2 s11400_7(wires_2850_6[0], addr_2850_6, addr_positional[45603:45600], addr_11400_7);

wire[31:0] addr_11401_7;

Selector_2 s11401_7(wires_2850_6[1], addr_2850_6, addr_positional[45607:45604], addr_11401_7);

wire[31:0] addr_11402_7;

Selector_2 s11402_7(wires_2850_6[2], addr_2850_6, addr_positional[45611:45608], addr_11402_7);

wire[31:0] addr_11403_7;

Selector_2 s11403_7(wires_2850_6[3], addr_2850_6, addr_positional[45615:45612], addr_11403_7);

wire[31:0] addr_11404_7;

Selector_2 s11404_7(wires_2851_6[0], addr_2851_6, addr_positional[45619:45616], addr_11404_7);

wire[31:0] addr_11405_7;

Selector_2 s11405_7(wires_2851_6[1], addr_2851_6, addr_positional[45623:45620], addr_11405_7);

wire[31:0] addr_11406_7;

Selector_2 s11406_7(wires_2851_6[2], addr_2851_6, addr_positional[45627:45624], addr_11406_7);

wire[31:0] addr_11407_7;

Selector_2 s11407_7(wires_2851_6[3], addr_2851_6, addr_positional[45631:45628], addr_11407_7);

wire[31:0] addr_11408_7;

Selector_2 s11408_7(wires_2852_6[0], addr_2852_6, addr_positional[45635:45632], addr_11408_7);

wire[31:0] addr_11409_7;

Selector_2 s11409_7(wires_2852_6[1], addr_2852_6, addr_positional[45639:45636], addr_11409_7);

wire[31:0] addr_11410_7;

Selector_2 s11410_7(wires_2852_6[2], addr_2852_6, addr_positional[45643:45640], addr_11410_7);

wire[31:0] addr_11411_7;

Selector_2 s11411_7(wires_2852_6[3], addr_2852_6, addr_positional[45647:45644], addr_11411_7);

wire[31:0] addr_11412_7;

Selector_2 s11412_7(wires_2853_6[0], addr_2853_6, addr_positional[45651:45648], addr_11412_7);

wire[31:0] addr_11413_7;

Selector_2 s11413_7(wires_2853_6[1], addr_2853_6, addr_positional[45655:45652], addr_11413_7);

wire[31:0] addr_11414_7;

Selector_2 s11414_7(wires_2853_6[2], addr_2853_6, addr_positional[45659:45656], addr_11414_7);

wire[31:0] addr_11415_7;

Selector_2 s11415_7(wires_2853_6[3], addr_2853_6, addr_positional[45663:45660], addr_11415_7);

wire[31:0] addr_11416_7;

Selector_2 s11416_7(wires_2854_6[0], addr_2854_6, addr_positional[45667:45664], addr_11416_7);

wire[31:0] addr_11417_7;

Selector_2 s11417_7(wires_2854_6[1], addr_2854_6, addr_positional[45671:45668], addr_11417_7);

wire[31:0] addr_11418_7;

Selector_2 s11418_7(wires_2854_6[2], addr_2854_6, addr_positional[45675:45672], addr_11418_7);

wire[31:0] addr_11419_7;

Selector_2 s11419_7(wires_2854_6[3], addr_2854_6, addr_positional[45679:45676], addr_11419_7);

wire[31:0] addr_11420_7;

Selector_2 s11420_7(wires_2855_6[0], addr_2855_6, addr_positional[45683:45680], addr_11420_7);

wire[31:0] addr_11421_7;

Selector_2 s11421_7(wires_2855_6[1], addr_2855_6, addr_positional[45687:45684], addr_11421_7);

wire[31:0] addr_11422_7;

Selector_2 s11422_7(wires_2855_6[2], addr_2855_6, addr_positional[45691:45688], addr_11422_7);

wire[31:0] addr_11423_7;

Selector_2 s11423_7(wires_2855_6[3], addr_2855_6, addr_positional[45695:45692], addr_11423_7);

wire[31:0] addr_11424_7;

Selector_2 s11424_7(wires_2856_6[0], addr_2856_6, addr_positional[45699:45696], addr_11424_7);

wire[31:0] addr_11425_7;

Selector_2 s11425_7(wires_2856_6[1], addr_2856_6, addr_positional[45703:45700], addr_11425_7);

wire[31:0] addr_11426_7;

Selector_2 s11426_7(wires_2856_6[2], addr_2856_6, addr_positional[45707:45704], addr_11426_7);

wire[31:0] addr_11427_7;

Selector_2 s11427_7(wires_2856_6[3], addr_2856_6, addr_positional[45711:45708], addr_11427_7);

wire[31:0] addr_11428_7;

Selector_2 s11428_7(wires_2857_6[0], addr_2857_6, addr_positional[45715:45712], addr_11428_7);

wire[31:0] addr_11429_7;

Selector_2 s11429_7(wires_2857_6[1], addr_2857_6, addr_positional[45719:45716], addr_11429_7);

wire[31:0] addr_11430_7;

Selector_2 s11430_7(wires_2857_6[2], addr_2857_6, addr_positional[45723:45720], addr_11430_7);

wire[31:0] addr_11431_7;

Selector_2 s11431_7(wires_2857_6[3], addr_2857_6, addr_positional[45727:45724], addr_11431_7);

wire[31:0] addr_11432_7;

Selector_2 s11432_7(wires_2858_6[0], addr_2858_6, addr_positional[45731:45728], addr_11432_7);

wire[31:0] addr_11433_7;

Selector_2 s11433_7(wires_2858_6[1], addr_2858_6, addr_positional[45735:45732], addr_11433_7);

wire[31:0] addr_11434_7;

Selector_2 s11434_7(wires_2858_6[2], addr_2858_6, addr_positional[45739:45736], addr_11434_7);

wire[31:0] addr_11435_7;

Selector_2 s11435_7(wires_2858_6[3], addr_2858_6, addr_positional[45743:45740], addr_11435_7);

wire[31:0] addr_11436_7;

Selector_2 s11436_7(wires_2859_6[0], addr_2859_6, addr_positional[45747:45744], addr_11436_7);

wire[31:0] addr_11437_7;

Selector_2 s11437_7(wires_2859_6[1], addr_2859_6, addr_positional[45751:45748], addr_11437_7);

wire[31:0] addr_11438_7;

Selector_2 s11438_7(wires_2859_6[2], addr_2859_6, addr_positional[45755:45752], addr_11438_7);

wire[31:0] addr_11439_7;

Selector_2 s11439_7(wires_2859_6[3], addr_2859_6, addr_positional[45759:45756], addr_11439_7);

wire[31:0] addr_11440_7;

Selector_2 s11440_7(wires_2860_6[0], addr_2860_6, addr_positional[45763:45760], addr_11440_7);

wire[31:0] addr_11441_7;

Selector_2 s11441_7(wires_2860_6[1], addr_2860_6, addr_positional[45767:45764], addr_11441_7);

wire[31:0] addr_11442_7;

Selector_2 s11442_7(wires_2860_6[2], addr_2860_6, addr_positional[45771:45768], addr_11442_7);

wire[31:0] addr_11443_7;

Selector_2 s11443_7(wires_2860_6[3], addr_2860_6, addr_positional[45775:45772], addr_11443_7);

wire[31:0] addr_11444_7;

Selector_2 s11444_7(wires_2861_6[0], addr_2861_6, addr_positional[45779:45776], addr_11444_7);

wire[31:0] addr_11445_7;

Selector_2 s11445_7(wires_2861_6[1], addr_2861_6, addr_positional[45783:45780], addr_11445_7);

wire[31:0] addr_11446_7;

Selector_2 s11446_7(wires_2861_6[2], addr_2861_6, addr_positional[45787:45784], addr_11446_7);

wire[31:0] addr_11447_7;

Selector_2 s11447_7(wires_2861_6[3], addr_2861_6, addr_positional[45791:45788], addr_11447_7);

wire[31:0] addr_11448_7;

Selector_2 s11448_7(wires_2862_6[0], addr_2862_6, addr_positional[45795:45792], addr_11448_7);

wire[31:0] addr_11449_7;

Selector_2 s11449_7(wires_2862_6[1], addr_2862_6, addr_positional[45799:45796], addr_11449_7);

wire[31:0] addr_11450_7;

Selector_2 s11450_7(wires_2862_6[2], addr_2862_6, addr_positional[45803:45800], addr_11450_7);

wire[31:0] addr_11451_7;

Selector_2 s11451_7(wires_2862_6[3], addr_2862_6, addr_positional[45807:45804], addr_11451_7);

wire[31:0] addr_11452_7;

Selector_2 s11452_7(wires_2863_6[0], addr_2863_6, addr_positional[45811:45808], addr_11452_7);

wire[31:0] addr_11453_7;

Selector_2 s11453_7(wires_2863_6[1], addr_2863_6, addr_positional[45815:45812], addr_11453_7);

wire[31:0] addr_11454_7;

Selector_2 s11454_7(wires_2863_6[2], addr_2863_6, addr_positional[45819:45816], addr_11454_7);

wire[31:0] addr_11455_7;

Selector_2 s11455_7(wires_2863_6[3], addr_2863_6, addr_positional[45823:45820], addr_11455_7);

wire[31:0] addr_11456_7;

Selector_2 s11456_7(wires_2864_6[0], addr_2864_6, addr_positional[45827:45824], addr_11456_7);

wire[31:0] addr_11457_7;

Selector_2 s11457_7(wires_2864_6[1], addr_2864_6, addr_positional[45831:45828], addr_11457_7);

wire[31:0] addr_11458_7;

Selector_2 s11458_7(wires_2864_6[2], addr_2864_6, addr_positional[45835:45832], addr_11458_7);

wire[31:0] addr_11459_7;

Selector_2 s11459_7(wires_2864_6[3], addr_2864_6, addr_positional[45839:45836], addr_11459_7);

wire[31:0] addr_11460_7;

Selector_2 s11460_7(wires_2865_6[0], addr_2865_6, addr_positional[45843:45840], addr_11460_7);

wire[31:0] addr_11461_7;

Selector_2 s11461_7(wires_2865_6[1], addr_2865_6, addr_positional[45847:45844], addr_11461_7);

wire[31:0] addr_11462_7;

Selector_2 s11462_7(wires_2865_6[2], addr_2865_6, addr_positional[45851:45848], addr_11462_7);

wire[31:0] addr_11463_7;

Selector_2 s11463_7(wires_2865_6[3], addr_2865_6, addr_positional[45855:45852], addr_11463_7);

wire[31:0] addr_11464_7;

Selector_2 s11464_7(wires_2866_6[0], addr_2866_6, addr_positional[45859:45856], addr_11464_7);

wire[31:0] addr_11465_7;

Selector_2 s11465_7(wires_2866_6[1], addr_2866_6, addr_positional[45863:45860], addr_11465_7);

wire[31:0] addr_11466_7;

Selector_2 s11466_7(wires_2866_6[2], addr_2866_6, addr_positional[45867:45864], addr_11466_7);

wire[31:0] addr_11467_7;

Selector_2 s11467_7(wires_2866_6[3], addr_2866_6, addr_positional[45871:45868], addr_11467_7);

wire[31:0] addr_11468_7;

Selector_2 s11468_7(wires_2867_6[0], addr_2867_6, addr_positional[45875:45872], addr_11468_7);

wire[31:0] addr_11469_7;

Selector_2 s11469_7(wires_2867_6[1], addr_2867_6, addr_positional[45879:45876], addr_11469_7);

wire[31:0] addr_11470_7;

Selector_2 s11470_7(wires_2867_6[2], addr_2867_6, addr_positional[45883:45880], addr_11470_7);

wire[31:0] addr_11471_7;

Selector_2 s11471_7(wires_2867_6[3], addr_2867_6, addr_positional[45887:45884], addr_11471_7);

wire[31:0] addr_11472_7;

Selector_2 s11472_7(wires_2868_6[0], addr_2868_6, addr_positional[45891:45888], addr_11472_7);

wire[31:0] addr_11473_7;

Selector_2 s11473_7(wires_2868_6[1], addr_2868_6, addr_positional[45895:45892], addr_11473_7);

wire[31:0] addr_11474_7;

Selector_2 s11474_7(wires_2868_6[2], addr_2868_6, addr_positional[45899:45896], addr_11474_7);

wire[31:0] addr_11475_7;

Selector_2 s11475_7(wires_2868_6[3], addr_2868_6, addr_positional[45903:45900], addr_11475_7);

wire[31:0] addr_11476_7;

Selector_2 s11476_7(wires_2869_6[0], addr_2869_6, addr_positional[45907:45904], addr_11476_7);

wire[31:0] addr_11477_7;

Selector_2 s11477_7(wires_2869_6[1], addr_2869_6, addr_positional[45911:45908], addr_11477_7);

wire[31:0] addr_11478_7;

Selector_2 s11478_7(wires_2869_6[2], addr_2869_6, addr_positional[45915:45912], addr_11478_7);

wire[31:0] addr_11479_7;

Selector_2 s11479_7(wires_2869_6[3], addr_2869_6, addr_positional[45919:45916], addr_11479_7);

wire[31:0] addr_11480_7;

Selector_2 s11480_7(wires_2870_6[0], addr_2870_6, addr_positional[45923:45920], addr_11480_7);

wire[31:0] addr_11481_7;

Selector_2 s11481_7(wires_2870_6[1], addr_2870_6, addr_positional[45927:45924], addr_11481_7);

wire[31:0] addr_11482_7;

Selector_2 s11482_7(wires_2870_6[2], addr_2870_6, addr_positional[45931:45928], addr_11482_7);

wire[31:0] addr_11483_7;

Selector_2 s11483_7(wires_2870_6[3], addr_2870_6, addr_positional[45935:45932], addr_11483_7);

wire[31:0] addr_11484_7;

Selector_2 s11484_7(wires_2871_6[0], addr_2871_6, addr_positional[45939:45936], addr_11484_7);

wire[31:0] addr_11485_7;

Selector_2 s11485_7(wires_2871_6[1], addr_2871_6, addr_positional[45943:45940], addr_11485_7);

wire[31:0] addr_11486_7;

Selector_2 s11486_7(wires_2871_6[2], addr_2871_6, addr_positional[45947:45944], addr_11486_7);

wire[31:0] addr_11487_7;

Selector_2 s11487_7(wires_2871_6[3], addr_2871_6, addr_positional[45951:45948], addr_11487_7);

wire[31:0] addr_11488_7;

Selector_2 s11488_7(wires_2872_6[0], addr_2872_6, addr_positional[45955:45952], addr_11488_7);

wire[31:0] addr_11489_7;

Selector_2 s11489_7(wires_2872_6[1], addr_2872_6, addr_positional[45959:45956], addr_11489_7);

wire[31:0] addr_11490_7;

Selector_2 s11490_7(wires_2872_6[2], addr_2872_6, addr_positional[45963:45960], addr_11490_7);

wire[31:0] addr_11491_7;

Selector_2 s11491_7(wires_2872_6[3], addr_2872_6, addr_positional[45967:45964], addr_11491_7);

wire[31:0] addr_11492_7;

Selector_2 s11492_7(wires_2873_6[0], addr_2873_6, addr_positional[45971:45968], addr_11492_7);

wire[31:0] addr_11493_7;

Selector_2 s11493_7(wires_2873_6[1], addr_2873_6, addr_positional[45975:45972], addr_11493_7);

wire[31:0] addr_11494_7;

Selector_2 s11494_7(wires_2873_6[2], addr_2873_6, addr_positional[45979:45976], addr_11494_7);

wire[31:0] addr_11495_7;

Selector_2 s11495_7(wires_2873_6[3], addr_2873_6, addr_positional[45983:45980], addr_11495_7);

wire[31:0] addr_11496_7;

Selector_2 s11496_7(wires_2874_6[0], addr_2874_6, addr_positional[45987:45984], addr_11496_7);

wire[31:0] addr_11497_7;

Selector_2 s11497_7(wires_2874_6[1], addr_2874_6, addr_positional[45991:45988], addr_11497_7);

wire[31:0] addr_11498_7;

Selector_2 s11498_7(wires_2874_6[2], addr_2874_6, addr_positional[45995:45992], addr_11498_7);

wire[31:0] addr_11499_7;

Selector_2 s11499_7(wires_2874_6[3], addr_2874_6, addr_positional[45999:45996], addr_11499_7);

wire[31:0] addr_11500_7;

Selector_2 s11500_7(wires_2875_6[0], addr_2875_6, addr_positional[46003:46000], addr_11500_7);

wire[31:0] addr_11501_7;

Selector_2 s11501_7(wires_2875_6[1], addr_2875_6, addr_positional[46007:46004], addr_11501_7);

wire[31:0] addr_11502_7;

Selector_2 s11502_7(wires_2875_6[2], addr_2875_6, addr_positional[46011:46008], addr_11502_7);

wire[31:0] addr_11503_7;

Selector_2 s11503_7(wires_2875_6[3], addr_2875_6, addr_positional[46015:46012], addr_11503_7);

wire[31:0] addr_11504_7;

Selector_2 s11504_7(wires_2876_6[0], addr_2876_6, addr_positional[46019:46016], addr_11504_7);

wire[31:0] addr_11505_7;

Selector_2 s11505_7(wires_2876_6[1], addr_2876_6, addr_positional[46023:46020], addr_11505_7);

wire[31:0] addr_11506_7;

Selector_2 s11506_7(wires_2876_6[2], addr_2876_6, addr_positional[46027:46024], addr_11506_7);

wire[31:0] addr_11507_7;

Selector_2 s11507_7(wires_2876_6[3], addr_2876_6, addr_positional[46031:46028], addr_11507_7);

wire[31:0] addr_11508_7;

Selector_2 s11508_7(wires_2877_6[0], addr_2877_6, addr_positional[46035:46032], addr_11508_7);

wire[31:0] addr_11509_7;

Selector_2 s11509_7(wires_2877_6[1], addr_2877_6, addr_positional[46039:46036], addr_11509_7);

wire[31:0] addr_11510_7;

Selector_2 s11510_7(wires_2877_6[2], addr_2877_6, addr_positional[46043:46040], addr_11510_7);

wire[31:0] addr_11511_7;

Selector_2 s11511_7(wires_2877_6[3], addr_2877_6, addr_positional[46047:46044], addr_11511_7);

wire[31:0] addr_11512_7;

Selector_2 s11512_7(wires_2878_6[0], addr_2878_6, addr_positional[46051:46048], addr_11512_7);

wire[31:0] addr_11513_7;

Selector_2 s11513_7(wires_2878_6[1], addr_2878_6, addr_positional[46055:46052], addr_11513_7);

wire[31:0] addr_11514_7;

Selector_2 s11514_7(wires_2878_6[2], addr_2878_6, addr_positional[46059:46056], addr_11514_7);

wire[31:0] addr_11515_7;

Selector_2 s11515_7(wires_2878_6[3], addr_2878_6, addr_positional[46063:46060], addr_11515_7);

wire[31:0] addr_11516_7;

Selector_2 s11516_7(wires_2879_6[0], addr_2879_6, addr_positional[46067:46064], addr_11516_7);

wire[31:0] addr_11517_7;

Selector_2 s11517_7(wires_2879_6[1], addr_2879_6, addr_positional[46071:46068], addr_11517_7);

wire[31:0] addr_11518_7;

Selector_2 s11518_7(wires_2879_6[2], addr_2879_6, addr_positional[46075:46072], addr_11518_7);

wire[31:0] addr_11519_7;

Selector_2 s11519_7(wires_2879_6[3], addr_2879_6, addr_positional[46079:46076], addr_11519_7);

wire[31:0] addr_11520_7;

Selector_2 s11520_7(wires_2880_6[0], addr_2880_6, addr_positional[46083:46080], addr_11520_7);

wire[31:0] addr_11521_7;

Selector_2 s11521_7(wires_2880_6[1], addr_2880_6, addr_positional[46087:46084], addr_11521_7);

wire[31:0] addr_11522_7;

Selector_2 s11522_7(wires_2880_6[2], addr_2880_6, addr_positional[46091:46088], addr_11522_7);

wire[31:0] addr_11523_7;

Selector_2 s11523_7(wires_2880_6[3], addr_2880_6, addr_positional[46095:46092], addr_11523_7);

wire[31:0] addr_11524_7;

Selector_2 s11524_7(wires_2881_6[0], addr_2881_6, addr_positional[46099:46096], addr_11524_7);

wire[31:0] addr_11525_7;

Selector_2 s11525_7(wires_2881_6[1], addr_2881_6, addr_positional[46103:46100], addr_11525_7);

wire[31:0] addr_11526_7;

Selector_2 s11526_7(wires_2881_6[2], addr_2881_6, addr_positional[46107:46104], addr_11526_7);

wire[31:0] addr_11527_7;

Selector_2 s11527_7(wires_2881_6[3], addr_2881_6, addr_positional[46111:46108], addr_11527_7);

wire[31:0] addr_11528_7;

Selector_2 s11528_7(wires_2882_6[0], addr_2882_6, addr_positional[46115:46112], addr_11528_7);

wire[31:0] addr_11529_7;

Selector_2 s11529_7(wires_2882_6[1], addr_2882_6, addr_positional[46119:46116], addr_11529_7);

wire[31:0] addr_11530_7;

Selector_2 s11530_7(wires_2882_6[2], addr_2882_6, addr_positional[46123:46120], addr_11530_7);

wire[31:0] addr_11531_7;

Selector_2 s11531_7(wires_2882_6[3], addr_2882_6, addr_positional[46127:46124], addr_11531_7);

wire[31:0] addr_11532_7;

Selector_2 s11532_7(wires_2883_6[0], addr_2883_6, addr_positional[46131:46128], addr_11532_7);

wire[31:0] addr_11533_7;

Selector_2 s11533_7(wires_2883_6[1], addr_2883_6, addr_positional[46135:46132], addr_11533_7);

wire[31:0] addr_11534_7;

Selector_2 s11534_7(wires_2883_6[2], addr_2883_6, addr_positional[46139:46136], addr_11534_7);

wire[31:0] addr_11535_7;

Selector_2 s11535_7(wires_2883_6[3], addr_2883_6, addr_positional[46143:46140], addr_11535_7);

wire[31:0] addr_11536_7;

Selector_2 s11536_7(wires_2884_6[0], addr_2884_6, addr_positional[46147:46144], addr_11536_7);

wire[31:0] addr_11537_7;

Selector_2 s11537_7(wires_2884_6[1], addr_2884_6, addr_positional[46151:46148], addr_11537_7);

wire[31:0] addr_11538_7;

Selector_2 s11538_7(wires_2884_6[2], addr_2884_6, addr_positional[46155:46152], addr_11538_7);

wire[31:0] addr_11539_7;

Selector_2 s11539_7(wires_2884_6[3], addr_2884_6, addr_positional[46159:46156], addr_11539_7);

wire[31:0] addr_11540_7;

Selector_2 s11540_7(wires_2885_6[0], addr_2885_6, addr_positional[46163:46160], addr_11540_7);

wire[31:0] addr_11541_7;

Selector_2 s11541_7(wires_2885_6[1], addr_2885_6, addr_positional[46167:46164], addr_11541_7);

wire[31:0] addr_11542_7;

Selector_2 s11542_7(wires_2885_6[2], addr_2885_6, addr_positional[46171:46168], addr_11542_7);

wire[31:0] addr_11543_7;

Selector_2 s11543_7(wires_2885_6[3], addr_2885_6, addr_positional[46175:46172], addr_11543_7);

wire[31:0] addr_11544_7;

Selector_2 s11544_7(wires_2886_6[0], addr_2886_6, addr_positional[46179:46176], addr_11544_7);

wire[31:0] addr_11545_7;

Selector_2 s11545_7(wires_2886_6[1], addr_2886_6, addr_positional[46183:46180], addr_11545_7);

wire[31:0] addr_11546_7;

Selector_2 s11546_7(wires_2886_6[2], addr_2886_6, addr_positional[46187:46184], addr_11546_7);

wire[31:0] addr_11547_7;

Selector_2 s11547_7(wires_2886_6[3], addr_2886_6, addr_positional[46191:46188], addr_11547_7);

wire[31:0] addr_11548_7;

Selector_2 s11548_7(wires_2887_6[0], addr_2887_6, addr_positional[46195:46192], addr_11548_7);

wire[31:0] addr_11549_7;

Selector_2 s11549_7(wires_2887_6[1], addr_2887_6, addr_positional[46199:46196], addr_11549_7);

wire[31:0] addr_11550_7;

Selector_2 s11550_7(wires_2887_6[2], addr_2887_6, addr_positional[46203:46200], addr_11550_7);

wire[31:0] addr_11551_7;

Selector_2 s11551_7(wires_2887_6[3], addr_2887_6, addr_positional[46207:46204], addr_11551_7);

wire[31:0] addr_11552_7;

Selector_2 s11552_7(wires_2888_6[0], addr_2888_6, addr_positional[46211:46208], addr_11552_7);

wire[31:0] addr_11553_7;

Selector_2 s11553_7(wires_2888_6[1], addr_2888_6, addr_positional[46215:46212], addr_11553_7);

wire[31:0] addr_11554_7;

Selector_2 s11554_7(wires_2888_6[2], addr_2888_6, addr_positional[46219:46216], addr_11554_7);

wire[31:0] addr_11555_7;

Selector_2 s11555_7(wires_2888_6[3], addr_2888_6, addr_positional[46223:46220], addr_11555_7);

wire[31:0] addr_11556_7;

Selector_2 s11556_7(wires_2889_6[0], addr_2889_6, addr_positional[46227:46224], addr_11556_7);

wire[31:0] addr_11557_7;

Selector_2 s11557_7(wires_2889_6[1], addr_2889_6, addr_positional[46231:46228], addr_11557_7);

wire[31:0] addr_11558_7;

Selector_2 s11558_7(wires_2889_6[2], addr_2889_6, addr_positional[46235:46232], addr_11558_7);

wire[31:0] addr_11559_7;

Selector_2 s11559_7(wires_2889_6[3], addr_2889_6, addr_positional[46239:46236], addr_11559_7);

wire[31:0] addr_11560_7;

Selector_2 s11560_7(wires_2890_6[0], addr_2890_6, addr_positional[46243:46240], addr_11560_7);

wire[31:0] addr_11561_7;

Selector_2 s11561_7(wires_2890_6[1], addr_2890_6, addr_positional[46247:46244], addr_11561_7);

wire[31:0] addr_11562_7;

Selector_2 s11562_7(wires_2890_6[2], addr_2890_6, addr_positional[46251:46248], addr_11562_7);

wire[31:0] addr_11563_7;

Selector_2 s11563_7(wires_2890_6[3], addr_2890_6, addr_positional[46255:46252], addr_11563_7);

wire[31:0] addr_11564_7;

Selector_2 s11564_7(wires_2891_6[0], addr_2891_6, addr_positional[46259:46256], addr_11564_7);

wire[31:0] addr_11565_7;

Selector_2 s11565_7(wires_2891_6[1], addr_2891_6, addr_positional[46263:46260], addr_11565_7);

wire[31:0] addr_11566_7;

Selector_2 s11566_7(wires_2891_6[2], addr_2891_6, addr_positional[46267:46264], addr_11566_7);

wire[31:0] addr_11567_7;

Selector_2 s11567_7(wires_2891_6[3], addr_2891_6, addr_positional[46271:46268], addr_11567_7);

wire[31:0] addr_11568_7;

Selector_2 s11568_7(wires_2892_6[0], addr_2892_6, addr_positional[46275:46272], addr_11568_7);

wire[31:0] addr_11569_7;

Selector_2 s11569_7(wires_2892_6[1], addr_2892_6, addr_positional[46279:46276], addr_11569_7);

wire[31:0] addr_11570_7;

Selector_2 s11570_7(wires_2892_6[2], addr_2892_6, addr_positional[46283:46280], addr_11570_7);

wire[31:0] addr_11571_7;

Selector_2 s11571_7(wires_2892_6[3], addr_2892_6, addr_positional[46287:46284], addr_11571_7);

wire[31:0] addr_11572_7;

Selector_2 s11572_7(wires_2893_6[0], addr_2893_6, addr_positional[46291:46288], addr_11572_7);

wire[31:0] addr_11573_7;

Selector_2 s11573_7(wires_2893_6[1], addr_2893_6, addr_positional[46295:46292], addr_11573_7);

wire[31:0] addr_11574_7;

Selector_2 s11574_7(wires_2893_6[2], addr_2893_6, addr_positional[46299:46296], addr_11574_7);

wire[31:0] addr_11575_7;

Selector_2 s11575_7(wires_2893_6[3], addr_2893_6, addr_positional[46303:46300], addr_11575_7);

wire[31:0] addr_11576_7;

Selector_2 s11576_7(wires_2894_6[0], addr_2894_6, addr_positional[46307:46304], addr_11576_7);

wire[31:0] addr_11577_7;

Selector_2 s11577_7(wires_2894_6[1], addr_2894_6, addr_positional[46311:46308], addr_11577_7);

wire[31:0] addr_11578_7;

Selector_2 s11578_7(wires_2894_6[2], addr_2894_6, addr_positional[46315:46312], addr_11578_7);

wire[31:0] addr_11579_7;

Selector_2 s11579_7(wires_2894_6[3], addr_2894_6, addr_positional[46319:46316], addr_11579_7);

wire[31:0] addr_11580_7;

Selector_2 s11580_7(wires_2895_6[0], addr_2895_6, addr_positional[46323:46320], addr_11580_7);

wire[31:0] addr_11581_7;

Selector_2 s11581_7(wires_2895_6[1], addr_2895_6, addr_positional[46327:46324], addr_11581_7);

wire[31:0] addr_11582_7;

Selector_2 s11582_7(wires_2895_6[2], addr_2895_6, addr_positional[46331:46328], addr_11582_7);

wire[31:0] addr_11583_7;

Selector_2 s11583_7(wires_2895_6[3], addr_2895_6, addr_positional[46335:46332], addr_11583_7);

wire[31:0] addr_11584_7;

Selector_2 s11584_7(wires_2896_6[0], addr_2896_6, addr_positional[46339:46336], addr_11584_7);

wire[31:0] addr_11585_7;

Selector_2 s11585_7(wires_2896_6[1], addr_2896_6, addr_positional[46343:46340], addr_11585_7);

wire[31:0] addr_11586_7;

Selector_2 s11586_7(wires_2896_6[2], addr_2896_6, addr_positional[46347:46344], addr_11586_7);

wire[31:0] addr_11587_7;

Selector_2 s11587_7(wires_2896_6[3], addr_2896_6, addr_positional[46351:46348], addr_11587_7);

wire[31:0] addr_11588_7;

Selector_2 s11588_7(wires_2897_6[0], addr_2897_6, addr_positional[46355:46352], addr_11588_7);

wire[31:0] addr_11589_7;

Selector_2 s11589_7(wires_2897_6[1], addr_2897_6, addr_positional[46359:46356], addr_11589_7);

wire[31:0] addr_11590_7;

Selector_2 s11590_7(wires_2897_6[2], addr_2897_6, addr_positional[46363:46360], addr_11590_7);

wire[31:0] addr_11591_7;

Selector_2 s11591_7(wires_2897_6[3], addr_2897_6, addr_positional[46367:46364], addr_11591_7);

wire[31:0] addr_11592_7;

Selector_2 s11592_7(wires_2898_6[0], addr_2898_6, addr_positional[46371:46368], addr_11592_7);

wire[31:0] addr_11593_7;

Selector_2 s11593_7(wires_2898_6[1], addr_2898_6, addr_positional[46375:46372], addr_11593_7);

wire[31:0] addr_11594_7;

Selector_2 s11594_7(wires_2898_6[2], addr_2898_6, addr_positional[46379:46376], addr_11594_7);

wire[31:0] addr_11595_7;

Selector_2 s11595_7(wires_2898_6[3], addr_2898_6, addr_positional[46383:46380], addr_11595_7);

wire[31:0] addr_11596_7;

Selector_2 s11596_7(wires_2899_6[0], addr_2899_6, addr_positional[46387:46384], addr_11596_7);

wire[31:0] addr_11597_7;

Selector_2 s11597_7(wires_2899_6[1], addr_2899_6, addr_positional[46391:46388], addr_11597_7);

wire[31:0] addr_11598_7;

Selector_2 s11598_7(wires_2899_6[2], addr_2899_6, addr_positional[46395:46392], addr_11598_7);

wire[31:0] addr_11599_7;

Selector_2 s11599_7(wires_2899_6[3], addr_2899_6, addr_positional[46399:46396], addr_11599_7);

wire[31:0] addr_11600_7;

Selector_2 s11600_7(wires_2900_6[0], addr_2900_6, addr_positional[46403:46400], addr_11600_7);

wire[31:0] addr_11601_7;

Selector_2 s11601_7(wires_2900_6[1], addr_2900_6, addr_positional[46407:46404], addr_11601_7);

wire[31:0] addr_11602_7;

Selector_2 s11602_7(wires_2900_6[2], addr_2900_6, addr_positional[46411:46408], addr_11602_7);

wire[31:0] addr_11603_7;

Selector_2 s11603_7(wires_2900_6[3], addr_2900_6, addr_positional[46415:46412], addr_11603_7);

wire[31:0] addr_11604_7;

Selector_2 s11604_7(wires_2901_6[0], addr_2901_6, addr_positional[46419:46416], addr_11604_7);

wire[31:0] addr_11605_7;

Selector_2 s11605_7(wires_2901_6[1], addr_2901_6, addr_positional[46423:46420], addr_11605_7);

wire[31:0] addr_11606_7;

Selector_2 s11606_7(wires_2901_6[2], addr_2901_6, addr_positional[46427:46424], addr_11606_7);

wire[31:0] addr_11607_7;

Selector_2 s11607_7(wires_2901_6[3], addr_2901_6, addr_positional[46431:46428], addr_11607_7);

wire[31:0] addr_11608_7;

Selector_2 s11608_7(wires_2902_6[0], addr_2902_6, addr_positional[46435:46432], addr_11608_7);

wire[31:0] addr_11609_7;

Selector_2 s11609_7(wires_2902_6[1], addr_2902_6, addr_positional[46439:46436], addr_11609_7);

wire[31:0] addr_11610_7;

Selector_2 s11610_7(wires_2902_6[2], addr_2902_6, addr_positional[46443:46440], addr_11610_7);

wire[31:0] addr_11611_7;

Selector_2 s11611_7(wires_2902_6[3], addr_2902_6, addr_positional[46447:46444], addr_11611_7);

wire[31:0] addr_11612_7;

Selector_2 s11612_7(wires_2903_6[0], addr_2903_6, addr_positional[46451:46448], addr_11612_7);

wire[31:0] addr_11613_7;

Selector_2 s11613_7(wires_2903_6[1], addr_2903_6, addr_positional[46455:46452], addr_11613_7);

wire[31:0] addr_11614_7;

Selector_2 s11614_7(wires_2903_6[2], addr_2903_6, addr_positional[46459:46456], addr_11614_7);

wire[31:0] addr_11615_7;

Selector_2 s11615_7(wires_2903_6[3], addr_2903_6, addr_positional[46463:46460], addr_11615_7);

wire[31:0] addr_11616_7;

Selector_2 s11616_7(wires_2904_6[0], addr_2904_6, addr_positional[46467:46464], addr_11616_7);

wire[31:0] addr_11617_7;

Selector_2 s11617_7(wires_2904_6[1], addr_2904_6, addr_positional[46471:46468], addr_11617_7);

wire[31:0] addr_11618_7;

Selector_2 s11618_7(wires_2904_6[2], addr_2904_6, addr_positional[46475:46472], addr_11618_7);

wire[31:0] addr_11619_7;

Selector_2 s11619_7(wires_2904_6[3], addr_2904_6, addr_positional[46479:46476], addr_11619_7);

wire[31:0] addr_11620_7;

Selector_2 s11620_7(wires_2905_6[0], addr_2905_6, addr_positional[46483:46480], addr_11620_7);

wire[31:0] addr_11621_7;

Selector_2 s11621_7(wires_2905_6[1], addr_2905_6, addr_positional[46487:46484], addr_11621_7);

wire[31:0] addr_11622_7;

Selector_2 s11622_7(wires_2905_6[2], addr_2905_6, addr_positional[46491:46488], addr_11622_7);

wire[31:0] addr_11623_7;

Selector_2 s11623_7(wires_2905_6[3], addr_2905_6, addr_positional[46495:46492], addr_11623_7);

wire[31:0] addr_11624_7;

Selector_2 s11624_7(wires_2906_6[0], addr_2906_6, addr_positional[46499:46496], addr_11624_7);

wire[31:0] addr_11625_7;

Selector_2 s11625_7(wires_2906_6[1], addr_2906_6, addr_positional[46503:46500], addr_11625_7);

wire[31:0] addr_11626_7;

Selector_2 s11626_7(wires_2906_6[2], addr_2906_6, addr_positional[46507:46504], addr_11626_7);

wire[31:0] addr_11627_7;

Selector_2 s11627_7(wires_2906_6[3], addr_2906_6, addr_positional[46511:46508], addr_11627_7);

wire[31:0] addr_11628_7;

Selector_2 s11628_7(wires_2907_6[0], addr_2907_6, addr_positional[46515:46512], addr_11628_7);

wire[31:0] addr_11629_7;

Selector_2 s11629_7(wires_2907_6[1], addr_2907_6, addr_positional[46519:46516], addr_11629_7);

wire[31:0] addr_11630_7;

Selector_2 s11630_7(wires_2907_6[2], addr_2907_6, addr_positional[46523:46520], addr_11630_7);

wire[31:0] addr_11631_7;

Selector_2 s11631_7(wires_2907_6[3], addr_2907_6, addr_positional[46527:46524], addr_11631_7);

wire[31:0] addr_11632_7;

Selector_2 s11632_7(wires_2908_6[0], addr_2908_6, addr_positional[46531:46528], addr_11632_7);

wire[31:0] addr_11633_7;

Selector_2 s11633_7(wires_2908_6[1], addr_2908_6, addr_positional[46535:46532], addr_11633_7);

wire[31:0] addr_11634_7;

Selector_2 s11634_7(wires_2908_6[2], addr_2908_6, addr_positional[46539:46536], addr_11634_7);

wire[31:0] addr_11635_7;

Selector_2 s11635_7(wires_2908_6[3], addr_2908_6, addr_positional[46543:46540], addr_11635_7);

wire[31:0] addr_11636_7;

Selector_2 s11636_7(wires_2909_6[0], addr_2909_6, addr_positional[46547:46544], addr_11636_7);

wire[31:0] addr_11637_7;

Selector_2 s11637_7(wires_2909_6[1], addr_2909_6, addr_positional[46551:46548], addr_11637_7);

wire[31:0] addr_11638_7;

Selector_2 s11638_7(wires_2909_6[2], addr_2909_6, addr_positional[46555:46552], addr_11638_7);

wire[31:0] addr_11639_7;

Selector_2 s11639_7(wires_2909_6[3], addr_2909_6, addr_positional[46559:46556], addr_11639_7);

wire[31:0] addr_11640_7;

Selector_2 s11640_7(wires_2910_6[0], addr_2910_6, addr_positional[46563:46560], addr_11640_7);

wire[31:0] addr_11641_7;

Selector_2 s11641_7(wires_2910_6[1], addr_2910_6, addr_positional[46567:46564], addr_11641_7);

wire[31:0] addr_11642_7;

Selector_2 s11642_7(wires_2910_6[2], addr_2910_6, addr_positional[46571:46568], addr_11642_7);

wire[31:0] addr_11643_7;

Selector_2 s11643_7(wires_2910_6[3], addr_2910_6, addr_positional[46575:46572], addr_11643_7);

wire[31:0] addr_11644_7;

Selector_2 s11644_7(wires_2911_6[0], addr_2911_6, addr_positional[46579:46576], addr_11644_7);

wire[31:0] addr_11645_7;

Selector_2 s11645_7(wires_2911_6[1], addr_2911_6, addr_positional[46583:46580], addr_11645_7);

wire[31:0] addr_11646_7;

Selector_2 s11646_7(wires_2911_6[2], addr_2911_6, addr_positional[46587:46584], addr_11646_7);

wire[31:0] addr_11647_7;

Selector_2 s11647_7(wires_2911_6[3], addr_2911_6, addr_positional[46591:46588], addr_11647_7);

wire[31:0] addr_11648_7;

Selector_2 s11648_7(wires_2912_6[0], addr_2912_6, addr_positional[46595:46592], addr_11648_7);

wire[31:0] addr_11649_7;

Selector_2 s11649_7(wires_2912_6[1], addr_2912_6, addr_positional[46599:46596], addr_11649_7);

wire[31:0] addr_11650_7;

Selector_2 s11650_7(wires_2912_6[2], addr_2912_6, addr_positional[46603:46600], addr_11650_7);

wire[31:0] addr_11651_7;

Selector_2 s11651_7(wires_2912_6[3], addr_2912_6, addr_positional[46607:46604], addr_11651_7);

wire[31:0] addr_11652_7;

Selector_2 s11652_7(wires_2913_6[0], addr_2913_6, addr_positional[46611:46608], addr_11652_7);

wire[31:0] addr_11653_7;

Selector_2 s11653_7(wires_2913_6[1], addr_2913_6, addr_positional[46615:46612], addr_11653_7);

wire[31:0] addr_11654_7;

Selector_2 s11654_7(wires_2913_6[2], addr_2913_6, addr_positional[46619:46616], addr_11654_7);

wire[31:0] addr_11655_7;

Selector_2 s11655_7(wires_2913_6[3], addr_2913_6, addr_positional[46623:46620], addr_11655_7);

wire[31:0] addr_11656_7;

Selector_2 s11656_7(wires_2914_6[0], addr_2914_6, addr_positional[46627:46624], addr_11656_7);

wire[31:0] addr_11657_7;

Selector_2 s11657_7(wires_2914_6[1], addr_2914_6, addr_positional[46631:46628], addr_11657_7);

wire[31:0] addr_11658_7;

Selector_2 s11658_7(wires_2914_6[2], addr_2914_6, addr_positional[46635:46632], addr_11658_7);

wire[31:0] addr_11659_7;

Selector_2 s11659_7(wires_2914_6[3], addr_2914_6, addr_positional[46639:46636], addr_11659_7);

wire[31:0] addr_11660_7;

Selector_2 s11660_7(wires_2915_6[0], addr_2915_6, addr_positional[46643:46640], addr_11660_7);

wire[31:0] addr_11661_7;

Selector_2 s11661_7(wires_2915_6[1], addr_2915_6, addr_positional[46647:46644], addr_11661_7);

wire[31:0] addr_11662_7;

Selector_2 s11662_7(wires_2915_6[2], addr_2915_6, addr_positional[46651:46648], addr_11662_7);

wire[31:0] addr_11663_7;

Selector_2 s11663_7(wires_2915_6[3], addr_2915_6, addr_positional[46655:46652], addr_11663_7);

wire[31:0] addr_11664_7;

Selector_2 s11664_7(wires_2916_6[0], addr_2916_6, addr_positional[46659:46656], addr_11664_7);

wire[31:0] addr_11665_7;

Selector_2 s11665_7(wires_2916_6[1], addr_2916_6, addr_positional[46663:46660], addr_11665_7);

wire[31:0] addr_11666_7;

Selector_2 s11666_7(wires_2916_6[2], addr_2916_6, addr_positional[46667:46664], addr_11666_7);

wire[31:0] addr_11667_7;

Selector_2 s11667_7(wires_2916_6[3], addr_2916_6, addr_positional[46671:46668], addr_11667_7);

wire[31:0] addr_11668_7;

Selector_2 s11668_7(wires_2917_6[0], addr_2917_6, addr_positional[46675:46672], addr_11668_7);

wire[31:0] addr_11669_7;

Selector_2 s11669_7(wires_2917_6[1], addr_2917_6, addr_positional[46679:46676], addr_11669_7);

wire[31:0] addr_11670_7;

Selector_2 s11670_7(wires_2917_6[2], addr_2917_6, addr_positional[46683:46680], addr_11670_7);

wire[31:0] addr_11671_7;

Selector_2 s11671_7(wires_2917_6[3], addr_2917_6, addr_positional[46687:46684], addr_11671_7);

wire[31:0] addr_11672_7;

Selector_2 s11672_7(wires_2918_6[0], addr_2918_6, addr_positional[46691:46688], addr_11672_7);

wire[31:0] addr_11673_7;

Selector_2 s11673_7(wires_2918_6[1], addr_2918_6, addr_positional[46695:46692], addr_11673_7);

wire[31:0] addr_11674_7;

Selector_2 s11674_7(wires_2918_6[2], addr_2918_6, addr_positional[46699:46696], addr_11674_7);

wire[31:0] addr_11675_7;

Selector_2 s11675_7(wires_2918_6[3], addr_2918_6, addr_positional[46703:46700], addr_11675_7);

wire[31:0] addr_11676_7;

Selector_2 s11676_7(wires_2919_6[0], addr_2919_6, addr_positional[46707:46704], addr_11676_7);

wire[31:0] addr_11677_7;

Selector_2 s11677_7(wires_2919_6[1], addr_2919_6, addr_positional[46711:46708], addr_11677_7);

wire[31:0] addr_11678_7;

Selector_2 s11678_7(wires_2919_6[2], addr_2919_6, addr_positional[46715:46712], addr_11678_7);

wire[31:0] addr_11679_7;

Selector_2 s11679_7(wires_2919_6[3], addr_2919_6, addr_positional[46719:46716], addr_11679_7);

wire[31:0] addr_11680_7;

Selector_2 s11680_7(wires_2920_6[0], addr_2920_6, addr_positional[46723:46720], addr_11680_7);

wire[31:0] addr_11681_7;

Selector_2 s11681_7(wires_2920_6[1], addr_2920_6, addr_positional[46727:46724], addr_11681_7);

wire[31:0] addr_11682_7;

Selector_2 s11682_7(wires_2920_6[2], addr_2920_6, addr_positional[46731:46728], addr_11682_7);

wire[31:0] addr_11683_7;

Selector_2 s11683_7(wires_2920_6[3], addr_2920_6, addr_positional[46735:46732], addr_11683_7);

wire[31:0] addr_11684_7;

Selector_2 s11684_7(wires_2921_6[0], addr_2921_6, addr_positional[46739:46736], addr_11684_7);

wire[31:0] addr_11685_7;

Selector_2 s11685_7(wires_2921_6[1], addr_2921_6, addr_positional[46743:46740], addr_11685_7);

wire[31:0] addr_11686_7;

Selector_2 s11686_7(wires_2921_6[2], addr_2921_6, addr_positional[46747:46744], addr_11686_7);

wire[31:0] addr_11687_7;

Selector_2 s11687_7(wires_2921_6[3], addr_2921_6, addr_positional[46751:46748], addr_11687_7);

wire[31:0] addr_11688_7;

Selector_2 s11688_7(wires_2922_6[0], addr_2922_6, addr_positional[46755:46752], addr_11688_7);

wire[31:0] addr_11689_7;

Selector_2 s11689_7(wires_2922_6[1], addr_2922_6, addr_positional[46759:46756], addr_11689_7);

wire[31:0] addr_11690_7;

Selector_2 s11690_7(wires_2922_6[2], addr_2922_6, addr_positional[46763:46760], addr_11690_7);

wire[31:0] addr_11691_7;

Selector_2 s11691_7(wires_2922_6[3], addr_2922_6, addr_positional[46767:46764], addr_11691_7);

wire[31:0] addr_11692_7;

Selector_2 s11692_7(wires_2923_6[0], addr_2923_6, addr_positional[46771:46768], addr_11692_7);

wire[31:0] addr_11693_7;

Selector_2 s11693_7(wires_2923_6[1], addr_2923_6, addr_positional[46775:46772], addr_11693_7);

wire[31:0] addr_11694_7;

Selector_2 s11694_7(wires_2923_6[2], addr_2923_6, addr_positional[46779:46776], addr_11694_7);

wire[31:0] addr_11695_7;

Selector_2 s11695_7(wires_2923_6[3], addr_2923_6, addr_positional[46783:46780], addr_11695_7);

wire[31:0] addr_11696_7;

Selector_2 s11696_7(wires_2924_6[0], addr_2924_6, addr_positional[46787:46784], addr_11696_7);

wire[31:0] addr_11697_7;

Selector_2 s11697_7(wires_2924_6[1], addr_2924_6, addr_positional[46791:46788], addr_11697_7);

wire[31:0] addr_11698_7;

Selector_2 s11698_7(wires_2924_6[2], addr_2924_6, addr_positional[46795:46792], addr_11698_7);

wire[31:0] addr_11699_7;

Selector_2 s11699_7(wires_2924_6[3], addr_2924_6, addr_positional[46799:46796], addr_11699_7);

wire[31:0] addr_11700_7;

Selector_2 s11700_7(wires_2925_6[0], addr_2925_6, addr_positional[46803:46800], addr_11700_7);

wire[31:0] addr_11701_7;

Selector_2 s11701_7(wires_2925_6[1], addr_2925_6, addr_positional[46807:46804], addr_11701_7);

wire[31:0] addr_11702_7;

Selector_2 s11702_7(wires_2925_6[2], addr_2925_6, addr_positional[46811:46808], addr_11702_7);

wire[31:0] addr_11703_7;

Selector_2 s11703_7(wires_2925_6[3], addr_2925_6, addr_positional[46815:46812], addr_11703_7);

wire[31:0] addr_11704_7;

Selector_2 s11704_7(wires_2926_6[0], addr_2926_6, addr_positional[46819:46816], addr_11704_7);

wire[31:0] addr_11705_7;

Selector_2 s11705_7(wires_2926_6[1], addr_2926_6, addr_positional[46823:46820], addr_11705_7);

wire[31:0] addr_11706_7;

Selector_2 s11706_7(wires_2926_6[2], addr_2926_6, addr_positional[46827:46824], addr_11706_7);

wire[31:0] addr_11707_7;

Selector_2 s11707_7(wires_2926_6[3], addr_2926_6, addr_positional[46831:46828], addr_11707_7);

wire[31:0] addr_11708_7;

Selector_2 s11708_7(wires_2927_6[0], addr_2927_6, addr_positional[46835:46832], addr_11708_7);

wire[31:0] addr_11709_7;

Selector_2 s11709_7(wires_2927_6[1], addr_2927_6, addr_positional[46839:46836], addr_11709_7);

wire[31:0] addr_11710_7;

Selector_2 s11710_7(wires_2927_6[2], addr_2927_6, addr_positional[46843:46840], addr_11710_7);

wire[31:0] addr_11711_7;

Selector_2 s11711_7(wires_2927_6[3], addr_2927_6, addr_positional[46847:46844], addr_11711_7);

wire[31:0] addr_11712_7;

Selector_2 s11712_7(wires_2928_6[0], addr_2928_6, addr_positional[46851:46848], addr_11712_7);

wire[31:0] addr_11713_7;

Selector_2 s11713_7(wires_2928_6[1], addr_2928_6, addr_positional[46855:46852], addr_11713_7);

wire[31:0] addr_11714_7;

Selector_2 s11714_7(wires_2928_6[2], addr_2928_6, addr_positional[46859:46856], addr_11714_7);

wire[31:0] addr_11715_7;

Selector_2 s11715_7(wires_2928_6[3], addr_2928_6, addr_positional[46863:46860], addr_11715_7);

wire[31:0] addr_11716_7;

Selector_2 s11716_7(wires_2929_6[0], addr_2929_6, addr_positional[46867:46864], addr_11716_7);

wire[31:0] addr_11717_7;

Selector_2 s11717_7(wires_2929_6[1], addr_2929_6, addr_positional[46871:46868], addr_11717_7);

wire[31:0] addr_11718_7;

Selector_2 s11718_7(wires_2929_6[2], addr_2929_6, addr_positional[46875:46872], addr_11718_7);

wire[31:0] addr_11719_7;

Selector_2 s11719_7(wires_2929_6[3], addr_2929_6, addr_positional[46879:46876], addr_11719_7);

wire[31:0] addr_11720_7;

Selector_2 s11720_7(wires_2930_6[0], addr_2930_6, addr_positional[46883:46880], addr_11720_7);

wire[31:0] addr_11721_7;

Selector_2 s11721_7(wires_2930_6[1], addr_2930_6, addr_positional[46887:46884], addr_11721_7);

wire[31:0] addr_11722_7;

Selector_2 s11722_7(wires_2930_6[2], addr_2930_6, addr_positional[46891:46888], addr_11722_7);

wire[31:0] addr_11723_7;

Selector_2 s11723_7(wires_2930_6[3], addr_2930_6, addr_positional[46895:46892], addr_11723_7);

wire[31:0] addr_11724_7;

Selector_2 s11724_7(wires_2931_6[0], addr_2931_6, addr_positional[46899:46896], addr_11724_7);

wire[31:0] addr_11725_7;

Selector_2 s11725_7(wires_2931_6[1], addr_2931_6, addr_positional[46903:46900], addr_11725_7);

wire[31:0] addr_11726_7;

Selector_2 s11726_7(wires_2931_6[2], addr_2931_6, addr_positional[46907:46904], addr_11726_7);

wire[31:0] addr_11727_7;

Selector_2 s11727_7(wires_2931_6[3], addr_2931_6, addr_positional[46911:46908], addr_11727_7);

wire[31:0] addr_11728_7;

Selector_2 s11728_7(wires_2932_6[0], addr_2932_6, addr_positional[46915:46912], addr_11728_7);

wire[31:0] addr_11729_7;

Selector_2 s11729_7(wires_2932_6[1], addr_2932_6, addr_positional[46919:46916], addr_11729_7);

wire[31:0] addr_11730_7;

Selector_2 s11730_7(wires_2932_6[2], addr_2932_6, addr_positional[46923:46920], addr_11730_7);

wire[31:0] addr_11731_7;

Selector_2 s11731_7(wires_2932_6[3], addr_2932_6, addr_positional[46927:46924], addr_11731_7);

wire[31:0] addr_11732_7;

Selector_2 s11732_7(wires_2933_6[0], addr_2933_6, addr_positional[46931:46928], addr_11732_7);

wire[31:0] addr_11733_7;

Selector_2 s11733_7(wires_2933_6[1], addr_2933_6, addr_positional[46935:46932], addr_11733_7);

wire[31:0] addr_11734_7;

Selector_2 s11734_7(wires_2933_6[2], addr_2933_6, addr_positional[46939:46936], addr_11734_7);

wire[31:0] addr_11735_7;

Selector_2 s11735_7(wires_2933_6[3], addr_2933_6, addr_positional[46943:46940], addr_11735_7);

wire[31:0] addr_11736_7;

Selector_2 s11736_7(wires_2934_6[0], addr_2934_6, addr_positional[46947:46944], addr_11736_7);

wire[31:0] addr_11737_7;

Selector_2 s11737_7(wires_2934_6[1], addr_2934_6, addr_positional[46951:46948], addr_11737_7);

wire[31:0] addr_11738_7;

Selector_2 s11738_7(wires_2934_6[2], addr_2934_6, addr_positional[46955:46952], addr_11738_7);

wire[31:0] addr_11739_7;

Selector_2 s11739_7(wires_2934_6[3], addr_2934_6, addr_positional[46959:46956], addr_11739_7);

wire[31:0] addr_11740_7;

Selector_2 s11740_7(wires_2935_6[0], addr_2935_6, addr_positional[46963:46960], addr_11740_7);

wire[31:0] addr_11741_7;

Selector_2 s11741_7(wires_2935_6[1], addr_2935_6, addr_positional[46967:46964], addr_11741_7);

wire[31:0] addr_11742_7;

Selector_2 s11742_7(wires_2935_6[2], addr_2935_6, addr_positional[46971:46968], addr_11742_7);

wire[31:0] addr_11743_7;

Selector_2 s11743_7(wires_2935_6[3], addr_2935_6, addr_positional[46975:46972], addr_11743_7);

wire[31:0] addr_11744_7;

Selector_2 s11744_7(wires_2936_6[0], addr_2936_6, addr_positional[46979:46976], addr_11744_7);

wire[31:0] addr_11745_7;

Selector_2 s11745_7(wires_2936_6[1], addr_2936_6, addr_positional[46983:46980], addr_11745_7);

wire[31:0] addr_11746_7;

Selector_2 s11746_7(wires_2936_6[2], addr_2936_6, addr_positional[46987:46984], addr_11746_7);

wire[31:0] addr_11747_7;

Selector_2 s11747_7(wires_2936_6[3], addr_2936_6, addr_positional[46991:46988], addr_11747_7);

wire[31:0] addr_11748_7;

Selector_2 s11748_7(wires_2937_6[0], addr_2937_6, addr_positional[46995:46992], addr_11748_7);

wire[31:0] addr_11749_7;

Selector_2 s11749_7(wires_2937_6[1], addr_2937_6, addr_positional[46999:46996], addr_11749_7);

wire[31:0] addr_11750_7;

Selector_2 s11750_7(wires_2937_6[2], addr_2937_6, addr_positional[47003:47000], addr_11750_7);

wire[31:0] addr_11751_7;

Selector_2 s11751_7(wires_2937_6[3], addr_2937_6, addr_positional[47007:47004], addr_11751_7);

wire[31:0] addr_11752_7;

Selector_2 s11752_7(wires_2938_6[0], addr_2938_6, addr_positional[47011:47008], addr_11752_7);

wire[31:0] addr_11753_7;

Selector_2 s11753_7(wires_2938_6[1], addr_2938_6, addr_positional[47015:47012], addr_11753_7);

wire[31:0] addr_11754_7;

Selector_2 s11754_7(wires_2938_6[2], addr_2938_6, addr_positional[47019:47016], addr_11754_7);

wire[31:0] addr_11755_7;

Selector_2 s11755_7(wires_2938_6[3], addr_2938_6, addr_positional[47023:47020], addr_11755_7);

wire[31:0] addr_11756_7;

Selector_2 s11756_7(wires_2939_6[0], addr_2939_6, addr_positional[47027:47024], addr_11756_7);

wire[31:0] addr_11757_7;

Selector_2 s11757_7(wires_2939_6[1], addr_2939_6, addr_positional[47031:47028], addr_11757_7);

wire[31:0] addr_11758_7;

Selector_2 s11758_7(wires_2939_6[2], addr_2939_6, addr_positional[47035:47032], addr_11758_7);

wire[31:0] addr_11759_7;

Selector_2 s11759_7(wires_2939_6[3], addr_2939_6, addr_positional[47039:47036], addr_11759_7);

wire[31:0] addr_11760_7;

Selector_2 s11760_7(wires_2940_6[0], addr_2940_6, addr_positional[47043:47040], addr_11760_7);

wire[31:0] addr_11761_7;

Selector_2 s11761_7(wires_2940_6[1], addr_2940_6, addr_positional[47047:47044], addr_11761_7);

wire[31:0] addr_11762_7;

Selector_2 s11762_7(wires_2940_6[2], addr_2940_6, addr_positional[47051:47048], addr_11762_7);

wire[31:0] addr_11763_7;

Selector_2 s11763_7(wires_2940_6[3], addr_2940_6, addr_positional[47055:47052], addr_11763_7);

wire[31:0] addr_11764_7;

Selector_2 s11764_7(wires_2941_6[0], addr_2941_6, addr_positional[47059:47056], addr_11764_7);

wire[31:0] addr_11765_7;

Selector_2 s11765_7(wires_2941_6[1], addr_2941_6, addr_positional[47063:47060], addr_11765_7);

wire[31:0] addr_11766_7;

Selector_2 s11766_7(wires_2941_6[2], addr_2941_6, addr_positional[47067:47064], addr_11766_7);

wire[31:0] addr_11767_7;

Selector_2 s11767_7(wires_2941_6[3], addr_2941_6, addr_positional[47071:47068], addr_11767_7);

wire[31:0] addr_11768_7;

Selector_2 s11768_7(wires_2942_6[0], addr_2942_6, addr_positional[47075:47072], addr_11768_7);

wire[31:0] addr_11769_7;

Selector_2 s11769_7(wires_2942_6[1], addr_2942_6, addr_positional[47079:47076], addr_11769_7);

wire[31:0] addr_11770_7;

Selector_2 s11770_7(wires_2942_6[2], addr_2942_6, addr_positional[47083:47080], addr_11770_7);

wire[31:0] addr_11771_7;

Selector_2 s11771_7(wires_2942_6[3], addr_2942_6, addr_positional[47087:47084], addr_11771_7);

wire[31:0] addr_11772_7;

Selector_2 s11772_7(wires_2943_6[0], addr_2943_6, addr_positional[47091:47088], addr_11772_7);

wire[31:0] addr_11773_7;

Selector_2 s11773_7(wires_2943_6[1], addr_2943_6, addr_positional[47095:47092], addr_11773_7);

wire[31:0] addr_11774_7;

Selector_2 s11774_7(wires_2943_6[2], addr_2943_6, addr_positional[47099:47096], addr_11774_7);

wire[31:0] addr_11775_7;

Selector_2 s11775_7(wires_2943_6[3], addr_2943_6, addr_positional[47103:47100], addr_11775_7);

wire[31:0] addr_11776_7;

Selector_2 s11776_7(wires_2944_6[0], addr_2944_6, addr_positional[47107:47104], addr_11776_7);

wire[31:0] addr_11777_7;

Selector_2 s11777_7(wires_2944_6[1], addr_2944_6, addr_positional[47111:47108], addr_11777_7);

wire[31:0] addr_11778_7;

Selector_2 s11778_7(wires_2944_6[2], addr_2944_6, addr_positional[47115:47112], addr_11778_7);

wire[31:0] addr_11779_7;

Selector_2 s11779_7(wires_2944_6[3], addr_2944_6, addr_positional[47119:47116], addr_11779_7);

wire[31:0] addr_11780_7;

Selector_2 s11780_7(wires_2945_6[0], addr_2945_6, addr_positional[47123:47120], addr_11780_7);

wire[31:0] addr_11781_7;

Selector_2 s11781_7(wires_2945_6[1], addr_2945_6, addr_positional[47127:47124], addr_11781_7);

wire[31:0] addr_11782_7;

Selector_2 s11782_7(wires_2945_6[2], addr_2945_6, addr_positional[47131:47128], addr_11782_7);

wire[31:0] addr_11783_7;

Selector_2 s11783_7(wires_2945_6[3], addr_2945_6, addr_positional[47135:47132], addr_11783_7);

wire[31:0] addr_11784_7;

Selector_2 s11784_7(wires_2946_6[0], addr_2946_6, addr_positional[47139:47136], addr_11784_7);

wire[31:0] addr_11785_7;

Selector_2 s11785_7(wires_2946_6[1], addr_2946_6, addr_positional[47143:47140], addr_11785_7);

wire[31:0] addr_11786_7;

Selector_2 s11786_7(wires_2946_6[2], addr_2946_6, addr_positional[47147:47144], addr_11786_7);

wire[31:0] addr_11787_7;

Selector_2 s11787_7(wires_2946_6[3], addr_2946_6, addr_positional[47151:47148], addr_11787_7);

wire[31:0] addr_11788_7;

Selector_2 s11788_7(wires_2947_6[0], addr_2947_6, addr_positional[47155:47152], addr_11788_7);

wire[31:0] addr_11789_7;

Selector_2 s11789_7(wires_2947_6[1], addr_2947_6, addr_positional[47159:47156], addr_11789_7);

wire[31:0] addr_11790_7;

Selector_2 s11790_7(wires_2947_6[2], addr_2947_6, addr_positional[47163:47160], addr_11790_7);

wire[31:0] addr_11791_7;

Selector_2 s11791_7(wires_2947_6[3], addr_2947_6, addr_positional[47167:47164], addr_11791_7);

wire[31:0] addr_11792_7;

Selector_2 s11792_7(wires_2948_6[0], addr_2948_6, addr_positional[47171:47168], addr_11792_7);

wire[31:0] addr_11793_7;

Selector_2 s11793_7(wires_2948_6[1], addr_2948_6, addr_positional[47175:47172], addr_11793_7);

wire[31:0] addr_11794_7;

Selector_2 s11794_7(wires_2948_6[2], addr_2948_6, addr_positional[47179:47176], addr_11794_7);

wire[31:0] addr_11795_7;

Selector_2 s11795_7(wires_2948_6[3], addr_2948_6, addr_positional[47183:47180], addr_11795_7);

wire[31:0] addr_11796_7;

Selector_2 s11796_7(wires_2949_6[0], addr_2949_6, addr_positional[47187:47184], addr_11796_7);

wire[31:0] addr_11797_7;

Selector_2 s11797_7(wires_2949_6[1], addr_2949_6, addr_positional[47191:47188], addr_11797_7);

wire[31:0] addr_11798_7;

Selector_2 s11798_7(wires_2949_6[2], addr_2949_6, addr_positional[47195:47192], addr_11798_7);

wire[31:0] addr_11799_7;

Selector_2 s11799_7(wires_2949_6[3], addr_2949_6, addr_positional[47199:47196], addr_11799_7);

wire[31:0] addr_11800_7;

Selector_2 s11800_7(wires_2950_6[0], addr_2950_6, addr_positional[47203:47200], addr_11800_7);

wire[31:0] addr_11801_7;

Selector_2 s11801_7(wires_2950_6[1], addr_2950_6, addr_positional[47207:47204], addr_11801_7);

wire[31:0] addr_11802_7;

Selector_2 s11802_7(wires_2950_6[2], addr_2950_6, addr_positional[47211:47208], addr_11802_7);

wire[31:0] addr_11803_7;

Selector_2 s11803_7(wires_2950_6[3], addr_2950_6, addr_positional[47215:47212], addr_11803_7);

wire[31:0] addr_11804_7;

Selector_2 s11804_7(wires_2951_6[0], addr_2951_6, addr_positional[47219:47216], addr_11804_7);

wire[31:0] addr_11805_7;

Selector_2 s11805_7(wires_2951_6[1], addr_2951_6, addr_positional[47223:47220], addr_11805_7);

wire[31:0] addr_11806_7;

Selector_2 s11806_7(wires_2951_6[2], addr_2951_6, addr_positional[47227:47224], addr_11806_7);

wire[31:0] addr_11807_7;

Selector_2 s11807_7(wires_2951_6[3], addr_2951_6, addr_positional[47231:47228], addr_11807_7);

wire[31:0] addr_11808_7;

Selector_2 s11808_7(wires_2952_6[0], addr_2952_6, addr_positional[47235:47232], addr_11808_7);

wire[31:0] addr_11809_7;

Selector_2 s11809_7(wires_2952_6[1], addr_2952_6, addr_positional[47239:47236], addr_11809_7);

wire[31:0] addr_11810_7;

Selector_2 s11810_7(wires_2952_6[2], addr_2952_6, addr_positional[47243:47240], addr_11810_7);

wire[31:0] addr_11811_7;

Selector_2 s11811_7(wires_2952_6[3], addr_2952_6, addr_positional[47247:47244], addr_11811_7);

wire[31:0] addr_11812_7;

Selector_2 s11812_7(wires_2953_6[0], addr_2953_6, addr_positional[47251:47248], addr_11812_7);

wire[31:0] addr_11813_7;

Selector_2 s11813_7(wires_2953_6[1], addr_2953_6, addr_positional[47255:47252], addr_11813_7);

wire[31:0] addr_11814_7;

Selector_2 s11814_7(wires_2953_6[2], addr_2953_6, addr_positional[47259:47256], addr_11814_7);

wire[31:0] addr_11815_7;

Selector_2 s11815_7(wires_2953_6[3], addr_2953_6, addr_positional[47263:47260], addr_11815_7);

wire[31:0] addr_11816_7;

Selector_2 s11816_7(wires_2954_6[0], addr_2954_6, addr_positional[47267:47264], addr_11816_7);

wire[31:0] addr_11817_7;

Selector_2 s11817_7(wires_2954_6[1], addr_2954_6, addr_positional[47271:47268], addr_11817_7);

wire[31:0] addr_11818_7;

Selector_2 s11818_7(wires_2954_6[2], addr_2954_6, addr_positional[47275:47272], addr_11818_7);

wire[31:0] addr_11819_7;

Selector_2 s11819_7(wires_2954_6[3], addr_2954_6, addr_positional[47279:47276], addr_11819_7);

wire[31:0] addr_11820_7;

Selector_2 s11820_7(wires_2955_6[0], addr_2955_6, addr_positional[47283:47280], addr_11820_7);

wire[31:0] addr_11821_7;

Selector_2 s11821_7(wires_2955_6[1], addr_2955_6, addr_positional[47287:47284], addr_11821_7);

wire[31:0] addr_11822_7;

Selector_2 s11822_7(wires_2955_6[2], addr_2955_6, addr_positional[47291:47288], addr_11822_7);

wire[31:0] addr_11823_7;

Selector_2 s11823_7(wires_2955_6[3], addr_2955_6, addr_positional[47295:47292], addr_11823_7);

wire[31:0] addr_11824_7;

Selector_2 s11824_7(wires_2956_6[0], addr_2956_6, addr_positional[47299:47296], addr_11824_7);

wire[31:0] addr_11825_7;

Selector_2 s11825_7(wires_2956_6[1], addr_2956_6, addr_positional[47303:47300], addr_11825_7);

wire[31:0] addr_11826_7;

Selector_2 s11826_7(wires_2956_6[2], addr_2956_6, addr_positional[47307:47304], addr_11826_7);

wire[31:0] addr_11827_7;

Selector_2 s11827_7(wires_2956_6[3], addr_2956_6, addr_positional[47311:47308], addr_11827_7);

wire[31:0] addr_11828_7;

Selector_2 s11828_7(wires_2957_6[0], addr_2957_6, addr_positional[47315:47312], addr_11828_7);

wire[31:0] addr_11829_7;

Selector_2 s11829_7(wires_2957_6[1], addr_2957_6, addr_positional[47319:47316], addr_11829_7);

wire[31:0] addr_11830_7;

Selector_2 s11830_7(wires_2957_6[2], addr_2957_6, addr_positional[47323:47320], addr_11830_7);

wire[31:0] addr_11831_7;

Selector_2 s11831_7(wires_2957_6[3], addr_2957_6, addr_positional[47327:47324], addr_11831_7);

wire[31:0] addr_11832_7;

Selector_2 s11832_7(wires_2958_6[0], addr_2958_6, addr_positional[47331:47328], addr_11832_7);

wire[31:0] addr_11833_7;

Selector_2 s11833_7(wires_2958_6[1], addr_2958_6, addr_positional[47335:47332], addr_11833_7);

wire[31:0] addr_11834_7;

Selector_2 s11834_7(wires_2958_6[2], addr_2958_6, addr_positional[47339:47336], addr_11834_7);

wire[31:0] addr_11835_7;

Selector_2 s11835_7(wires_2958_6[3], addr_2958_6, addr_positional[47343:47340], addr_11835_7);

wire[31:0] addr_11836_7;

Selector_2 s11836_7(wires_2959_6[0], addr_2959_6, addr_positional[47347:47344], addr_11836_7);

wire[31:0] addr_11837_7;

Selector_2 s11837_7(wires_2959_6[1], addr_2959_6, addr_positional[47351:47348], addr_11837_7);

wire[31:0] addr_11838_7;

Selector_2 s11838_7(wires_2959_6[2], addr_2959_6, addr_positional[47355:47352], addr_11838_7);

wire[31:0] addr_11839_7;

Selector_2 s11839_7(wires_2959_6[3], addr_2959_6, addr_positional[47359:47356], addr_11839_7);

wire[31:0] addr_11840_7;

Selector_2 s11840_7(wires_2960_6[0], addr_2960_6, addr_positional[47363:47360], addr_11840_7);

wire[31:0] addr_11841_7;

Selector_2 s11841_7(wires_2960_6[1], addr_2960_6, addr_positional[47367:47364], addr_11841_7);

wire[31:0] addr_11842_7;

Selector_2 s11842_7(wires_2960_6[2], addr_2960_6, addr_positional[47371:47368], addr_11842_7);

wire[31:0] addr_11843_7;

Selector_2 s11843_7(wires_2960_6[3], addr_2960_6, addr_positional[47375:47372], addr_11843_7);

wire[31:0] addr_11844_7;

Selector_2 s11844_7(wires_2961_6[0], addr_2961_6, addr_positional[47379:47376], addr_11844_7);

wire[31:0] addr_11845_7;

Selector_2 s11845_7(wires_2961_6[1], addr_2961_6, addr_positional[47383:47380], addr_11845_7);

wire[31:0] addr_11846_7;

Selector_2 s11846_7(wires_2961_6[2], addr_2961_6, addr_positional[47387:47384], addr_11846_7);

wire[31:0] addr_11847_7;

Selector_2 s11847_7(wires_2961_6[3], addr_2961_6, addr_positional[47391:47388], addr_11847_7);

wire[31:0] addr_11848_7;

Selector_2 s11848_7(wires_2962_6[0], addr_2962_6, addr_positional[47395:47392], addr_11848_7);

wire[31:0] addr_11849_7;

Selector_2 s11849_7(wires_2962_6[1], addr_2962_6, addr_positional[47399:47396], addr_11849_7);

wire[31:0] addr_11850_7;

Selector_2 s11850_7(wires_2962_6[2], addr_2962_6, addr_positional[47403:47400], addr_11850_7);

wire[31:0] addr_11851_7;

Selector_2 s11851_7(wires_2962_6[3], addr_2962_6, addr_positional[47407:47404], addr_11851_7);

wire[31:0] addr_11852_7;

Selector_2 s11852_7(wires_2963_6[0], addr_2963_6, addr_positional[47411:47408], addr_11852_7);

wire[31:0] addr_11853_7;

Selector_2 s11853_7(wires_2963_6[1], addr_2963_6, addr_positional[47415:47412], addr_11853_7);

wire[31:0] addr_11854_7;

Selector_2 s11854_7(wires_2963_6[2], addr_2963_6, addr_positional[47419:47416], addr_11854_7);

wire[31:0] addr_11855_7;

Selector_2 s11855_7(wires_2963_6[3], addr_2963_6, addr_positional[47423:47420], addr_11855_7);

wire[31:0] addr_11856_7;

Selector_2 s11856_7(wires_2964_6[0], addr_2964_6, addr_positional[47427:47424], addr_11856_7);

wire[31:0] addr_11857_7;

Selector_2 s11857_7(wires_2964_6[1], addr_2964_6, addr_positional[47431:47428], addr_11857_7);

wire[31:0] addr_11858_7;

Selector_2 s11858_7(wires_2964_6[2], addr_2964_6, addr_positional[47435:47432], addr_11858_7);

wire[31:0] addr_11859_7;

Selector_2 s11859_7(wires_2964_6[3], addr_2964_6, addr_positional[47439:47436], addr_11859_7);

wire[31:0] addr_11860_7;

Selector_2 s11860_7(wires_2965_6[0], addr_2965_6, addr_positional[47443:47440], addr_11860_7);

wire[31:0] addr_11861_7;

Selector_2 s11861_7(wires_2965_6[1], addr_2965_6, addr_positional[47447:47444], addr_11861_7);

wire[31:0] addr_11862_7;

Selector_2 s11862_7(wires_2965_6[2], addr_2965_6, addr_positional[47451:47448], addr_11862_7);

wire[31:0] addr_11863_7;

Selector_2 s11863_7(wires_2965_6[3], addr_2965_6, addr_positional[47455:47452], addr_11863_7);

wire[31:0] addr_11864_7;

Selector_2 s11864_7(wires_2966_6[0], addr_2966_6, addr_positional[47459:47456], addr_11864_7);

wire[31:0] addr_11865_7;

Selector_2 s11865_7(wires_2966_6[1], addr_2966_6, addr_positional[47463:47460], addr_11865_7);

wire[31:0] addr_11866_7;

Selector_2 s11866_7(wires_2966_6[2], addr_2966_6, addr_positional[47467:47464], addr_11866_7);

wire[31:0] addr_11867_7;

Selector_2 s11867_7(wires_2966_6[3], addr_2966_6, addr_positional[47471:47468], addr_11867_7);

wire[31:0] addr_11868_7;

Selector_2 s11868_7(wires_2967_6[0], addr_2967_6, addr_positional[47475:47472], addr_11868_7);

wire[31:0] addr_11869_7;

Selector_2 s11869_7(wires_2967_6[1], addr_2967_6, addr_positional[47479:47476], addr_11869_7);

wire[31:0] addr_11870_7;

Selector_2 s11870_7(wires_2967_6[2], addr_2967_6, addr_positional[47483:47480], addr_11870_7);

wire[31:0] addr_11871_7;

Selector_2 s11871_7(wires_2967_6[3], addr_2967_6, addr_positional[47487:47484], addr_11871_7);

wire[31:0] addr_11872_7;

Selector_2 s11872_7(wires_2968_6[0], addr_2968_6, addr_positional[47491:47488], addr_11872_7);

wire[31:0] addr_11873_7;

Selector_2 s11873_7(wires_2968_6[1], addr_2968_6, addr_positional[47495:47492], addr_11873_7);

wire[31:0] addr_11874_7;

Selector_2 s11874_7(wires_2968_6[2], addr_2968_6, addr_positional[47499:47496], addr_11874_7);

wire[31:0] addr_11875_7;

Selector_2 s11875_7(wires_2968_6[3], addr_2968_6, addr_positional[47503:47500], addr_11875_7);

wire[31:0] addr_11876_7;

Selector_2 s11876_7(wires_2969_6[0], addr_2969_6, addr_positional[47507:47504], addr_11876_7);

wire[31:0] addr_11877_7;

Selector_2 s11877_7(wires_2969_6[1], addr_2969_6, addr_positional[47511:47508], addr_11877_7);

wire[31:0] addr_11878_7;

Selector_2 s11878_7(wires_2969_6[2], addr_2969_6, addr_positional[47515:47512], addr_11878_7);

wire[31:0] addr_11879_7;

Selector_2 s11879_7(wires_2969_6[3], addr_2969_6, addr_positional[47519:47516], addr_11879_7);

wire[31:0] addr_11880_7;

Selector_2 s11880_7(wires_2970_6[0], addr_2970_6, addr_positional[47523:47520], addr_11880_7);

wire[31:0] addr_11881_7;

Selector_2 s11881_7(wires_2970_6[1], addr_2970_6, addr_positional[47527:47524], addr_11881_7);

wire[31:0] addr_11882_7;

Selector_2 s11882_7(wires_2970_6[2], addr_2970_6, addr_positional[47531:47528], addr_11882_7);

wire[31:0] addr_11883_7;

Selector_2 s11883_7(wires_2970_6[3], addr_2970_6, addr_positional[47535:47532], addr_11883_7);

wire[31:0] addr_11884_7;

Selector_2 s11884_7(wires_2971_6[0], addr_2971_6, addr_positional[47539:47536], addr_11884_7);

wire[31:0] addr_11885_7;

Selector_2 s11885_7(wires_2971_6[1], addr_2971_6, addr_positional[47543:47540], addr_11885_7);

wire[31:0] addr_11886_7;

Selector_2 s11886_7(wires_2971_6[2], addr_2971_6, addr_positional[47547:47544], addr_11886_7);

wire[31:0] addr_11887_7;

Selector_2 s11887_7(wires_2971_6[3], addr_2971_6, addr_positional[47551:47548], addr_11887_7);

wire[31:0] addr_11888_7;

Selector_2 s11888_7(wires_2972_6[0], addr_2972_6, addr_positional[47555:47552], addr_11888_7);

wire[31:0] addr_11889_7;

Selector_2 s11889_7(wires_2972_6[1], addr_2972_6, addr_positional[47559:47556], addr_11889_7);

wire[31:0] addr_11890_7;

Selector_2 s11890_7(wires_2972_6[2], addr_2972_6, addr_positional[47563:47560], addr_11890_7);

wire[31:0] addr_11891_7;

Selector_2 s11891_7(wires_2972_6[3], addr_2972_6, addr_positional[47567:47564], addr_11891_7);

wire[31:0] addr_11892_7;

Selector_2 s11892_7(wires_2973_6[0], addr_2973_6, addr_positional[47571:47568], addr_11892_7);

wire[31:0] addr_11893_7;

Selector_2 s11893_7(wires_2973_6[1], addr_2973_6, addr_positional[47575:47572], addr_11893_7);

wire[31:0] addr_11894_7;

Selector_2 s11894_7(wires_2973_6[2], addr_2973_6, addr_positional[47579:47576], addr_11894_7);

wire[31:0] addr_11895_7;

Selector_2 s11895_7(wires_2973_6[3], addr_2973_6, addr_positional[47583:47580], addr_11895_7);

wire[31:0] addr_11896_7;

Selector_2 s11896_7(wires_2974_6[0], addr_2974_6, addr_positional[47587:47584], addr_11896_7);

wire[31:0] addr_11897_7;

Selector_2 s11897_7(wires_2974_6[1], addr_2974_6, addr_positional[47591:47588], addr_11897_7);

wire[31:0] addr_11898_7;

Selector_2 s11898_7(wires_2974_6[2], addr_2974_6, addr_positional[47595:47592], addr_11898_7);

wire[31:0] addr_11899_7;

Selector_2 s11899_7(wires_2974_6[3], addr_2974_6, addr_positional[47599:47596], addr_11899_7);

wire[31:0] addr_11900_7;

Selector_2 s11900_7(wires_2975_6[0], addr_2975_6, addr_positional[47603:47600], addr_11900_7);

wire[31:0] addr_11901_7;

Selector_2 s11901_7(wires_2975_6[1], addr_2975_6, addr_positional[47607:47604], addr_11901_7);

wire[31:0] addr_11902_7;

Selector_2 s11902_7(wires_2975_6[2], addr_2975_6, addr_positional[47611:47608], addr_11902_7);

wire[31:0] addr_11903_7;

Selector_2 s11903_7(wires_2975_6[3], addr_2975_6, addr_positional[47615:47612], addr_11903_7);

wire[31:0] addr_11904_7;

Selector_2 s11904_7(wires_2976_6[0], addr_2976_6, addr_positional[47619:47616], addr_11904_7);

wire[31:0] addr_11905_7;

Selector_2 s11905_7(wires_2976_6[1], addr_2976_6, addr_positional[47623:47620], addr_11905_7);

wire[31:0] addr_11906_7;

Selector_2 s11906_7(wires_2976_6[2], addr_2976_6, addr_positional[47627:47624], addr_11906_7);

wire[31:0] addr_11907_7;

Selector_2 s11907_7(wires_2976_6[3], addr_2976_6, addr_positional[47631:47628], addr_11907_7);

wire[31:0] addr_11908_7;

Selector_2 s11908_7(wires_2977_6[0], addr_2977_6, addr_positional[47635:47632], addr_11908_7);

wire[31:0] addr_11909_7;

Selector_2 s11909_7(wires_2977_6[1], addr_2977_6, addr_positional[47639:47636], addr_11909_7);

wire[31:0] addr_11910_7;

Selector_2 s11910_7(wires_2977_6[2], addr_2977_6, addr_positional[47643:47640], addr_11910_7);

wire[31:0] addr_11911_7;

Selector_2 s11911_7(wires_2977_6[3], addr_2977_6, addr_positional[47647:47644], addr_11911_7);

wire[31:0] addr_11912_7;

Selector_2 s11912_7(wires_2978_6[0], addr_2978_6, addr_positional[47651:47648], addr_11912_7);

wire[31:0] addr_11913_7;

Selector_2 s11913_7(wires_2978_6[1], addr_2978_6, addr_positional[47655:47652], addr_11913_7);

wire[31:0] addr_11914_7;

Selector_2 s11914_7(wires_2978_6[2], addr_2978_6, addr_positional[47659:47656], addr_11914_7);

wire[31:0] addr_11915_7;

Selector_2 s11915_7(wires_2978_6[3], addr_2978_6, addr_positional[47663:47660], addr_11915_7);

wire[31:0] addr_11916_7;

Selector_2 s11916_7(wires_2979_6[0], addr_2979_6, addr_positional[47667:47664], addr_11916_7);

wire[31:0] addr_11917_7;

Selector_2 s11917_7(wires_2979_6[1], addr_2979_6, addr_positional[47671:47668], addr_11917_7);

wire[31:0] addr_11918_7;

Selector_2 s11918_7(wires_2979_6[2], addr_2979_6, addr_positional[47675:47672], addr_11918_7);

wire[31:0] addr_11919_7;

Selector_2 s11919_7(wires_2979_6[3], addr_2979_6, addr_positional[47679:47676], addr_11919_7);

wire[31:0] addr_11920_7;

Selector_2 s11920_7(wires_2980_6[0], addr_2980_6, addr_positional[47683:47680], addr_11920_7);

wire[31:0] addr_11921_7;

Selector_2 s11921_7(wires_2980_6[1], addr_2980_6, addr_positional[47687:47684], addr_11921_7);

wire[31:0] addr_11922_7;

Selector_2 s11922_7(wires_2980_6[2], addr_2980_6, addr_positional[47691:47688], addr_11922_7);

wire[31:0] addr_11923_7;

Selector_2 s11923_7(wires_2980_6[3], addr_2980_6, addr_positional[47695:47692], addr_11923_7);

wire[31:0] addr_11924_7;

Selector_2 s11924_7(wires_2981_6[0], addr_2981_6, addr_positional[47699:47696], addr_11924_7);

wire[31:0] addr_11925_7;

Selector_2 s11925_7(wires_2981_6[1], addr_2981_6, addr_positional[47703:47700], addr_11925_7);

wire[31:0] addr_11926_7;

Selector_2 s11926_7(wires_2981_6[2], addr_2981_6, addr_positional[47707:47704], addr_11926_7);

wire[31:0] addr_11927_7;

Selector_2 s11927_7(wires_2981_6[3], addr_2981_6, addr_positional[47711:47708], addr_11927_7);

wire[31:0] addr_11928_7;

Selector_2 s11928_7(wires_2982_6[0], addr_2982_6, addr_positional[47715:47712], addr_11928_7);

wire[31:0] addr_11929_7;

Selector_2 s11929_7(wires_2982_6[1], addr_2982_6, addr_positional[47719:47716], addr_11929_7);

wire[31:0] addr_11930_7;

Selector_2 s11930_7(wires_2982_6[2], addr_2982_6, addr_positional[47723:47720], addr_11930_7);

wire[31:0] addr_11931_7;

Selector_2 s11931_7(wires_2982_6[3], addr_2982_6, addr_positional[47727:47724], addr_11931_7);

wire[31:0] addr_11932_7;

Selector_2 s11932_7(wires_2983_6[0], addr_2983_6, addr_positional[47731:47728], addr_11932_7);

wire[31:0] addr_11933_7;

Selector_2 s11933_7(wires_2983_6[1], addr_2983_6, addr_positional[47735:47732], addr_11933_7);

wire[31:0] addr_11934_7;

Selector_2 s11934_7(wires_2983_6[2], addr_2983_6, addr_positional[47739:47736], addr_11934_7);

wire[31:0] addr_11935_7;

Selector_2 s11935_7(wires_2983_6[3], addr_2983_6, addr_positional[47743:47740], addr_11935_7);

wire[31:0] addr_11936_7;

Selector_2 s11936_7(wires_2984_6[0], addr_2984_6, addr_positional[47747:47744], addr_11936_7);

wire[31:0] addr_11937_7;

Selector_2 s11937_7(wires_2984_6[1], addr_2984_6, addr_positional[47751:47748], addr_11937_7);

wire[31:0] addr_11938_7;

Selector_2 s11938_7(wires_2984_6[2], addr_2984_6, addr_positional[47755:47752], addr_11938_7);

wire[31:0] addr_11939_7;

Selector_2 s11939_7(wires_2984_6[3], addr_2984_6, addr_positional[47759:47756], addr_11939_7);

wire[31:0] addr_11940_7;

Selector_2 s11940_7(wires_2985_6[0], addr_2985_6, addr_positional[47763:47760], addr_11940_7);

wire[31:0] addr_11941_7;

Selector_2 s11941_7(wires_2985_6[1], addr_2985_6, addr_positional[47767:47764], addr_11941_7);

wire[31:0] addr_11942_7;

Selector_2 s11942_7(wires_2985_6[2], addr_2985_6, addr_positional[47771:47768], addr_11942_7);

wire[31:0] addr_11943_7;

Selector_2 s11943_7(wires_2985_6[3], addr_2985_6, addr_positional[47775:47772], addr_11943_7);

wire[31:0] addr_11944_7;

Selector_2 s11944_7(wires_2986_6[0], addr_2986_6, addr_positional[47779:47776], addr_11944_7);

wire[31:0] addr_11945_7;

Selector_2 s11945_7(wires_2986_6[1], addr_2986_6, addr_positional[47783:47780], addr_11945_7);

wire[31:0] addr_11946_7;

Selector_2 s11946_7(wires_2986_6[2], addr_2986_6, addr_positional[47787:47784], addr_11946_7);

wire[31:0] addr_11947_7;

Selector_2 s11947_7(wires_2986_6[3], addr_2986_6, addr_positional[47791:47788], addr_11947_7);

wire[31:0] addr_11948_7;

Selector_2 s11948_7(wires_2987_6[0], addr_2987_6, addr_positional[47795:47792], addr_11948_7);

wire[31:0] addr_11949_7;

Selector_2 s11949_7(wires_2987_6[1], addr_2987_6, addr_positional[47799:47796], addr_11949_7);

wire[31:0] addr_11950_7;

Selector_2 s11950_7(wires_2987_6[2], addr_2987_6, addr_positional[47803:47800], addr_11950_7);

wire[31:0] addr_11951_7;

Selector_2 s11951_7(wires_2987_6[3], addr_2987_6, addr_positional[47807:47804], addr_11951_7);

wire[31:0] addr_11952_7;

Selector_2 s11952_7(wires_2988_6[0], addr_2988_6, addr_positional[47811:47808], addr_11952_7);

wire[31:0] addr_11953_7;

Selector_2 s11953_7(wires_2988_6[1], addr_2988_6, addr_positional[47815:47812], addr_11953_7);

wire[31:0] addr_11954_7;

Selector_2 s11954_7(wires_2988_6[2], addr_2988_6, addr_positional[47819:47816], addr_11954_7);

wire[31:0] addr_11955_7;

Selector_2 s11955_7(wires_2988_6[3], addr_2988_6, addr_positional[47823:47820], addr_11955_7);

wire[31:0] addr_11956_7;

Selector_2 s11956_7(wires_2989_6[0], addr_2989_6, addr_positional[47827:47824], addr_11956_7);

wire[31:0] addr_11957_7;

Selector_2 s11957_7(wires_2989_6[1], addr_2989_6, addr_positional[47831:47828], addr_11957_7);

wire[31:0] addr_11958_7;

Selector_2 s11958_7(wires_2989_6[2], addr_2989_6, addr_positional[47835:47832], addr_11958_7);

wire[31:0] addr_11959_7;

Selector_2 s11959_7(wires_2989_6[3], addr_2989_6, addr_positional[47839:47836], addr_11959_7);

wire[31:0] addr_11960_7;

Selector_2 s11960_7(wires_2990_6[0], addr_2990_6, addr_positional[47843:47840], addr_11960_7);

wire[31:0] addr_11961_7;

Selector_2 s11961_7(wires_2990_6[1], addr_2990_6, addr_positional[47847:47844], addr_11961_7);

wire[31:0] addr_11962_7;

Selector_2 s11962_7(wires_2990_6[2], addr_2990_6, addr_positional[47851:47848], addr_11962_7);

wire[31:0] addr_11963_7;

Selector_2 s11963_7(wires_2990_6[3], addr_2990_6, addr_positional[47855:47852], addr_11963_7);

wire[31:0] addr_11964_7;

Selector_2 s11964_7(wires_2991_6[0], addr_2991_6, addr_positional[47859:47856], addr_11964_7);

wire[31:0] addr_11965_7;

Selector_2 s11965_7(wires_2991_6[1], addr_2991_6, addr_positional[47863:47860], addr_11965_7);

wire[31:0] addr_11966_7;

Selector_2 s11966_7(wires_2991_6[2], addr_2991_6, addr_positional[47867:47864], addr_11966_7);

wire[31:0] addr_11967_7;

Selector_2 s11967_7(wires_2991_6[3], addr_2991_6, addr_positional[47871:47868], addr_11967_7);

wire[31:0] addr_11968_7;

Selector_2 s11968_7(wires_2992_6[0], addr_2992_6, addr_positional[47875:47872], addr_11968_7);

wire[31:0] addr_11969_7;

Selector_2 s11969_7(wires_2992_6[1], addr_2992_6, addr_positional[47879:47876], addr_11969_7);

wire[31:0] addr_11970_7;

Selector_2 s11970_7(wires_2992_6[2], addr_2992_6, addr_positional[47883:47880], addr_11970_7);

wire[31:0] addr_11971_7;

Selector_2 s11971_7(wires_2992_6[3], addr_2992_6, addr_positional[47887:47884], addr_11971_7);

wire[31:0] addr_11972_7;

Selector_2 s11972_7(wires_2993_6[0], addr_2993_6, addr_positional[47891:47888], addr_11972_7);

wire[31:0] addr_11973_7;

Selector_2 s11973_7(wires_2993_6[1], addr_2993_6, addr_positional[47895:47892], addr_11973_7);

wire[31:0] addr_11974_7;

Selector_2 s11974_7(wires_2993_6[2], addr_2993_6, addr_positional[47899:47896], addr_11974_7);

wire[31:0] addr_11975_7;

Selector_2 s11975_7(wires_2993_6[3], addr_2993_6, addr_positional[47903:47900], addr_11975_7);

wire[31:0] addr_11976_7;

Selector_2 s11976_7(wires_2994_6[0], addr_2994_6, addr_positional[47907:47904], addr_11976_7);

wire[31:0] addr_11977_7;

Selector_2 s11977_7(wires_2994_6[1], addr_2994_6, addr_positional[47911:47908], addr_11977_7);

wire[31:0] addr_11978_7;

Selector_2 s11978_7(wires_2994_6[2], addr_2994_6, addr_positional[47915:47912], addr_11978_7);

wire[31:0] addr_11979_7;

Selector_2 s11979_7(wires_2994_6[3], addr_2994_6, addr_positional[47919:47916], addr_11979_7);

wire[31:0] addr_11980_7;

Selector_2 s11980_7(wires_2995_6[0], addr_2995_6, addr_positional[47923:47920], addr_11980_7);

wire[31:0] addr_11981_7;

Selector_2 s11981_7(wires_2995_6[1], addr_2995_6, addr_positional[47927:47924], addr_11981_7);

wire[31:0] addr_11982_7;

Selector_2 s11982_7(wires_2995_6[2], addr_2995_6, addr_positional[47931:47928], addr_11982_7);

wire[31:0] addr_11983_7;

Selector_2 s11983_7(wires_2995_6[3], addr_2995_6, addr_positional[47935:47932], addr_11983_7);

wire[31:0] addr_11984_7;

Selector_2 s11984_7(wires_2996_6[0], addr_2996_6, addr_positional[47939:47936], addr_11984_7);

wire[31:0] addr_11985_7;

Selector_2 s11985_7(wires_2996_6[1], addr_2996_6, addr_positional[47943:47940], addr_11985_7);

wire[31:0] addr_11986_7;

Selector_2 s11986_7(wires_2996_6[2], addr_2996_6, addr_positional[47947:47944], addr_11986_7);

wire[31:0] addr_11987_7;

Selector_2 s11987_7(wires_2996_6[3], addr_2996_6, addr_positional[47951:47948], addr_11987_7);

wire[31:0] addr_11988_7;

Selector_2 s11988_7(wires_2997_6[0], addr_2997_6, addr_positional[47955:47952], addr_11988_7);

wire[31:0] addr_11989_7;

Selector_2 s11989_7(wires_2997_6[1], addr_2997_6, addr_positional[47959:47956], addr_11989_7);

wire[31:0] addr_11990_7;

Selector_2 s11990_7(wires_2997_6[2], addr_2997_6, addr_positional[47963:47960], addr_11990_7);

wire[31:0] addr_11991_7;

Selector_2 s11991_7(wires_2997_6[3], addr_2997_6, addr_positional[47967:47964], addr_11991_7);

wire[31:0] addr_11992_7;

Selector_2 s11992_7(wires_2998_6[0], addr_2998_6, addr_positional[47971:47968], addr_11992_7);

wire[31:0] addr_11993_7;

Selector_2 s11993_7(wires_2998_6[1], addr_2998_6, addr_positional[47975:47972], addr_11993_7);

wire[31:0] addr_11994_7;

Selector_2 s11994_7(wires_2998_6[2], addr_2998_6, addr_positional[47979:47976], addr_11994_7);

wire[31:0] addr_11995_7;

Selector_2 s11995_7(wires_2998_6[3], addr_2998_6, addr_positional[47983:47980], addr_11995_7);

wire[31:0] addr_11996_7;

Selector_2 s11996_7(wires_2999_6[0], addr_2999_6, addr_positional[47987:47984], addr_11996_7);

wire[31:0] addr_11997_7;

Selector_2 s11997_7(wires_2999_6[1], addr_2999_6, addr_positional[47991:47988], addr_11997_7);

wire[31:0] addr_11998_7;

Selector_2 s11998_7(wires_2999_6[2], addr_2999_6, addr_positional[47995:47992], addr_11998_7);

wire[31:0] addr_11999_7;

Selector_2 s11999_7(wires_2999_6[3], addr_2999_6, addr_positional[47999:47996], addr_11999_7);

wire[31:0] addr_12000_7;

Selector_2 s12000_7(wires_3000_6[0], addr_3000_6, addr_positional[48003:48000], addr_12000_7);

wire[31:0] addr_12001_7;

Selector_2 s12001_7(wires_3000_6[1], addr_3000_6, addr_positional[48007:48004], addr_12001_7);

wire[31:0] addr_12002_7;

Selector_2 s12002_7(wires_3000_6[2], addr_3000_6, addr_positional[48011:48008], addr_12002_7);

wire[31:0] addr_12003_7;

Selector_2 s12003_7(wires_3000_6[3], addr_3000_6, addr_positional[48015:48012], addr_12003_7);

wire[31:0] addr_12004_7;

Selector_2 s12004_7(wires_3001_6[0], addr_3001_6, addr_positional[48019:48016], addr_12004_7);

wire[31:0] addr_12005_7;

Selector_2 s12005_7(wires_3001_6[1], addr_3001_6, addr_positional[48023:48020], addr_12005_7);

wire[31:0] addr_12006_7;

Selector_2 s12006_7(wires_3001_6[2], addr_3001_6, addr_positional[48027:48024], addr_12006_7);

wire[31:0] addr_12007_7;

Selector_2 s12007_7(wires_3001_6[3], addr_3001_6, addr_positional[48031:48028], addr_12007_7);

wire[31:0] addr_12008_7;

Selector_2 s12008_7(wires_3002_6[0], addr_3002_6, addr_positional[48035:48032], addr_12008_7);

wire[31:0] addr_12009_7;

Selector_2 s12009_7(wires_3002_6[1], addr_3002_6, addr_positional[48039:48036], addr_12009_7);

wire[31:0] addr_12010_7;

Selector_2 s12010_7(wires_3002_6[2], addr_3002_6, addr_positional[48043:48040], addr_12010_7);

wire[31:0] addr_12011_7;

Selector_2 s12011_7(wires_3002_6[3], addr_3002_6, addr_positional[48047:48044], addr_12011_7);

wire[31:0] addr_12012_7;

Selector_2 s12012_7(wires_3003_6[0], addr_3003_6, addr_positional[48051:48048], addr_12012_7);

wire[31:0] addr_12013_7;

Selector_2 s12013_7(wires_3003_6[1], addr_3003_6, addr_positional[48055:48052], addr_12013_7);

wire[31:0] addr_12014_7;

Selector_2 s12014_7(wires_3003_6[2], addr_3003_6, addr_positional[48059:48056], addr_12014_7);

wire[31:0] addr_12015_7;

Selector_2 s12015_7(wires_3003_6[3], addr_3003_6, addr_positional[48063:48060], addr_12015_7);

wire[31:0] addr_12016_7;

Selector_2 s12016_7(wires_3004_6[0], addr_3004_6, addr_positional[48067:48064], addr_12016_7);

wire[31:0] addr_12017_7;

Selector_2 s12017_7(wires_3004_6[1], addr_3004_6, addr_positional[48071:48068], addr_12017_7);

wire[31:0] addr_12018_7;

Selector_2 s12018_7(wires_3004_6[2], addr_3004_6, addr_positional[48075:48072], addr_12018_7);

wire[31:0] addr_12019_7;

Selector_2 s12019_7(wires_3004_6[3], addr_3004_6, addr_positional[48079:48076], addr_12019_7);

wire[31:0] addr_12020_7;

Selector_2 s12020_7(wires_3005_6[0], addr_3005_6, addr_positional[48083:48080], addr_12020_7);

wire[31:0] addr_12021_7;

Selector_2 s12021_7(wires_3005_6[1], addr_3005_6, addr_positional[48087:48084], addr_12021_7);

wire[31:0] addr_12022_7;

Selector_2 s12022_7(wires_3005_6[2], addr_3005_6, addr_positional[48091:48088], addr_12022_7);

wire[31:0] addr_12023_7;

Selector_2 s12023_7(wires_3005_6[3], addr_3005_6, addr_positional[48095:48092], addr_12023_7);

wire[31:0] addr_12024_7;

Selector_2 s12024_7(wires_3006_6[0], addr_3006_6, addr_positional[48099:48096], addr_12024_7);

wire[31:0] addr_12025_7;

Selector_2 s12025_7(wires_3006_6[1], addr_3006_6, addr_positional[48103:48100], addr_12025_7);

wire[31:0] addr_12026_7;

Selector_2 s12026_7(wires_3006_6[2], addr_3006_6, addr_positional[48107:48104], addr_12026_7);

wire[31:0] addr_12027_7;

Selector_2 s12027_7(wires_3006_6[3], addr_3006_6, addr_positional[48111:48108], addr_12027_7);

wire[31:0] addr_12028_7;

Selector_2 s12028_7(wires_3007_6[0], addr_3007_6, addr_positional[48115:48112], addr_12028_7);

wire[31:0] addr_12029_7;

Selector_2 s12029_7(wires_3007_6[1], addr_3007_6, addr_positional[48119:48116], addr_12029_7);

wire[31:0] addr_12030_7;

Selector_2 s12030_7(wires_3007_6[2], addr_3007_6, addr_positional[48123:48120], addr_12030_7);

wire[31:0] addr_12031_7;

Selector_2 s12031_7(wires_3007_6[3], addr_3007_6, addr_positional[48127:48124], addr_12031_7);

wire[31:0] addr_12032_7;

Selector_2 s12032_7(wires_3008_6[0], addr_3008_6, addr_positional[48131:48128], addr_12032_7);

wire[31:0] addr_12033_7;

Selector_2 s12033_7(wires_3008_6[1], addr_3008_6, addr_positional[48135:48132], addr_12033_7);

wire[31:0] addr_12034_7;

Selector_2 s12034_7(wires_3008_6[2], addr_3008_6, addr_positional[48139:48136], addr_12034_7);

wire[31:0] addr_12035_7;

Selector_2 s12035_7(wires_3008_6[3], addr_3008_6, addr_positional[48143:48140], addr_12035_7);

wire[31:0] addr_12036_7;

Selector_2 s12036_7(wires_3009_6[0], addr_3009_6, addr_positional[48147:48144], addr_12036_7);

wire[31:0] addr_12037_7;

Selector_2 s12037_7(wires_3009_6[1], addr_3009_6, addr_positional[48151:48148], addr_12037_7);

wire[31:0] addr_12038_7;

Selector_2 s12038_7(wires_3009_6[2], addr_3009_6, addr_positional[48155:48152], addr_12038_7);

wire[31:0] addr_12039_7;

Selector_2 s12039_7(wires_3009_6[3], addr_3009_6, addr_positional[48159:48156], addr_12039_7);

wire[31:0] addr_12040_7;

Selector_2 s12040_7(wires_3010_6[0], addr_3010_6, addr_positional[48163:48160], addr_12040_7);

wire[31:0] addr_12041_7;

Selector_2 s12041_7(wires_3010_6[1], addr_3010_6, addr_positional[48167:48164], addr_12041_7);

wire[31:0] addr_12042_7;

Selector_2 s12042_7(wires_3010_6[2], addr_3010_6, addr_positional[48171:48168], addr_12042_7);

wire[31:0] addr_12043_7;

Selector_2 s12043_7(wires_3010_6[3], addr_3010_6, addr_positional[48175:48172], addr_12043_7);

wire[31:0] addr_12044_7;

Selector_2 s12044_7(wires_3011_6[0], addr_3011_6, addr_positional[48179:48176], addr_12044_7);

wire[31:0] addr_12045_7;

Selector_2 s12045_7(wires_3011_6[1], addr_3011_6, addr_positional[48183:48180], addr_12045_7);

wire[31:0] addr_12046_7;

Selector_2 s12046_7(wires_3011_6[2], addr_3011_6, addr_positional[48187:48184], addr_12046_7);

wire[31:0] addr_12047_7;

Selector_2 s12047_7(wires_3011_6[3], addr_3011_6, addr_positional[48191:48188], addr_12047_7);

wire[31:0] addr_12048_7;

Selector_2 s12048_7(wires_3012_6[0], addr_3012_6, addr_positional[48195:48192], addr_12048_7);

wire[31:0] addr_12049_7;

Selector_2 s12049_7(wires_3012_6[1], addr_3012_6, addr_positional[48199:48196], addr_12049_7);

wire[31:0] addr_12050_7;

Selector_2 s12050_7(wires_3012_6[2], addr_3012_6, addr_positional[48203:48200], addr_12050_7);

wire[31:0] addr_12051_7;

Selector_2 s12051_7(wires_3012_6[3], addr_3012_6, addr_positional[48207:48204], addr_12051_7);

wire[31:0] addr_12052_7;

Selector_2 s12052_7(wires_3013_6[0], addr_3013_6, addr_positional[48211:48208], addr_12052_7);

wire[31:0] addr_12053_7;

Selector_2 s12053_7(wires_3013_6[1], addr_3013_6, addr_positional[48215:48212], addr_12053_7);

wire[31:0] addr_12054_7;

Selector_2 s12054_7(wires_3013_6[2], addr_3013_6, addr_positional[48219:48216], addr_12054_7);

wire[31:0] addr_12055_7;

Selector_2 s12055_7(wires_3013_6[3], addr_3013_6, addr_positional[48223:48220], addr_12055_7);

wire[31:0] addr_12056_7;

Selector_2 s12056_7(wires_3014_6[0], addr_3014_6, addr_positional[48227:48224], addr_12056_7);

wire[31:0] addr_12057_7;

Selector_2 s12057_7(wires_3014_6[1], addr_3014_6, addr_positional[48231:48228], addr_12057_7);

wire[31:0] addr_12058_7;

Selector_2 s12058_7(wires_3014_6[2], addr_3014_6, addr_positional[48235:48232], addr_12058_7);

wire[31:0] addr_12059_7;

Selector_2 s12059_7(wires_3014_6[3], addr_3014_6, addr_positional[48239:48236], addr_12059_7);

wire[31:0] addr_12060_7;

Selector_2 s12060_7(wires_3015_6[0], addr_3015_6, addr_positional[48243:48240], addr_12060_7);

wire[31:0] addr_12061_7;

Selector_2 s12061_7(wires_3015_6[1], addr_3015_6, addr_positional[48247:48244], addr_12061_7);

wire[31:0] addr_12062_7;

Selector_2 s12062_7(wires_3015_6[2], addr_3015_6, addr_positional[48251:48248], addr_12062_7);

wire[31:0] addr_12063_7;

Selector_2 s12063_7(wires_3015_6[3], addr_3015_6, addr_positional[48255:48252], addr_12063_7);

wire[31:0] addr_12064_7;

Selector_2 s12064_7(wires_3016_6[0], addr_3016_6, addr_positional[48259:48256], addr_12064_7);

wire[31:0] addr_12065_7;

Selector_2 s12065_7(wires_3016_6[1], addr_3016_6, addr_positional[48263:48260], addr_12065_7);

wire[31:0] addr_12066_7;

Selector_2 s12066_7(wires_3016_6[2], addr_3016_6, addr_positional[48267:48264], addr_12066_7);

wire[31:0] addr_12067_7;

Selector_2 s12067_7(wires_3016_6[3], addr_3016_6, addr_positional[48271:48268], addr_12067_7);

wire[31:0] addr_12068_7;

Selector_2 s12068_7(wires_3017_6[0], addr_3017_6, addr_positional[48275:48272], addr_12068_7);

wire[31:0] addr_12069_7;

Selector_2 s12069_7(wires_3017_6[1], addr_3017_6, addr_positional[48279:48276], addr_12069_7);

wire[31:0] addr_12070_7;

Selector_2 s12070_7(wires_3017_6[2], addr_3017_6, addr_positional[48283:48280], addr_12070_7);

wire[31:0] addr_12071_7;

Selector_2 s12071_7(wires_3017_6[3], addr_3017_6, addr_positional[48287:48284], addr_12071_7);

wire[31:0] addr_12072_7;

Selector_2 s12072_7(wires_3018_6[0], addr_3018_6, addr_positional[48291:48288], addr_12072_7);

wire[31:0] addr_12073_7;

Selector_2 s12073_7(wires_3018_6[1], addr_3018_6, addr_positional[48295:48292], addr_12073_7);

wire[31:0] addr_12074_7;

Selector_2 s12074_7(wires_3018_6[2], addr_3018_6, addr_positional[48299:48296], addr_12074_7);

wire[31:0] addr_12075_7;

Selector_2 s12075_7(wires_3018_6[3], addr_3018_6, addr_positional[48303:48300], addr_12075_7);

wire[31:0] addr_12076_7;

Selector_2 s12076_7(wires_3019_6[0], addr_3019_6, addr_positional[48307:48304], addr_12076_7);

wire[31:0] addr_12077_7;

Selector_2 s12077_7(wires_3019_6[1], addr_3019_6, addr_positional[48311:48308], addr_12077_7);

wire[31:0] addr_12078_7;

Selector_2 s12078_7(wires_3019_6[2], addr_3019_6, addr_positional[48315:48312], addr_12078_7);

wire[31:0] addr_12079_7;

Selector_2 s12079_7(wires_3019_6[3], addr_3019_6, addr_positional[48319:48316], addr_12079_7);

wire[31:0] addr_12080_7;

Selector_2 s12080_7(wires_3020_6[0], addr_3020_6, addr_positional[48323:48320], addr_12080_7);

wire[31:0] addr_12081_7;

Selector_2 s12081_7(wires_3020_6[1], addr_3020_6, addr_positional[48327:48324], addr_12081_7);

wire[31:0] addr_12082_7;

Selector_2 s12082_7(wires_3020_6[2], addr_3020_6, addr_positional[48331:48328], addr_12082_7);

wire[31:0] addr_12083_7;

Selector_2 s12083_7(wires_3020_6[3], addr_3020_6, addr_positional[48335:48332], addr_12083_7);

wire[31:0] addr_12084_7;

Selector_2 s12084_7(wires_3021_6[0], addr_3021_6, addr_positional[48339:48336], addr_12084_7);

wire[31:0] addr_12085_7;

Selector_2 s12085_7(wires_3021_6[1], addr_3021_6, addr_positional[48343:48340], addr_12085_7);

wire[31:0] addr_12086_7;

Selector_2 s12086_7(wires_3021_6[2], addr_3021_6, addr_positional[48347:48344], addr_12086_7);

wire[31:0] addr_12087_7;

Selector_2 s12087_7(wires_3021_6[3], addr_3021_6, addr_positional[48351:48348], addr_12087_7);

wire[31:0] addr_12088_7;

Selector_2 s12088_7(wires_3022_6[0], addr_3022_6, addr_positional[48355:48352], addr_12088_7);

wire[31:0] addr_12089_7;

Selector_2 s12089_7(wires_3022_6[1], addr_3022_6, addr_positional[48359:48356], addr_12089_7);

wire[31:0] addr_12090_7;

Selector_2 s12090_7(wires_3022_6[2], addr_3022_6, addr_positional[48363:48360], addr_12090_7);

wire[31:0] addr_12091_7;

Selector_2 s12091_7(wires_3022_6[3], addr_3022_6, addr_positional[48367:48364], addr_12091_7);

wire[31:0] addr_12092_7;

Selector_2 s12092_7(wires_3023_6[0], addr_3023_6, addr_positional[48371:48368], addr_12092_7);

wire[31:0] addr_12093_7;

Selector_2 s12093_7(wires_3023_6[1], addr_3023_6, addr_positional[48375:48372], addr_12093_7);

wire[31:0] addr_12094_7;

Selector_2 s12094_7(wires_3023_6[2], addr_3023_6, addr_positional[48379:48376], addr_12094_7);

wire[31:0] addr_12095_7;

Selector_2 s12095_7(wires_3023_6[3], addr_3023_6, addr_positional[48383:48380], addr_12095_7);

wire[31:0] addr_12096_7;

Selector_2 s12096_7(wires_3024_6[0], addr_3024_6, addr_positional[48387:48384], addr_12096_7);

wire[31:0] addr_12097_7;

Selector_2 s12097_7(wires_3024_6[1], addr_3024_6, addr_positional[48391:48388], addr_12097_7);

wire[31:0] addr_12098_7;

Selector_2 s12098_7(wires_3024_6[2], addr_3024_6, addr_positional[48395:48392], addr_12098_7);

wire[31:0] addr_12099_7;

Selector_2 s12099_7(wires_3024_6[3], addr_3024_6, addr_positional[48399:48396], addr_12099_7);

wire[31:0] addr_12100_7;

Selector_2 s12100_7(wires_3025_6[0], addr_3025_6, addr_positional[48403:48400], addr_12100_7);

wire[31:0] addr_12101_7;

Selector_2 s12101_7(wires_3025_6[1], addr_3025_6, addr_positional[48407:48404], addr_12101_7);

wire[31:0] addr_12102_7;

Selector_2 s12102_7(wires_3025_6[2], addr_3025_6, addr_positional[48411:48408], addr_12102_7);

wire[31:0] addr_12103_7;

Selector_2 s12103_7(wires_3025_6[3], addr_3025_6, addr_positional[48415:48412], addr_12103_7);

wire[31:0] addr_12104_7;

Selector_2 s12104_7(wires_3026_6[0], addr_3026_6, addr_positional[48419:48416], addr_12104_7);

wire[31:0] addr_12105_7;

Selector_2 s12105_7(wires_3026_6[1], addr_3026_6, addr_positional[48423:48420], addr_12105_7);

wire[31:0] addr_12106_7;

Selector_2 s12106_7(wires_3026_6[2], addr_3026_6, addr_positional[48427:48424], addr_12106_7);

wire[31:0] addr_12107_7;

Selector_2 s12107_7(wires_3026_6[3], addr_3026_6, addr_positional[48431:48428], addr_12107_7);

wire[31:0] addr_12108_7;

Selector_2 s12108_7(wires_3027_6[0], addr_3027_6, addr_positional[48435:48432], addr_12108_7);

wire[31:0] addr_12109_7;

Selector_2 s12109_7(wires_3027_6[1], addr_3027_6, addr_positional[48439:48436], addr_12109_7);

wire[31:0] addr_12110_7;

Selector_2 s12110_7(wires_3027_6[2], addr_3027_6, addr_positional[48443:48440], addr_12110_7);

wire[31:0] addr_12111_7;

Selector_2 s12111_7(wires_3027_6[3], addr_3027_6, addr_positional[48447:48444], addr_12111_7);

wire[31:0] addr_12112_7;

Selector_2 s12112_7(wires_3028_6[0], addr_3028_6, addr_positional[48451:48448], addr_12112_7);

wire[31:0] addr_12113_7;

Selector_2 s12113_7(wires_3028_6[1], addr_3028_6, addr_positional[48455:48452], addr_12113_7);

wire[31:0] addr_12114_7;

Selector_2 s12114_7(wires_3028_6[2], addr_3028_6, addr_positional[48459:48456], addr_12114_7);

wire[31:0] addr_12115_7;

Selector_2 s12115_7(wires_3028_6[3], addr_3028_6, addr_positional[48463:48460], addr_12115_7);

wire[31:0] addr_12116_7;

Selector_2 s12116_7(wires_3029_6[0], addr_3029_6, addr_positional[48467:48464], addr_12116_7);

wire[31:0] addr_12117_7;

Selector_2 s12117_7(wires_3029_6[1], addr_3029_6, addr_positional[48471:48468], addr_12117_7);

wire[31:0] addr_12118_7;

Selector_2 s12118_7(wires_3029_6[2], addr_3029_6, addr_positional[48475:48472], addr_12118_7);

wire[31:0] addr_12119_7;

Selector_2 s12119_7(wires_3029_6[3], addr_3029_6, addr_positional[48479:48476], addr_12119_7);

wire[31:0] addr_12120_7;

Selector_2 s12120_7(wires_3030_6[0], addr_3030_6, addr_positional[48483:48480], addr_12120_7);

wire[31:0] addr_12121_7;

Selector_2 s12121_7(wires_3030_6[1], addr_3030_6, addr_positional[48487:48484], addr_12121_7);

wire[31:0] addr_12122_7;

Selector_2 s12122_7(wires_3030_6[2], addr_3030_6, addr_positional[48491:48488], addr_12122_7);

wire[31:0] addr_12123_7;

Selector_2 s12123_7(wires_3030_6[3], addr_3030_6, addr_positional[48495:48492], addr_12123_7);

wire[31:0] addr_12124_7;

Selector_2 s12124_7(wires_3031_6[0], addr_3031_6, addr_positional[48499:48496], addr_12124_7);

wire[31:0] addr_12125_7;

Selector_2 s12125_7(wires_3031_6[1], addr_3031_6, addr_positional[48503:48500], addr_12125_7);

wire[31:0] addr_12126_7;

Selector_2 s12126_7(wires_3031_6[2], addr_3031_6, addr_positional[48507:48504], addr_12126_7);

wire[31:0] addr_12127_7;

Selector_2 s12127_7(wires_3031_6[3], addr_3031_6, addr_positional[48511:48508], addr_12127_7);

wire[31:0] addr_12128_7;

Selector_2 s12128_7(wires_3032_6[0], addr_3032_6, addr_positional[48515:48512], addr_12128_7);

wire[31:0] addr_12129_7;

Selector_2 s12129_7(wires_3032_6[1], addr_3032_6, addr_positional[48519:48516], addr_12129_7);

wire[31:0] addr_12130_7;

Selector_2 s12130_7(wires_3032_6[2], addr_3032_6, addr_positional[48523:48520], addr_12130_7);

wire[31:0] addr_12131_7;

Selector_2 s12131_7(wires_3032_6[3], addr_3032_6, addr_positional[48527:48524], addr_12131_7);

wire[31:0] addr_12132_7;

Selector_2 s12132_7(wires_3033_6[0], addr_3033_6, addr_positional[48531:48528], addr_12132_7);

wire[31:0] addr_12133_7;

Selector_2 s12133_7(wires_3033_6[1], addr_3033_6, addr_positional[48535:48532], addr_12133_7);

wire[31:0] addr_12134_7;

Selector_2 s12134_7(wires_3033_6[2], addr_3033_6, addr_positional[48539:48536], addr_12134_7);

wire[31:0] addr_12135_7;

Selector_2 s12135_7(wires_3033_6[3], addr_3033_6, addr_positional[48543:48540], addr_12135_7);

wire[31:0] addr_12136_7;

Selector_2 s12136_7(wires_3034_6[0], addr_3034_6, addr_positional[48547:48544], addr_12136_7);

wire[31:0] addr_12137_7;

Selector_2 s12137_7(wires_3034_6[1], addr_3034_6, addr_positional[48551:48548], addr_12137_7);

wire[31:0] addr_12138_7;

Selector_2 s12138_7(wires_3034_6[2], addr_3034_6, addr_positional[48555:48552], addr_12138_7);

wire[31:0] addr_12139_7;

Selector_2 s12139_7(wires_3034_6[3], addr_3034_6, addr_positional[48559:48556], addr_12139_7);

wire[31:0] addr_12140_7;

Selector_2 s12140_7(wires_3035_6[0], addr_3035_6, addr_positional[48563:48560], addr_12140_7);

wire[31:0] addr_12141_7;

Selector_2 s12141_7(wires_3035_6[1], addr_3035_6, addr_positional[48567:48564], addr_12141_7);

wire[31:0] addr_12142_7;

Selector_2 s12142_7(wires_3035_6[2], addr_3035_6, addr_positional[48571:48568], addr_12142_7);

wire[31:0] addr_12143_7;

Selector_2 s12143_7(wires_3035_6[3], addr_3035_6, addr_positional[48575:48572], addr_12143_7);

wire[31:0] addr_12144_7;

Selector_2 s12144_7(wires_3036_6[0], addr_3036_6, addr_positional[48579:48576], addr_12144_7);

wire[31:0] addr_12145_7;

Selector_2 s12145_7(wires_3036_6[1], addr_3036_6, addr_positional[48583:48580], addr_12145_7);

wire[31:0] addr_12146_7;

Selector_2 s12146_7(wires_3036_6[2], addr_3036_6, addr_positional[48587:48584], addr_12146_7);

wire[31:0] addr_12147_7;

Selector_2 s12147_7(wires_3036_6[3], addr_3036_6, addr_positional[48591:48588], addr_12147_7);

wire[31:0] addr_12148_7;

Selector_2 s12148_7(wires_3037_6[0], addr_3037_6, addr_positional[48595:48592], addr_12148_7);

wire[31:0] addr_12149_7;

Selector_2 s12149_7(wires_3037_6[1], addr_3037_6, addr_positional[48599:48596], addr_12149_7);

wire[31:0] addr_12150_7;

Selector_2 s12150_7(wires_3037_6[2], addr_3037_6, addr_positional[48603:48600], addr_12150_7);

wire[31:0] addr_12151_7;

Selector_2 s12151_7(wires_3037_6[3], addr_3037_6, addr_positional[48607:48604], addr_12151_7);

wire[31:0] addr_12152_7;

Selector_2 s12152_7(wires_3038_6[0], addr_3038_6, addr_positional[48611:48608], addr_12152_7);

wire[31:0] addr_12153_7;

Selector_2 s12153_7(wires_3038_6[1], addr_3038_6, addr_positional[48615:48612], addr_12153_7);

wire[31:0] addr_12154_7;

Selector_2 s12154_7(wires_3038_6[2], addr_3038_6, addr_positional[48619:48616], addr_12154_7);

wire[31:0] addr_12155_7;

Selector_2 s12155_7(wires_3038_6[3], addr_3038_6, addr_positional[48623:48620], addr_12155_7);

wire[31:0] addr_12156_7;

Selector_2 s12156_7(wires_3039_6[0], addr_3039_6, addr_positional[48627:48624], addr_12156_7);

wire[31:0] addr_12157_7;

Selector_2 s12157_7(wires_3039_6[1], addr_3039_6, addr_positional[48631:48628], addr_12157_7);

wire[31:0] addr_12158_7;

Selector_2 s12158_7(wires_3039_6[2], addr_3039_6, addr_positional[48635:48632], addr_12158_7);

wire[31:0] addr_12159_7;

Selector_2 s12159_7(wires_3039_6[3], addr_3039_6, addr_positional[48639:48636], addr_12159_7);

wire[31:0] addr_12160_7;

Selector_2 s12160_7(wires_3040_6[0], addr_3040_6, addr_positional[48643:48640], addr_12160_7);

wire[31:0] addr_12161_7;

Selector_2 s12161_7(wires_3040_6[1], addr_3040_6, addr_positional[48647:48644], addr_12161_7);

wire[31:0] addr_12162_7;

Selector_2 s12162_7(wires_3040_6[2], addr_3040_6, addr_positional[48651:48648], addr_12162_7);

wire[31:0] addr_12163_7;

Selector_2 s12163_7(wires_3040_6[3], addr_3040_6, addr_positional[48655:48652], addr_12163_7);

wire[31:0] addr_12164_7;

Selector_2 s12164_7(wires_3041_6[0], addr_3041_6, addr_positional[48659:48656], addr_12164_7);

wire[31:0] addr_12165_7;

Selector_2 s12165_7(wires_3041_6[1], addr_3041_6, addr_positional[48663:48660], addr_12165_7);

wire[31:0] addr_12166_7;

Selector_2 s12166_7(wires_3041_6[2], addr_3041_6, addr_positional[48667:48664], addr_12166_7);

wire[31:0] addr_12167_7;

Selector_2 s12167_7(wires_3041_6[3], addr_3041_6, addr_positional[48671:48668], addr_12167_7);

wire[31:0] addr_12168_7;

Selector_2 s12168_7(wires_3042_6[0], addr_3042_6, addr_positional[48675:48672], addr_12168_7);

wire[31:0] addr_12169_7;

Selector_2 s12169_7(wires_3042_6[1], addr_3042_6, addr_positional[48679:48676], addr_12169_7);

wire[31:0] addr_12170_7;

Selector_2 s12170_7(wires_3042_6[2], addr_3042_6, addr_positional[48683:48680], addr_12170_7);

wire[31:0] addr_12171_7;

Selector_2 s12171_7(wires_3042_6[3], addr_3042_6, addr_positional[48687:48684], addr_12171_7);

wire[31:0] addr_12172_7;

Selector_2 s12172_7(wires_3043_6[0], addr_3043_6, addr_positional[48691:48688], addr_12172_7);

wire[31:0] addr_12173_7;

Selector_2 s12173_7(wires_3043_6[1], addr_3043_6, addr_positional[48695:48692], addr_12173_7);

wire[31:0] addr_12174_7;

Selector_2 s12174_7(wires_3043_6[2], addr_3043_6, addr_positional[48699:48696], addr_12174_7);

wire[31:0] addr_12175_7;

Selector_2 s12175_7(wires_3043_6[3], addr_3043_6, addr_positional[48703:48700], addr_12175_7);

wire[31:0] addr_12176_7;

Selector_2 s12176_7(wires_3044_6[0], addr_3044_6, addr_positional[48707:48704], addr_12176_7);

wire[31:0] addr_12177_7;

Selector_2 s12177_7(wires_3044_6[1], addr_3044_6, addr_positional[48711:48708], addr_12177_7);

wire[31:0] addr_12178_7;

Selector_2 s12178_7(wires_3044_6[2], addr_3044_6, addr_positional[48715:48712], addr_12178_7);

wire[31:0] addr_12179_7;

Selector_2 s12179_7(wires_3044_6[3], addr_3044_6, addr_positional[48719:48716], addr_12179_7);

wire[31:0] addr_12180_7;

Selector_2 s12180_7(wires_3045_6[0], addr_3045_6, addr_positional[48723:48720], addr_12180_7);

wire[31:0] addr_12181_7;

Selector_2 s12181_7(wires_3045_6[1], addr_3045_6, addr_positional[48727:48724], addr_12181_7);

wire[31:0] addr_12182_7;

Selector_2 s12182_7(wires_3045_6[2], addr_3045_6, addr_positional[48731:48728], addr_12182_7);

wire[31:0] addr_12183_7;

Selector_2 s12183_7(wires_3045_6[3], addr_3045_6, addr_positional[48735:48732], addr_12183_7);

wire[31:0] addr_12184_7;

Selector_2 s12184_7(wires_3046_6[0], addr_3046_6, addr_positional[48739:48736], addr_12184_7);

wire[31:0] addr_12185_7;

Selector_2 s12185_7(wires_3046_6[1], addr_3046_6, addr_positional[48743:48740], addr_12185_7);

wire[31:0] addr_12186_7;

Selector_2 s12186_7(wires_3046_6[2], addr_3046_6, addr_positional[48747:48744], addr_12186_7);

wire[31:0] addr_12187_7;

Selector_2 s12187_7(wires_3046_6[3], addr_3046_6, addr_positional[48751:48748], addr_12187_7);

wire[31:0] addr_12188_7;

Selector_2 s12188_7(wires_3047_6[0], addr_3047_6, addr_positional[48755:48752], addr_12188_7);

wire[31:0] addr_12189_7;

Selector_2 s12189_7(wires_3047_6[1], addr_3047_6, addr_positional[48759:48756], addr_12189_7);

wire[31:0] addr_12190_7;

Selector_2 s12190_7(wires_3047_6[2], addr_3047_6, addr_positional[48763:48760], addr_12190_7);

wire[31:0] addr_12191_7;

Selector_2 s12191_7(wires_3047_6[3], addr_3047_6, addr_positional[48767:48764], addr_12191_7);

wire[31:0] addr_12192_7;

Selector_2 s12192_7(wires_3048_6[0], addr_3048_6, addr_positional[48771:48768], addr_12192_7);

wire[31:0] addr_12193_7;

Selector_2 s12193_7(wires_3048_6[1], addr_3048_6, addr_positional[48775:48772], addr_12193_7);

wire[31:0] addr_12194_7;

Selector_2 s12194_7(wires_3048_6[2], addr_3048_6, addr_positional[48779:48776], addr_12194_7);

wire[31:0] addr_12195_7;

Selector_2 s12195_7(wires_3048_6[3], addr_3048_6, addr_positional[48783:48780], addr_12195_7);

wire[31:0] addr_12196_7;

Selector_2 s12196_7(wires_3049_6[0], addr_3049_6, addr_positional[48787:48784], addr_12196_7);

wire[31:0] addr_12197_7;

Selector_2 s12197_7(wires_3049_6[1], addr_3049_6, addr_positional[48791:48788], addr_12197_7);

wire[31:0] addr_12198_7;

Selector_2 s12198_7(wires_3049_6[2], addr_3049_6, addr_positional[48795:48792], addr_12198_7);

wire[31:0] addr_12199_7;

Selector_2 s12199_7(wires_3049_6[3], addr_3049_6, addr_positional[48799:48796], addr_12199_7);

wire[31:0] addr_12200_7;

Selector_2 s12200_7(wires_3050_6[0], addr_3050_6, addr_positional[48803:48800], addr_12200_7);

wire[31:0] addr_12201_7;

Selector_2 s12201_7(wires_3050_6[1], addr_3050_6, addr_positional[48807:48804], addr_12201_7);

wire[31:0] addr_12202_7;

Selector_2 s12202_7(wires_3050_6[2], addr_3050_6, addr_positional[48811:48808], addr_12202_7);

wire[31:0] addr_12203_7;

Selector_2 s12203_7(wires_3050_6[3], addr_3050_6, addr_positional[48815:48812], addr_12203_7);

wire[31:0] addr_12204_7;

Selector_2 s12204_7(wires_3051_6[0], addr_3051_6, addr_positional[48819:48816], addr_12204_7);

wire[31:0] addr_12205_7;

Selector_2 s12205_7(wires_3051_6[1], addr_3051_6, addr_positional[48823:48820], addr_12205_7);

wire[31:0] addr_12206_7;

Selector_2 s12206_7(wires_3051_6[2], addr_3051_6, addr_positional[48827:48824], addr_12206_7);

wire[31:0] addr_12207_7;

Selector_2 s12207_7(wires_3051_6[3], addr_3051_6, addr_positional[48831:48828], addr_12207_7);

wire[31:0] addr_12208_7;

Selector_2 s12208_7(wires_3052_6[0], addr_3052_6, addr_positional[48835:48832], addr_12208_7);

wire[31:0] addr_12209_7;

Selector_2 s12209_7(wires_3052_6[1], addr_3052_6, addr_positional[48839:48836], addr_12209_7);

wire[31:0] addr_12210_7;

Selector_2 s12210_7(wires_3052_6[2], addr_3052_6, addr_positional[48843:48840], addr_12210_7);

wire[31:0] addr_12211_7;

Selector_2 s12211_7(wires_3052_6[3], addr_3052_6, addr_positional[48847:48844], addr_12211_7);

wire[31:0] addr_12212_7;

Selector_2 s12212_7(wires_3053_6[0], addr_3053_6, addr_positional[48851:48848], addr_12212_7);

wire[31:0] addr_12213_7;

Selector_2 s12213_7(wires_3053_6[1], addr_3053_6, addr_positional[48855:48852], addr_12213_7);

wire[31:0] addr_12214_7;

Selector_2 s12214_7(wires_3053_6[2], addr_3053_6, addr_positional[48859:48856], addr_12214_7);

wire[31:0] addr_12215_7;

Selector_2 s12215_7(wires_3053_6[3], addr_3053_6, addr_positional[48863:48860], addr_12215_7);

wire[31:0] addr_12216_7;

Selector_2 s12216_7(wires_3054_6[0], addr_3054_6, addr_positional[48867:48864], addr_12216_7);

wire[31:0] addr_12217_7;

Selector_2 s12217_7(wires_3054_6[1], addr_3054_6, addr_positional[48871:48868], addr_12217_7);

wire[31:0] addr_12218_7;

Selector_2 s12218_7(wires_3054_6[2], addr_3054_6, addr_positional[48875:48872], addr_12218_7);

wire[31:0] addr_12219_7;

Selector_2 s12219_7(wires_3054_6[3], addr_3054_6, addr_positional[48879:48876], addr_12219_7);

wire[31:0] addr_12220_7;

Selector_2 s12220_7(wires_3055_6[0], addr_3055_6, addr_positional[48883:48880], addr_12220_7);

wire[31:0] addr_12221_7;

Selector_2 s12221_7(wires_3055_6[1], addr_3055_6, addr_positional[48887:48884], addr_12221_7);

wire[31:0] addr_12222_7;

Selector_2 s12222_7(wires_3055_6[2], addr_3055_6, addr_positional[48891:48888], addr_12222_7);

wire[31:0] addr_12223_7;

Selector_2 s12223_7(wires_3055_6[3], addr_3055_6, addr_positional[48895:48892], addr_12223_7);

wire[31:0] addr_12224_7;

Selector_2 s12224_7(wires_3056_6[0], addr_3056_6, addr_positional[48899:48896], addr_12224_7);

wire[31:0] addr_12225_7;

Selector_2 s12225_7(wires_3056_6[1], addr_3056_6, addr_positional[48903:48900], addr_12225_7);

wire[31:0] addr_12226_7;

Selector_2 s12226_7(wires_3056_6[2], addr_3056_6, addr_positional[48907:48904], addr_12226_7);

wire[31:0] addr_12227_7;

Selector_2 s12227_7(wires_3056_6[3], addr_3056_6, addr_positional[48911:48908], addr_12227_7);

wire[31:0] addr_12228_7;

Selector_2 s12228_7(wires_3057_6[0], addr_3057_6, addr_positional[48915:48912], addr_12228_7);

wire[31:0] addr_12229_7;

Selector_2 s12229_7(wires_3057_6[1], addr_3057_6, addr_positional[48919:48916], addr_12229_7);

wire[31:0] addr_12230_7;

Selector_2 s12230_7(wires_3057_6[2], addr_3057_6, addr_positional[48923:48920], addr_12230_7);

wire[31:0] addr_12231_7;

Selector_2 s12231_7(wires_3057_6[3], addr_3057_6, addr_positional[48927:48924], addr_12231_7);

wire[31:0] addr_12232_7;

Selector_2 s12232_7(wires_3058_6[0], addr_3058_6, addr_positional[48931:48928], addr_12232_7);

wire[31:0] addr_12233_7;

Selector_2 s12233_7(wires_3058_6[1], addr_3058_6, addr_positional[48935:48932], addr_12233_7);

wire[31:0] addr_12234_7;

Selector_2 s12234_7(wires_3058_6[2], addr_3058_6, addr_positional[48939:48936], addr_12234_7);

wire[31:0] addr_12235_7;

Selector_2 s12235_7(wires_3058_6[3], addr_3058_6, addr_positional[48943:48940], addr_12235_7);

wire[31:0] addr_12236_7;

Selector_2 s12236_7(wires_3059_6[0], addr_3059_6, addr_positional[48947:48944], addr_12236_7);

wire[31:0] addr_12237_7;

Selector_2 s12237_7(wires_3059_6[1], addr_3059_6, addr_positional[48951:48948], addr_12237_7);

wire[31:0] addr_12238_7;

Selector_2 s12238_7(wires_3059_6[2], addr_3059_6, addr_positional[48955:48952], addr_12238_7);

wire[31:0] addr_12239_7;

Selector_2 s12239_7(wires_3059_6[3], addr_3059_6, addr_positional[48959:48956], addr_12239_7);

wire[31:0] addr_12240_7;

Selector_2 s12240_7(wires_3060_6[0], addr_3060_6, addr_positional[48963:48960], addr_12240_7);

wire[31:0] addr_12241_7;

Selector_2 s12241_7(wires_3060_6[1], addr_3060_6, addr_positional[48967:48964], addr_12241_7);

wire[31:0] addr_12242_7;

Selector_2 s12242_7(wires_3060_6[2], addr_3060_6, addr_positional[48971:48968], addr_12242_7);

wire[31:0] addr_12243_7;

Selector_2 s12243_7(wires_3060_6[3], addr_3060_6, addr_positional[48975:48972], addr_12243_7);

wire[31:0] addr_12244_7;

Selector_2 s12244_7(wires_3061_6[0], addr_3061_6, addr_positional[48979:48976], addr_12244_7);

wire[31:0] addr_12245_7;

Selector_2 s12245_7(wires_3061_6[1], addr_3061_6, addr_positional[48983:48980], addr_12245_7);

wire[31:0] addr_12246_7;

Selector_2 s12246_7(wires_3061_6[2], addr_3061_6, addr_positional[48987:48984], addr_12246_7);

wire[31:0] addr_12247_7;

Selector_2 s12247_7(wires_3061_6[3], addr_3061_6, addr_positional[48991:48988], addr_12247_7);

wire[31:0] addr_12248_7;

Selector_2 s12248_7(wires_3062_6[0], addr_3062_6, addr_positional[48995:48992], addr_12248_7);

wire[31:0] addr_12249_7;

Selector_2 s12249_7(wires_3062_6[1], addr_3062_6, addr_positional[48999:48996], addr_12249_7);

wire[31:0] addr_12250_7;

Selector_2 s12250_7(wires_3062_6[2], addr_3062_6, addr_positional[49003:49000], addr_12250_7);

wire[31:0] addr_12251_7;

Selector_2 s12251_7(wires_3062_6[3], addr_3062_6, addr_positional[49007:49004], addr_12251_7);

wire[31:0] addr_12252_7;

Selector_2 s12252_7(wires_3063_6[0], addr_3063_6, addr_positional[49011:49008], addr_12252_7);

wire[31:0] addr_12253_7;

Selector_2 s12253_7(wires_3063_6[1], addr_3063_6, addr_positional[49015:49012], addr_12253_7);

wire[31:0] addr_12254_7;

Selector_2 s12254_7(wires_3063_6[2], addr_3063_6, addr_positional[49019:49016], addr_12254_7);

wire[31:0] addr_12255_7;

Selector_2 s12255_7(wires_3063_6[3], addr_3063_6, addr_positional[49023:49020], addr_12255_7);

wire[31:0] addr_12256_7;

Selector_2 s12256_7(wires_3064_6[0], addr_3064_6, addr_positional[49027:49024], addr_12256_7);

wire[31:0] addr_12257_7;

Selector_2 s12257_7(wires_3064_6[1], addr_3064_6, addr_positional[49031:49028], addr_12257_7);

wire[31:0] addr_12258_7;

Selector_2 s12258_7(wires_3064_6[2], addr_3064_6, addr_positional[49035:49032], addr_12258_7);

wire[31:0] addr_12259_7;

Selector_2 s12259_7(wires_3064_6[3], addr_3064_6, addr_positional[49039:49036], addr_12259_7);

wire[31:0] addr_12260_7;

Selector_2 s12260_7(wires_3065_6[0], addr_3065_6, addr_positional[49043:49040], addr_12260_7);

wire[31:0] addr_12261_7;

Selector_2 s12261_7(wires_3065_6[1], addr_3065_6, addr_positional[49047:49044], addr_12261_7);

wire[31:0] addr_12262_7;

Selector_2 s12262_7(wires_3065_6[2], addr_3065_6, addr_positional[49051:49048], addr_12262_7);

wire[31:0] addr_12263_7;

Selector_2 s12263_7(wires_3065_6[3], addr_3065_6, addr_positional[49055:49052], addr_12263_7);

wire[31:0] addr_12264_7;

Selector_2 s12264_7(wires_3066_6[0], addr_3066_6, addr_positional[49059:49056], addr_12264_7);

wire[31:0] addr_12265_7;

Selector_2 s12265_7(wires_3066_6[1], addr_3066_6, addr_positional[49063:49060], addr_12265_7);

wire[31:0] addr_12266_7;

Selector_2 s12266_7(wires_3066_6[2], addr_3066_6, addr_positional[49067:49064], addr_12266_7);

wire[31:0] addr_12267_7;

Selector_2 s12267_7(wires_3066_6[3], addr_3066_6, addr_positional[49071:49068], addr_12267_7);

wire[31:0] addr_12268_7;

Selector_2 s12268_7(wires_3067_6[0], addr_3067_6, addr_positional[49075:49072], addr_12268_7);

wire[31:0] addr_12269_7;

Selector_2 s12269_7(wires_3067_6[1], addr_3067_6, addr_positional[49079:49076], addr_12269_7);

wire[31:0] addr_12270_7;

Selector_2 s12270_7(wires_3067_6[2], addr_3067_6, addr_positional[49083:49080], addr_12270_7);

wire[31:0] addr_12271_7;

Selector_2 s12271_7(wires_3067_6[3], addr_3067_6, addr_positional[49087:49084], addr_12271_7);

wire[31:0] addr_12272_7;

Selector_2 s12272_7(wires_3068_6[0], addr_3068_6, addr_positional[49091:49088], addr_12272_7);

wire[31:0] addr_12273_7;

Selector_2 s12273_7(wires_3068_6[1], addr_3068_6, addr_positional[49095:49092], addr_12273_7);

wire[31:0] addr_12274_7;

Selector_2 s12274_7(wires_3068_6[2], addr_3068_6, addr_positional[49099:49096], addr_12274_7);

wire[31:0] addr_12275_7;

Selector_2 s12275_7(wires_3068_6[3], addr_3068_6, addr_positional[49103:49100], addr_12275_7);

wire[31:0] addr_12276_7;

Selector_2 s12276_7(wires_3069_6[0], addr_3069_6, addr_positional[49107:49104], addr_12276_7);

wire[31:0] addr_12277_7;

Selector_2 s12277_7(wires_3069_6[1], addr_3069_6, addr_positional[49111:49108], addr_12277_7);

wire[31:0] addr_12278_7;

Selector_2 s12278_7(wires_3069_6[2], addr_3069_6, addr_positional[49115:49112], addr_12278_7);

wire[31:0] addr_12279_7;

Selector_2 s12279_7(wires_3069_6[3], addr_3069_6, addr_positional[49119:49116], addr_12279_7);

wire[31:0] addr_12280_7;

Selector_2 s12280_7(wires_3070_6[0], addr_3070_6, addr_positional[49123:49120], addr_12280_7);

wire[31:0] addr_12281_7;

Selector_2 s12281_7(wires_3070_6[1], addr_3070_6, addr_positional[49127:49124], addr_12281_7);

wire[31:0] addr_12282_7;

Selector_2 s12282_7(wires_3070_6[2], addr_3070_6, addr_positional[49131:49128], addr_12282_7);

wire[31:0] addr_12283_7;

Selector_2 s12283_7(wires_3070_6[3], addr_3070_6, addr_positional[49135:49132], addr_12283_7);

wire[31:0] addr_12284_7;

Selector_2 s12284_7(wires_3071_6[0], addr_3071_6, addr_positional[49139:49136], addr_12284_7);

wire[31:0] addr_12285_7;

Selector_2 s12285_7(wires_3071_6[1], addr_3071_6, addr_positional[49143:49140], addr_12285_7);

wire[31:0] addr_12286_7;

Selector_2 s12286_7(wires_3071_6[2], addr_3071_6, addr_positional[49147:49144], addr_12286_7);

wire[31:0] addr_12287_7;

Selector_2 s12287_7(wires_3071_6[3], addr_3071_6, addr_positional[49151:49148], addr_12287_7);

wire[31:0] addr_12288_7;

Selector_2 s12288_7(wires_3072_6[0], addr_3072_6, addr_positional[49155:49152], addr_12288_7);

wire[31:0] addr_12289_7;

Selector_2 s12289_7(wires_3072_6[1], addr_3072_6, addr_positional[49159:49156], addr_12289_7);

wire[31:0] addr_12290_7;

Selector_2 s12290_7(wires_3072_6[2], addr_3072_6, addr_positional[49163:49160], addr_12290_7);

wire[31:0] addr_12291_7;

Selector_2 s12291_7(wires_3072_6[3], addr_3072_6, addr_positional[49167:49164], addr_12291_7);

wire[31:0] addr_12292_7;

Selector_2 s12292_7(wires_3073_6[0], addr_3073_6, addr_positional[49171:49168], addr_12292_7);

wire[31:0] addr_12293_7;

Selector_2 s12293_7(wires_3073_6[1], addr_3073_6, addr_positional[49175:49172], addr_12293_7);

wire[31:0] addr_12294_7;

Selector_2 s12294_7(wires_3073_6[2], addr_3073_6, addr_positional[49179:49176], addr_12294_7);

wire[31:0] addr_12295_7;

Selector_2 s12295_7(wires_3073_6[3], addr_3073_6, addr_positional[49183:49180], addr_12295_7);

wire[31:0] addr_12296_7;

Selector_2 s12296_7(wires_3074_6[0], addr_3074_6, addr_positional[49187:49184], addr_12296_7);

wire[31:0] addr_12297_7;

Selector_2 s12297_7(wires_3074_6[1], addr_3074_6, addr_positional[49191:49188], addr_12297_7);

wire[31:0] addr_12298_7;

Selector_2 s12298_7(wires_3074_6[2], addr_3074_6, addr_positional[49195:49192], addr_12298_7);

wire[31:0] addr_12299_7;

Selector_2 s12299_7(wires_3074_6[3], addr_3074_6, addr_positional[49199:49196], addr_12299_7);

wire[31:0] addr_12300_7;

Selector_2 s12300_7(wires_3075_6[0], addr_3075_6, addr_positional[49203:49200], addr_12300_7);

wire[31:0] addr_12301_7;

Selector_2 s12301_7(wires_3075_6[1], addr_3075_6, addr_positional[49207:49204], addr_12301_7);

wire[31:0] addr_12302_7;

Selector_2 s12302_7(wires_3075_6[2], addr_3075_6, addr_positional[49211:49208], addr_12302_7);

wire[31:0] addr_12303_7;

Selector_2 s12303_7(wires_3075_6[3], addr_3075_6, addr_positional[49215:49212], addr_12303_7);

wire[31:0] addr_12304_7;

Selector_2 s12304_7(wires_3076_6[0], addr_3076_6, addr_positional[49219:49216], addr_12304_7);

wire[31:0] addr_12305_7;

Selector_2 s12305_7(wires_3076_6[1], addr_3076_6, addr_positional[49223:49220], addr_12305_7);

wire[31:0] addr_12306_7;

Selector_2 s12306_7(wires_3076_6[2], addr_3076_6, addr_positional[49227:49224], addr_12306_7);

wire[31:0] addr_12307_7;

Selector_2 s12307_7(wires_3076_6[3], addr_3076_6, addr_positional[49231:49228], addr_12307_7);

wire[31:0] addr_12308_7;

Selector_2 s12308_7(wires_3077_6[0], addr_3077_6, addr_positional[49235:49232], addr_12308_7);

wire[31:0] addr_12309_7;

Selector_2 s12309_7(wires_3077_6[1], addr_3077_6, addr_positional[49239:49236], addr_12309_7);

wire[31:0] addr_12310_7;

Selector_2 s12310_7(wires_3077_6[2], addr_3077_6, addr_positional[49243:49240], addr_12310_7);

wire[31:0] addr_12311_7;

Selector_2 s12311_7(wires_3077_6[3], addr_3077_6, addr_positional[49247:49244], addr_12311_7);

wire[31:0] addr_12312_7;

Selector_2 s12312_7(wires_3078_6[0], addr_3078_6, addr_positional[49251:49248], addr_12312_7);

wire[31:0] addr_12313_7;

Selector_2 s12313_7(wires_3078_6[1], addr_3078_6, addr_positional[49255:49252], addr_12313_7);

wire[31:0] addr_12314_7;

Selector_2 s12314_7(wires_3078_6[2], addr_3078_6, addr_positional[49259:49256], addr_12314_7);

wire[31:0] addr_12315_7;

Selector_2 s12315_7(wires_3078_6[3], addr_3078_6, addr_positional[49263:49260], addr_12315_7);

wire[31:0] addr_12316_7;

Selector_2 s12316_7(wires_3079_6[0], addr_3079_6, addr_positional[49267:49264], addr_12316_7);

wire[31:0] addr_12317_7;

Selector_2 s12317_7(wires_3079_6[1], addr_3079_6, addr_positional[49271:49268], addr_12317_7);

wire[31:0] addr_12318_7;

Selector_2 s12318_7(wires_3079_6[2], addr_3079_6, addr_positional[49275:49272], addr_12318_7);

wire[31:0] addr_12319_7;

Selector_2 s12319_7(wires_3079_6[3], addr_3079_6, addr_positional[49279:49276], addr_12319_7);

wire[31:0] addr_12320_7;

Selector_2 s12320_7(wires_3080_6[0], addr_3080_6, addr_positional[49283:49280], addr_12320_7);

wire[31:0] addr_12321_7;

Selector_2 s12321_7(wires_3080_6[1], addr_3080_6, addr_positional[49287:49284], addr_12321_7);

wire[31:0] addr_12322_7;

Selector_2 s12322_7(wires_3080_6[2], addr_3080_6, addr_positional[49291:49288], addr_12322_7);

wire[31:0] addr_12323_7;

Selector_2 s12323_7(wires_3080_6[3], addr_3080_6, addr_positional[49295:49292], addr_12323_7);

wire[31:0] addr_12324_7;

Selector_2 s12324_7(wires_3081_6[0], addr_3081_6, addr_positional[49299:49296], addr_12324_7);

wire[31:0] addr_12325_7;

Selector_2 s12325_7(wires_3081_6[1], addr_3081_6, addr_positional[49303:49300], addr_12325_7);

wire[31:0] addr_12326_7;

Selector_2 s12326_7(wires_3081_6[2], addr_3081_6, addr_positional[49307:49304], addr_12326_7);

wire[31:0] addr_12327_7;

Selector_2 s12327_7(wires_3081_6[3], addr_3081_6, addr_positional[49311:49308], addr_12327_7);

wire[31:0] addr_12328_7;

Selector_2 s12328_7(wires_3082_6[0], addr_3082_6, addr_positional[49315:49312], addr_12328_7);

wire[31:0] addr_12329_7;

Selector_2 s12329_7(wires_3082_6[1], addr_3082_6, addr_positional[49319:49316], addr_12329_7);

wire[31:0] addr_12330_7;

Selector_2 s12330_7(wires_3082_6[2], addr_3082_6, addr_positional[49323:49320], addr_12330_7);

wire[31:0] addr_12331_7;

Selector_2 s12331_7(wires_3082_6[3], addr_3082_6, addr_positional[49327:49324], addr_12331_7);

wire[31:0] addr_12332_7;

Selector_2 s12332_7(wires_3083_6[0], addr_3083_6, addr_positional[49331:49328], addr_12332_7);

wire[31:0] addr_12333_7;

Selector_2 s12333_7(wires_3083_6[1], addr_3083_6, addr_positional[49335:49332], addr_12333_7);

wire[31:0] addr_12334_7;

Selector_2 s12334_7(wires_3083_6[2], addr_3083_6, addr_positional[49339:49336], addr_12334_7);

wire[31:0] addr_12335_7;

Selector_2 s12335_7(wires_3083_6[3], addr_3083_6, addr_positional[49343:49340], addr_12335_7);

wire[31:0] addr_12336_7;

Selector_2 s12336_7(wires_3084_6[0], addr_3084_6, addr_positional[49347:49344], addr_12336_7);

wire[31:0] addr_12337_7;

Selector_2 s12337_7(wires_3084_6[1], addr_3084_6, addr_positional[49351:49348], addr_12337_7);

wire[31:0] addr_12338_7;

Selector_2 s12338_7(wires_3084_6[2], addr_3084_6, addr_positional[49355:49352], addr_12338_7);

wire[31:0] addr_12339_7;

Selector_2 s12339_7(wires_3084_6[3], addr_3084_6, addr_positional[49359:49356], addr_12339_7);

wire[31:0] addr_12340_7;

Selector_2 s12340_7(wires_3085_6[0], addr_3085_6, addr_positional[49363:49360], addr_12340_7);

wire[31:0] addr_12341_7;

Selector_2 s12341_7(wires_3085_6[1], addr_3085_6, addr_positional[49367:49364], addr_12341_7);

wire[31:0] addr_12342_7;

Selector_2 s12342_7(wires_3085_6[2], addr_3085_6, addr_positional[49371:49368], addr_12342_7);

wire[31:0] addr_12343_7;

Selector_2 s12343_7(wires_3085_6[3], addr_3085_6, addr_positional[49375:49372], addr_12343_7);

wire[31:0] addr_12344_7;

Selector_2 s12344_7(wires_3086_6[0], addr_3086_6, addr_positional[49379:49376], addr_12344_7);

wire[31:0] addr_12345_7;

Selector_2 s12345_7(wires_3086_6[1], addr_3086_6, addr_positional[49383:49380], addr_12345_7);

wire[31:0] addr_12346_7;

Selector_2 s12346_7(wires_3086_6[2], addr_3086_6, addr_positional[49387:49384], addr_12346_7);

wire[31:0] addr_12347_7;

Selector_2 s12347_7(wires_3086_6[3], addr_3086_6, addr_positional[49391:49388], addr_12347_7);

wire[31:0] addr_12348_7;

Selector_2 s12348_7(wires_3087_6[0], addr_3087_6, addr_positional[49395:49392], addr_12348_7);

wire[31:0] addr_12349_7;

Selector_2 s12349_7(wires_3087_6[1], addr_3087_6, addr_positional[49399:49396], addr_12349_7);

wire[31:0] addr_12350_7;

Selector_2 s12350_7(wires_3087_6[2], addr_3087_6, addr_positional[49403:49400], addr_12350_7);

wire[31:0] addr_12351_7;

Selector_2 s12351_7(wires_3087_6[3], addr_3087_6, addr_positional[49407:49404], addr_12351_7);

wire[31:0] addr_12352_7;

Selector_2 s12352_7(wires_3088_6[0], addr_3088_6, addr_positional[49411:49408], addr_12352_7);

wire[31:0] addr_12353_7;

Selector_2 s12353_7(wires_3088_6[1], addr_3088_6, addr_positional[49415:49412], addr_12353_7);

wire[31:0] addr_12354_7;

Selector_2 s12354_7(wires_3088_6[2], addr_3088_6, addr_positional[49419:49416], addr_12354_7);

wire[31:0] addr_12355_7;

Selector_2 s12355_7(wires_3088_6[3], addr_3088_6, addr_positional[49423:49420], addr_12355_7);

wire[31:0] addr_12356_7;

Selector_2 s12356_7(wires_3089_6[0], addr_3089_6, addr_positional[49427:49424], addr_12356_7);

wire[31:0] addr_12357_7;

Selector_2 s12357_7(wires_3089_6[1], addr_3089_6, addr_positional[49431:49428], addr_12357_7);

wire[31:0] addr_12358_7;

Selector_2 s12358_7(wires_3089_6[2], addr_3089_6, addr_positional[49435:49432], addr_12358_7);

wire[31:0] addr_12359_7;

Selector_2 s12359_7(wires_3089_6[3], addr_3089_6, addr_positional[49439:49436], addr_12359_7);

wire[31:0] addr_12360_7;

Selector_2 s12360_7(wires_3090_6[0], addr_3090_6, addr_positional[49443:49440], addr_12360_7);

wire[31:0] addr_12361_7;

Selector_2 s12361_7(wires_3090_6[1], addr_3090_6, addr_positional[49447:49444], addr_12361_7);

wire[31:0] addr_12362_7;

Selector_2 s12362_7(wires_3090_6[2], addr_3090_6, addr_positional[49451:49448], addr_12362_7);

wire[31:0] addr_12363_7;

Selector_2 s12363_7(wires_3090_6[3], addr_3090_6, addr_positional[49455:49452], addr_12363_7);

wire[31:0] addr_12364_7;

Selector_2 s12364_7(wires_3091_6[0], addr_3091_6, addr_positional[49459:49456], addr_12364_7);

wire[31:0] addr_12365_7;

Selector_2 s12365_7(wires_3091_6[1], addr_3091_6, addr_positional[49463:49460], addr_12365_7);

wire[31:0] addr_12366_7;

Selector_2 s12366_7(wires_3091_6[2], addr_3091_6, addr_positional[49467:49464], addr_12366_7);

wire[31:0] addr_12367_7;

Selector_2 s12367_7(wires_3091_6[3], addr_3091_6, addr_positional[49471:49468], addr_12367_7);

wire[31:0] addr_12368_7;

Selector_2 s12368_7(wires_3092_6[0], addr_3092_6, addr_positional[49475:49472], addr_12368_7);

wire[31:0] addr_12369_7;

Selector_2 s12369_7(wires_3092_6[1], addr_3092_6, addr_positional[49479:49476], addr_12369_7);

wire[31:0] addr_12370_7;

Selector_2 s12370_7(wires_3092_6[2], addr_3092_6, addr_positional[49483:49480], addr_12370_7);

wire[31:0] addr_12371_7;

Selector_2 s12371_7(wires_3092_6[3], addr_3092_6, addr_positional[49487:49484], addr_12371_7);

wire[31:0] addr_12372_7;

Selector_2 s12372_7(wires_3093_6[0], addr_3093_6, addr_positional[49491:49488], addr_12372_7);

wire[31:0] addr_12373_7;

Selector_2 s12373_7(wires_3093_6[1], addr_3093_6, addr_positional[49495:49492], addr_12373_7);

wire[31:0] addr_12374_7;

Selector_2 s12374_7(wires_3093_6[2], addr_3093_6, addr_positional[49499:49496], addr_12374_7);

wire[31:0] addr_12375_7;

Selector_2 s12375_7(wires_3093_6[3], addr_3093_6, addr_positional[49503:49500], addr_12375_7);

wire[31:0] addr_12376_7;

Selector_2 s12376_7(wires_3094_6[0], addr_3094_6, addr_positional[49507:49504], addr_12376_7);

wire[31:0] addr_12377_7;

Selector_2 s12377_7(wires_3094_6[1], addr_3094_6, addr_positional[49511:49508], addr_12377_7);

wire[31:0] addr_12378_7;

Selector_2 s12378_7(wires_3094_6[2], addr_3094_6, addr_positional[49515:49512], addr_12378_7);

wire[31:0] addr_12379_7;

Selector_2 s12379_7(wires_3094_6[3], addr_3094_6, addr_positional[49519:49516], addr_12379_7);

wire[31:0] addr_12380_7;

Selector_2 s12380_7(wires_3095_6[0], addr_3095_6, addr_positional[49523:49520], addr_12380_7);

wire[31:0] addr_12381_7;

Selector_2 s12381_7(wires_3095_6[1], addr_3095_6, addr_positional[49527:49524], addr_12381_7);

wire[31:0] addr_12382_7;

Selector_2 s12382_7(wires_3095_6[2], addr_3095_6, addr_positional[49531:49528], addr_12382_7);

wire[31:0] addr_12383_7;

Selector_2 s12383_7(wires_3095_6[3], addr_3095_6, addr_positional[49535:49532], addr_12383_7);

wire[31:0] addr_12384_7;

Selector_2 s12384_7(wires_3096_6[0], addr_3096_6, addr_positional[49539:49536], addr_12384_7);

wire[31:0] addr_12385_7;

Selector_2 s12385_7(wires_3096_6[1], addr_3096_6, addr_positional[49543:49540], addr_12385_7);

wire[31:0] addr_12386_7;

Selector_2 s12386_7(wires_3096_6[2], addr_3096_6, addr_positional[49547:49544], addr_12386_7);

wire[31:0] addr_12387_7;

Selector_2 s12387_7(wires_3096_6[3], addr_3096_6, addr_positional[49551:49548], addr_12387_7);

wire[31:0] addr_12388_7;

Selector_2 s12388_7(wires_3097_6[0], addr_3097_6, addr_positional[49555:49552], addr_12388_7);

wire[31:0] addr_12389_7;

Selector_2 s12389_7(wires_3097_6[1], addr_3097_6, addr_positional[49559:49556], addr_12389_7);

wire[31:0] addr_12390_7;

Selector_2 s12390_7(wires_3097_6[2], addr_3097_6, addr_positional[49563:49560], addr_12390_7);

wire[31:0] addr_12391_7;

Selector_2 s12391_7(wires_3097_6[3], addr_3097_6, addr_positional[49567:49564], addr_12391_7);

wire[31:0] addr_12392_7;

Selector_2 s12392_7(wires_3098_6[0], addr_3098_6, addr_positional[49571:49568], addr_12392_7);

wire[31:0] addr_12393_7;

Selector_2 s12393_7(wires_3098_6[1], addr_3098_6, addr_positional[49575:49572], addr_12393_7);

wire[31:0] addr_12394_7;

Selector_2 s12394_7(wires_3098_6[2], addr_3098_6, addr_positional[49579:49576], addr_12394_7);

wire[31:0] addr_12395_7;

Selector_2 s12395_7(wires_3098_6[3], addr_3098_6, addr_positional[49583:49580], addr_12395_7);

wire[31:0] addr_12396_7;

Selector_2 s12396_7(wires_3099_6[0], addr_3099_6, addr_positional[49587:49584], addr_12396_7);

wire[31:0] addr_12397_7;

Selector_2 s12397_7(wires_3099_6[1], addr_3099_6, addr_positional[49591:49588], addr_12397_7);

wire[31:0] addr_12398_7;

Selector_2 s12398_7(wires_3099_6[2], addr_3099_6, addr_positional[49595:49592], addr_12398_7);

wire[31:0] addr_12399_7;

Selector_2 s12399_7(wires_3099_6[3], addr_3099_6, addr_positional[49599:49596], addr_12399_7);

wire[31:0] addr_12400_7;

Selector_2 s12400_7(wires_3100_6[0], addr_3100_6, addr_positional[49603:49600], addr_12400_7);

wire[31:0] addr_12401_7;

Selector_2 s12401_7(wires_3100_6[1], addr_3100_6, addr_positional[49607:49604], addr_12401_7);

wire[31:0] addr_12402_7;

Selector_2 s12402_7(wires_3100_6[2], addr_3100_6, addr_positional[49611:49608], addr_12402_7);

wire[31:0] addr_12403_7;

Selector_2 s12403_7(wires_3100_6[3], addr_3100_6, addr_positional[49615:49612], addr_12403_7);

wire[31:0] addr_12404_7;

Selector_2 s12404_7(wires_3101_6[0], addr_3101_6, addr_positional[49619:49616], addr_12404_7);

wire[31:0] addr_12405_7;

Selector_2 s12405_7(wires_3101_6[1], addr_3101_6, addr_positional[49623:49620], addr_12405_7);

wire[31:0] addr_12406_7;

Selector_2 s12406_7(wires_3101_6[2], addr_3101_6, addr_positional[49627:49624], addr_12406_7);

wire[31:0] addr_12407_7;

Selector_2 s12407_7(wires_3101_6[3], addr_3101_6, addr_positional[49631:49628], addr_12407_7);

wire[31:0] addr_12408_7;

Selector_2 s12408_7(wires_3102_6[0], addr_3102_6, addr_positional[49635:49632], addr_12408_7);

wire[31:0] addr_12409_7;

Selector_2 s12409_7(wires_3102_6[1], addr_3102_6, addr_positional[49639:49636], addr_12409_7);

wire[31:0] addr_12410_7;

Selector_2 s12410_7(wires_3102_6[2], addr_3102_6, addr_positional[49643:49640], addr_12410_7);

wire[31:0] addr_12411_7;

Selector_2 s12411_7(wires_3102_6[3], addr_3102_6, addr_positional[49647:49644], addr_12411_7);

wire[31:0] addr_12412_7;

Selector_2 s12412_7(wires_3103_6[0], addr_3103_6, addr_positional[49651:49648], addr_12412_7);

wire[31:0] addr_12413_7;

Selector_2 s12413_7(wires_3103_6[1], addr_3103_6, addr_positional[49655:49652], addr_12413_7);

wire[31:0] addr_12414_7;

Selector_2 s12414_7(wires_3103_6[2], addr_3103_6, addr_positional[49659:49656], addr_12414_7);

wire[31:0] addr_12415_7;

Selector_2 s12415_7(wires_3103_6[3], addr_3103_6, addr_positional[49663:49660], addr_12415_7);

wire[31:0] addr_12416_7;

Selector_2 s12416_7(wires_3104_6[0], addr_3104_6, addr_positional[49667:49664], addr_12416_7);

wire[31:0] addr_12417_7;

Selector_2 s12417_7(wires_3104_6[1], addr_3104_6, addr_positional[49671:49668], addr_12417_7);

wire[31:0] addr_12418_7;

Selector_2 s12418_7(wires_3104_6[2], addr_3104_6, addr_positional[49675:49672], addr_12418_7);

wire[31:0] addr_12419_7;

Selector_2 s12419_7(wires_3104_6[3], addr_3104_6, addr_positional[49679:49676], addr_12419_7);

wire[31:0] addr_12420_7;

Selector_2 s12420_7(wires_3105_6[0], addr_3105_6, addr_positional[49683:49680], addr_12420_7);

wire[31:0] addr_12421_7;

Selector_2 s12421_7(wires_3105_6[1], addr_3105_6, addr_positional[49687:49684], addr_12421_7);

wire[31:0] addr_12422_7;

Selector_2 s12422_7(wires_3105_6[2], addr_3105_6, addr_positional[49691:49688], addr_12422_7);

wire[31:0] addr_12423_7;

Selector_2 s12423_7(wires_3105_6[3], addr_3105_6, addr_positional[49695:49692], addr_12423_7);

wire[31:0] addr_12424_7;

Selector_2 s12424_7(wires_3106_6[0], addr_3106_6, addr_positional[49699:49696], addr_12424_7);

wire[31:0] addr_12425_7;

Selector_2 s12425_7(wires_3106_6[1], addr_3106_6, addr_positional[49703:49700], addr_12425_7);

wire[31:0] addr_12426_7;

Selector_2 s12426_7(wires_3106_6[2], addr_3106_6, addr_positional[49707:49704], addr_12426_7);

wire[31:0] addr_12427_7;

Selector_2 s12427_7(wires_3106_6[3], addr_3106_6, addr_positional[49711:49708], addr_12427_7);

wire[31:0] addr_12428_7;

Selector_2 s12428_7(wires_3107_6[0], addr_3107_6, addr_positional[49715:49712], addr_12428_7);

wire[31:0] addr_12429_7;

Selector_2 s12429_7(wires_3107_6[1], addr_3107_6, addr_positional[49719:49716], addr_12429_7);

wire[31:0] addr_12430_7;

Selector_2 s12430_7(wires_3107_6[2], addr_3107_6, addr_positional[49723:49720], addr_12430_7);

wire[31:0] addr_12431_7;

Selector_2 s12431_7(wires_3107_6[3], addr_3107_6, addr_positional[49727:49724], addr_12431_7);

wire[31:0] addr_12432_7;

Selector_2 s12432_7(wires_3108_6[0], addr_3108_6, addr_positional[49731:49728], addr_12432_7);

wire[31:0] addr_12433_7;

Selector_2 s12433_7(wires_3108_6[1], addr_3108_6, addr_positional[49735:49732], addr_12433_7);

wire[31:0] addr_12434_7;

Selector_2 s12434_7(wires_3108_6[2], addr_3108_6, addr_positional[49739:49736], addr_12434_7);

wire[31:0] addr_12435_7;

Selector_2 s12435_7(wires_3108_6[3], addr_3108_6, addr_positional[49743:49740], addr_12435_7);

wire[31:0] addr_12436_7;

Selector_2 s12436_7(wires_3109_6[0], addr_3109_6, addr_positional[49747:49744], addr_12436_7);

wire[31:0] addr_12437_7;

Selector_2 s12437_7(wires_3109_6[1], addr_3109_6, addr_positional[49751:49748], addr_12437_7);

wire[31:0] addr_12438_7;

Selector_2 s12438_7(wires_3109_6[2], addr_3109_6, addr_positional[49755:49752], addr_12438_7);

wire[31:0] addr_12439_7;

Selector_2 s12439_7(wires_3109_6[3], addr_3109_6, addr_positional[49759:49756], addr_12439_7);

wire[31:0] addr_12440_7;

Selector_2 s12440_7(wires_3110_6[0], addr_3110_6, addr_positional[49763:49760], addr_12440_7);

wire[31:0] addr_12441_7;

Selector_2 s12441_7(wires_3110_6[1], addr_3110_6, addr_positional[49767:49764], addr_12441_7);

wire[31:0] addr_12442_7;

Selector_2 s12442_7(wires_3110_6[2], addr_3110_6, addr_positional[49771:49768], addr_12442_7);

wire[31:0] addr_12443_7;

Selector_2 s12443_7(wires_3110_6[3], addr_3110_6, addr_positional[49775:49772], addr_12443_7);

wire[31:0] addr_12444_7;

Selector_2 s12444_7(wires_3111_6[0], addr_3111_6, addr_positional[49779:49776], addr_12444_7);

wire[31:0] addr_12445_7;

Selector_2 s12445_7(wires_3111_6[1], addr_3111_6, addr_positional[49783:49780], addr_12445_7);

wire[31:0] addr_12446_7;

Selector_2 s12446_7(wires_3111_6[2], addr_3111_6, addr_positional[49787:49784], addr_12446_7);

wire[31:0] addr_12447_7;

Selector_2 s12447_7(wires_3111_6[3], addr_3111_6, addr_positional[49791:49788], addr_12447_7);

wire[31:0] addr_12448_7;

Selector_2 s12448_7(wires_3112_6[0], addr_3112_6, addr_positional[49795:49792], addr_12448_7);

wire[31:0] addr_12449_7;

Selector_2 s12449_7(wires_3112_6[1], addr_3112_6, addr_positional[49799:49796], addr_12449_7);

wire[31:0] addr_12450_7;

Selector_2 s12450_7(wires_3112_6[2], addr_3112_6, addr_positional[49803:49800], addr_12450_7);

wire[31:0] addr_12451_7;

Selector_2 s12451_7(wires_3112_6[3], addr_3112_6, addr_positional[49807:49804], addr_12451_7);

wire[31:0] addr_12452_7;

Selector_2 s12452_7(wires_3113_6[0], addr_3113_6, addr_positional[49811:49808], addr_12452_7);

wire[31:0] addr_12453_7;

Selector_2 s12453_7(wires_3113_6[1], addr_3113_6, addr_positional[49815:49812], addr_12453_7);

wire[31:0] addr_12454_7;

Selector_2 s12454_7(wires_3113_6[2], addr_3113_6, addr_positional[49819:49816], addr_12454_7);

wire[31:0] addr_12455_7;

Selector_2 s12455_7(wires_3113_6[3], addr_3113_6, addr_positional[49823:49820], addr_12455_7);

wire[31:0] addr_12456_7;

Selector_2 s12456_7(wires_3114_6[0], addr_3114_6, addr_positional[49827:49824], addr_12456_7);

wire[31:0] addr_12457_7;

Selector_2 s12457_7(wires_3114_6[1], addr_3114_6, addr_positional[49831:49828], addr_12457_7);

wire[31:0] addr_12458_7;

Selector_2 s12458_7(wires_3114_6[2], addr_3114_6, addr_positional[49835:49832], addr_12458_7);

wire[31:0] addr_12459_7;

Selector_2 s12459_7(wires_3114_6[3], addr_3114_6, addr_positional[49839:49836], addr_12459_7);

wire[31:0] addr_12460_7;

Selector_2 s12460_7(wires_3115_6[0], addr_3115_6, addr_positional[49843:49840], addr_12460_7);

wire[31:0] addr_12461_7;

Selector_2 s12461_7(wires_3115_6[1], addr_3115_6, addr_positional[49847:49844], addr_12461_7);

wire[31:0] addr_12462_7;

Selector_2 s12462_7(wires_3115_6[2], addr_3115_6, addr_positional[49851:49848], addr_12462_7);

wire[31:0] addr_12463_7;

Selector_2 s12463_7(wires_3115_6[3], addr_3115_6, addr_positional[49855:49852], addr_12463_7);

wire[31:0] addr_12464_7;

Selector_2 s12464_7(wires_3116_6[0], addr_3116_6, addr_positional[49859:49856], addr_12464_7);

wire[31:0] addr_12465_7;

Selector_2 s12465_7(wires_3116_6[1], addr_3116_6, addr_positional[49863:49860], addr_12465_7);

wire[31:0] addr_12466_7;

Selector_2 s12466_7(wires_3116_6[2], addr_3116_6, addr_positional[49867:49864], addr_12466_7);

wire[31:0] addr_12467_7;

Selector_2 s12467_7(wires_3116_6[3], addr_3116_6, addr_positional[49871:49868], addr_12467_7);

wire[31:0] addr_12468_7;

Selector_2 s12468_7(wires_3117_6[0], addr_3117_6, addr_positional[49875:49872], addr_12468_7);

wire[31:0] addr_12469_7;

Selector_2 s12469_7(wires_3117_6[1], addr_3117_6, addr_positional[49879:49876], addr_12469_7);

wire[31:0] addr_12470_7;

Selector_2 s12470_7(wires_3117_6[2], addr_3117_6, addr_positional[49883:49880], addr_12470_7);

wire[31:0] addr_12471_7;

Selector_2 s12471_7(wires_3117_6[3], addr_3117_6, addr_positional[49887:49884], addr_12471_7);

wire[31:0] addr_12472_7;

Selector_2 s12472_7(wires_3118_6[0], addr_3118_6, addr_positional[49891:49888], addr_12472_7);

wire[31:0] addr_12473_7;

Selector_2 s12473_7(wires_3118_6[1], addr_3118_6, addr_positional[49895:49892], addr_12473_7);

wire[31:0] addr_12474_7;

Selector_2 s12474_7(wires_3118_6[2], addr_3118_6, addr_positional[49899:49896], addr_12474_7);

wire[31:0] addr_12475_7;

Selector_2 s12475_7(wires_3118_6[3], addr_3118_6, addr_positional[49903:49900], addr_12475_7);

wire[31:0] addr_12476_7;

Selector_2 s12476_7(wires_3119_6[0], addr_3119_6, addr_positional[49907:49904], addr_12476_7);

wire[31:0] addr_12477_7;

Selector_2 s12477_7(wires_3119_6[1], addr_3119_6, addr_positional[49911:49908], addr_12477_7);

wire[31:0] addr_12478_7;

Selector_2 s12478_7(wires_3119_6[2], addr_3119_6, addr_positional[49915:49912], addr_12478_7);

wire[31:0] addr_12479_7;

Selector_2 s12479_7(wires_3119_6[3], addr_3119_6, addr_positional[49919:49916], addr_12479_7);

wire[31:0] addr_12480_7;

Selector_2 s12480_7(wires_3120_6[0], addr_3120_6, addr_positional[49923:49920], addr_12480_7);

wire[31:0] addr_12481_7;

Selector_2 s12481_7(wires_3120_6[1], addr_3120_6, addr_positional[49927:49924], addr_12481_7);

wire[31:0] addr_12482_7;

Selector_2 s12482_7(wires_3120_6[2], addr_3120_6, addr_positional[49931:49928], addr_12482_7);

wire[31:0] addr_12483_7;

Selector_2 s12483_7(wires_3120_6[3], addr_3120_6, addr_positional[49935:49932], addr_12483_7);

wire[31:0] addr_12484_7;

Selector_2 s12484_7(wires_3121_6[0], addr_3121_6, addr_positional[49939:49936], addr_12484_7);

wire[31:0] addr_12485_7;

Selector_2 s12485_7(wires_3121_6[1], addr_3121_6, addr_positional[49943:49940], addr_12485_7);

wire[31:0] addr_12486_7;

Selector_2 s12486_7(wires_3121_6[2], addr_3121_6, addr_positional[49947:49944], addr_12486_7);

wire[31:0] addr_12487_7;

Selector_2 s12487_7(wires_3121_6[3], addr_3121_6, addr_positional[49951:49948], addr_12487_7);

wire[31:0] addr_12488_7;

Selector_2 s12488_7(wires_3122_6[0], addr_3122_6, addr_positional[49955:49952], addr_12488_7);

wire[31:0] addr_12489_7;

Selector_2 s12489_7(wires_3122_6[1], addr_3122_6, addr_positional[49959:49956], addr_12489_7);

wire[31:0] addr_12490_7;

Selector_2 s12490_7(wires_3122_6[2], addr_3122_6, addr_positional[49963:49960], addr_12490_7);

wire[31:0] addr_12491_7;

Selector_2 s12491_7(wires_3122_6[3], addr_3122_6, addr_positional[49967:49964], addr_12491_7);

wire[31:0] addr_12492_7;

Selector_2 s12492_7(wires_3123_6[0], addr_3123_6, addr_positional[49971:49968], addr_12492_7);

wire[31:0] addr_12493_7;

Selector_2 s12493_7(wires_3123_6[1], addr_3123_6, addr_positional[49975:49972], addr_12493_7);

wire[31:0] addr_12494_7;

Selector_2 s12494_7(wires_3123_6[2], addr_3123_6, addr_positional[49979:49976], addr_12494_7);

wire[31:0] addr_12495_7;

Selector_2 s12495_7(wires_3123_6[3], addr_3123_6, addr_positional[49983:49980], addr_12495_7);

wire[31:0] addr_12496_7;

Selector_2 s12496_7(wires_3124_6[0], addr_3124_6, addr_positional[49987:49984], addr_12496_7);

wire[31:0] addr_12497_7;

Selector_2 s12497_7(wires_3124_6[1], addr_3124_6, addr_positional[49991:49988], addr_12497_7);

wire[31:0] addr_12498_7;

Selector_2 s12498_7(wires_3124_6[2], addr_3124_6, addr_positional[49995:49992], addr_12498_7);

wire[31:0] addr_12499_7;

Selector_2 s12499_7(wires_3124_6[3], addr_3124_6, addr_positional[49999:49996], addr_12499_7);

wire[31:0] addr_12500_7;

Selector_2 s12500_7(wires_3125_6[0], addr_3125_6, addr_positional[50003:50000], addr_12500_7);

wire[31:0] addr_12501_7;

Selector_2 s12501_7(wires_3125_6[1], addr_3125_6, addr_positional[50007:50004], addr_12501_7);

wire[31:0] addr_12502_7;

Selector_2 s12502_7(wires_3125_6[2], addr_3125_6, addr_positional[50011:50008], addr_12502_7);

wire[31:0] addr_12503_7;

Selector_2 s12503_7(wires_3125_6[3], addr_3125_6, addr_positional[50015:50012], addr_12503_7);

wire[31:0] addr_12504_7;

Selector_2 s12504_7(wires_3126_6[0], addr_3126_6, addr_positional[50019:50016], addr_12504_7);

wire[31:0] addr_12505_7;

Selector_2 s12505_7(wires_3126_6[1], addr_3126_6, addr_positional[50023:50020], addr_12505_7);

wire[31:0] addr_12506_7;

Selector_2 s12506_7(wires_3126_6[2], addr_3126_6, addr_positional[50027:50024], addr_12506_7);

wire[31:0] addr_12507_7;

Selector_2 s12507_7(wires_3126_6[3], addr_3126_6, addr_positional[50031:50028], addr_12507_7);

wire[31:0] addr_12508_7;

Selector_2 s12508_7(wires_3127_6[0], addr_3127_6, addr_positional[50035:50032], addr_12508_7);

wire[31:0] addr_12509_7;

Selector_2 s12509_7(wires_3127_6[1], addr_3127_6, addr_positional[50039:50036], addr_12509_7);

wire[31:0] addr_12510_7;

Selector_2 s12510_7(wires_3127_6[2], addr_3127_6, addr_positional[50043:50040], addr_12510_7);

wire[31:0] addr_12511_7;

Selector_2 s12511_7(wires_3127_6[3], addr_3127_6, addr_positional[50047:50044], addr_12511_7);

wire[31:0] addr_12512_7;

Selector_2 s12512_7(wires_3128_6[0], addr_3128_6, addr_positional[50051:50048], addr_12512_7);

wire[31:0] addr_12513_7;

Selector_2 s12513_7(wires_3128_6[1], addr_3128_6, addr_positional[50055:50052], addr_12513_7);

wire[31:0] addr_12514_7;

Selector_2 s12514_7(wires_3128_6[2], addr_3128_6, addr_positional[50059:50056], addr_12514_7);

wire[31:0] addr_12515_7;

Selector_2 s12515_7(wires_3128_6[3], addr_3128_6, addr_positional[50063:50060], addr_12515_7);

wire[31:0] addr_12516_7;

Selector_2 s12516_7(wires_3129_6[0], addr_3129_6, addr_positional[50067:50064], addr_12516_7);

wire[31:0] addr_12517_7;

Selector_2 s12517_7(wires_3129_6[1], addr_3129_6, addr_positional[50071:50068], addr_12517_7);

wire[31:0] addr_12518_7;

Selector_2 s12518_7(wires_3129_6[2], addr_3129_6, addr_positional[50075:50072], addr_12518_7);

wire[31:0] addr_12519_7;

Selector_2 s12519_7(wires_3129_6[3], addr_3129_6, addr_positional[50079:50076], addr_12519_7);

wire[31:0] addr_12520_7;

Selector_2 s12520_7(wires_3130_6[0], addr_3130_6, addr_positional[50083:50080], addr_12520_7);

wire[31:0] addr_12521_7;

Selector_2 s12521_7(wires_3130_6[1], addr_3130_6, addr_positional[50087:50084], addr_12521_7);

wire[31:0] addr_12522_7;

Selector_2 s12522_7(wires_3130_6[2], addr_3130_6, addr_positional[50091:50088], addr_12522_7);

wire[31:0] addr_12523_7;

Selector_2 s12523_7(wires_3130_6[3], addr_3130_6, addr_positional[50095:50092], addr_12523_7);

wire[31:0] addr_12524_7;

Selector_2 s12524_7(wires_3131_6[0], addr_3131_6, addr_positional[50099:50096], addr_12524_7);

wire[31:0] addr_12525_7;

Selector_2 s12525_7(wires_3131_6[1], addr_3131_6, addr_positional[50103:50100], addr_12525_7);

wire[31:0] addr_12526_7;

Selector_2 s12526_7(wires_3131_6[2], addr_3131_6, addr_positional[50107:50104], addr_12526_7);

wire[31:0] addr_12527_7;

Selector_2 s12527_7(wires_3131_6[3], addr_3131_6, addr_positional[50111:50108], addr_12527_7);

wire[31:0] addr_12528_7;

Selector_2 s12528_7(wires_3132_6[0], addr_3132_6, addr_positional[50115:50112], addr_12528_7);

wire[31:0] addr_12529_7;

Selector_2 s12529_7(wires_3132_6[1], addr_3132_6, addr_positional[50119:50116], addr_12529_7);

wire[31:0] addr_12530_7;

Selector_2 s12530_7(wires_3132_6[2], addr_3132_6, addr_positional[50123:50120], addr_12530_7);

wire[31:0] addr_12531_7;

Selector_2 s12531_7(wires_3132_6[3], addr_3132_6, addr_positional[50127:50124], addr_12531_7);

wire[31:0] addr_12532_7;

Selector_2 s12532_7(wires_3133_6[0], addr_3133_6, addr_positional[50131:50128], addr_12532_7);

wire[31:0] addr_12533_7;

Selector_2 s12533_7(wires_3133_6[1], addr_3133_6, addr_positional[50135:50132], addr_12533_7);

wire[31:0] addr_12534_7;

Selector_2 s12534_7(wires_3133_6[2], addr_3133_6, addr_positional[50139:50136], addr_12534_7);

wire[31:0] addr_12535_7;

Selector_2 s12535_7(wires_3133_6[3], addr_3133_6, addr_positional[50143:50140], addr_12535_7);

wire[31:0] addr_12536_7;

Selector_2 s12536_7(wires_3134_6[0], addr_3134_6, addr_positional[50147:50144], addr_12536_7);

wire[31:0] addr_12537_7;

Selector_2 s12537_7(wires_3134_6[1], addr_3134_6, addr_positional[50151:50148], addr_12537_7);

wire[31:0] addr_12538_7;

Selector_2 s12538_7(wires_3134_6[2], addr_3134_6, addr_positional[50155:50152], addr_12538_7);

wire[31:0] addr_12539_7;

Selector_2 s12539_7(wires_3134_6[3], addr_3134_6, addr_positional[50159:50156], addr_12539_7);

wire[31:0] addr_12540_7;

Selector_2 s12540_7(wires_3135_6[0], addr_3135_6, addr_positional[50163:50160], addr_12540_7);

wire[31:0] addr_12541_7;

Selector_2 s12541_7(wires_3135_6[1], addr_3135_6, addr_positional[50167:50164], addr_12541_7);

wire[31:0] addr_12542_7;

Selector_2 s12542_7(wires_3135_6[2], addr_3135_6, addr_positional[50171:50168], addr_12542_7);

wire[31:0] addr_12543_7;

Selector_2 s12543_7(wires_3135_6[3], addr_3135_6, addr_positional[50175:50172], addr_12543_7);

wire[31:0] addr_12544_7;

Selector_2 s12544_7(wires_3136_6[0], addr_3136_6, addr_positional[50179:50176], addr_12544_7);

wire[31:0] addr_12545_7;

Selector_2 s12545_7(wires_3136_6[1], addr_3136_6, addr_positional[50183:50180], addr_12545_7);

wire[31:0] addr_12546_7;

Selector_2 s12546_7(wires_3136_6[2], addr_3136_6, addr_positional[50187:50184], addr_12546_7);

wire[31:0] addr_12547_7;

Selector_2 s12547_7(wires_3136_6[3], addr_3136_6, addr_positional[50191:50188], addr_12547_7);

wire[31:0] addr_12548_7;

Selector_2 s12548_7(wires_3137_6[0], addr_3137_6, addr_positional[50195:50192], addr_12548_7);

wire[31:0] addr_12549_7;

Selector_2 s12549_7(wires_3137_6[1], addr_3137_6, addr_positional[50199:50196], addr_12549_7);

wire[31:0] addr_12550_7;

Selector_2 s12550_7(wires_3137_6[2], addr_3137_6, addr_positional[50203:50200], addr_12550_7);

wire[31:0] addr_12551_7;

Selector_2 s12551_7(wires_3137_6[3], addr_3137_6, addr_positional[50207:50204], addr_12551_7);

wire[31:0] addr_12552_7;

Selector_2 s12552_7(wires_3138_6[0], addr_3138_6, addr_positional[50211:50208], addr_12552_7);

wire[31:0] addr_12553_7;

Selector_2 s12553_7(wires_3138_6[1], addr_3138_6, addr_positional[50215:50212], addr_12553_7);

wire[31:0] addr_12554_7;

Selector_2 s12554_7(wires_3138_6[2], addr_3138_6, addr_positional[50219:50216], addr_12554_7);

wire[31:0] addr_12555_7;

Selector_2 s12555_7(wires_3138_6[3], addr_3138_6, addr_positional[50223:50220], addr_12555_7);

wire[31:0] addr_12556_7;

Selector_2 s12556_7(wires_3139_6[0], addr_3139_6, addr_positional[50227:50224], addr_12556_7);

wire[31:0] addr_12557_7;

Selector_2 s12557_7(wires_3139_6[1], addr_3139_6, addr_positional[50231:50228], addr_12557_7);

wire[31:0] addr_12558_7;

Selector_2 s12558_7(wires_3139_6[2], addr_3139_6, addr_positional[50235:50232], addr_12558_7);

wire[31:0] addr_12559_7;

Selector_2 s12559_7(wires_3139_6[3], addr_3139_6, addr_positional[50239:50236], addr_12559_7);

wire[31:0] addr_12560_7;

Selector_2 s12560_7(wires_3140_6[0], addr_3140_6, addr_positional[50243:50240], addr_12560_7);

wire[31:0] addr_12561_7;

Selector_2 s12561_7(wires_3140_6[1], addr_3140_6, addr_positional[50247:50244], addr_12561_7);

wire[31:0] addr_12562_7;

Selector_2 s12562_7(wires_3140_6[2], addr_3140_6, addr_positional[50251:50248], addr_12562_7);

wire[31:0] addr_12563_7;

Selector_2 s12563_7(wires_3140_6[3], addr_3140_6, addr_positional[50255:50252], addr_12563_7);

wire[31:0] addr_12564_7;

Selector_2 s12564_7(wires_3141_6[0], addr_3141_6, addr_positional[50259:50256], addr_12564_7);

wire[31:0] addr_12565_7;

Selector_2 s12565_7(wires_3141_6[1], addr_3141_6, addr_positional[50263:50260], addr_12565_7);

wire[31:0] addr_12566_7;

Selector_2 s12566_7(wires_3141_6[2], addr_3141_6, addr_positional[50267:50264], addr_12566_7);

wire[31:0] addr_12567_7;

Selector_2 s12567_7(wires_3141_6[3], addr_3141_6, addr_positional[50271:50268], addr_12567_7);

wire[31:0] addr_12568_7;

Selector_2 s12568_7(wires_3142_6[0], addr_3142_6, addr_positional[50275:50272], addr_12568_7);

wire[31:0] addr_12569_7;

Selector_2 s12569_7(wires_3142_6[1], addr_3142_6, addr_positional[50279:50276], addr_12569_7);

wire[31:0] addr_12570_7;

Selector_2 s12570_7(wires_3142_6[2], addr_3142_6, addr_positional[50283:50280], addr_12570_7);

wire[31:0] addr_12571_7;

Selector_2 s12571_7(wires_3142_6[3], addr_3142_6, addr_positional[50287:50284], addr_12571_7);

wire[31:0] addr_12572_7;

Selector_2 s12572_7(wires_3143_6[0], addr_3143_6, addr_positional[50291:50288], addr_12572_7);

wire[31:0] addr_12573_7;

Selector_2 s12573_7(wires_3143_6[1], addr_3143_6, addr_positional[50295:50292], addr_12573_7);

wire[31:0] addr_12574_7;

Selector_2 s12574_7(wires_3143_6[2], addr_3143_6, addr_positional[50299:50296], addr_12574_7);

wire[31:0] addr_12575_7;

Selector_2 s12575_7(wires_3143_6[3], addr_3143_6, addr_positional[50303:50300], addr_12575_7);

wire[31:0] addr_12576_7;

Selector_2 s12576_7(wires_3144_6[0], addr_3144_6, addr_positional[50307:50304], addr_12576_7);

wire[31:0] addr_12577_7;

Selector_2 s12577_7(wires_3144_6[1], addr_3144_6, addr_positional[50311:50308], addr_12577_7);

wire[31:0] addr_12578_7;

Selector_2 s12578_7(wires_3144_6[2], addr_3144_6, addr_positional[50315:50312], addr_12578_7);

wire[31:0] addr_12579_7;

Selector_2 s12579_7(wires_3144_6[3], addr_3144_6, addr_positional[50319:50316], addr_12579_7);

wire[31:0] addr_12580_7;

Selector_2 s12580_7(wires_3145_6[0], addr_3145_6, addr_positional[50323:50320], addr_12580_7);

wire[31:0] addr_12581_7;

Selector_2 s12581_7(wires_3145_6[1], addr_3145_6, addr_positional[50327:50324], addr_12581_7);

wire[31:0] addr_12582_7;

Selector_2 s12582_7(wires_3145_6[2], addr_3145_6, addr_positional[50331:50328], addr_12582_7);

wire[31:0] addr_12583_7;

Selector_2 s12583_7(wires_3145_6[3], addr_3145_6, addr_positional[50335:50332], addr_12583_7);

wire[31:0] addr_12584_7;

Selector_2 s12584_7(wires_3146_6[0], addr_3146_6, addr_positional[50339:50336], addr_12584_7);

wire[31:0] addr_12585_7;

Selector_2 s12585_7(wires_3146_6[1], addr_3146_6, addr_positional[50343:50340], addr_12585_7);

wire[31:0] addr_12586_7;

Selector_2 s12586_7(wires_3146_6[2], addr_3146_6, addr_positional[50347:50344], addr_12586_7);

wire[31:0] addr_12587_7;

Selector_2 s12587_7(wires_3146_6[3], addr_3146_6, addr_positional[50351:50348], addr_12587_7);

wire[31:0] addr_12588_7;

Selector_2 s12588_7(wires_3147_6[0], addr_3147_6, addr_positional[50355:50352], addr_12588_7);

wire[31:0] addr_12589_7;

Selector_2 s12589_7(wires_3147_6[1], addr_3147_6, addr_positional[50359:50356], addr_12589_7);

wire[31:0] addr_12590_7;

Selector_2 s12590_7(wires_3147_6[2], addr_3147_6, addr_positional[50363:50360], addr_12590_7);

wire[31:0] addr_12591_7;

Selector_2 s12591_7(wires_3147_6[3], addr_3147_6, addr_positional[50367:50364], addr_12591_7);

wire[31:0] addr_12592_7;

Selector_2 s12592_7(wires_3148_6[0], addr_3148_6, addr_positional[50371:50368], addr_12592_7);

wire[31:0] addr_12593_7;

Selector_2 s12593_7(wires_3148_6[1], addr_3148_6, addr_positional[50375:50372], addr_12593_7);

wire[31:0] addr_12594_7;

Selector_2 s12594_7(wires_3148_6[2], addr_3148_6, addr_positional[50379:50376], addr_12594_7);

wire[31:0] addr_12595_7;

Selector_2 s12595_7(wires_3148_6[3], addr_3148_6, addr_positional[50383:50380], addr_12595_7);

wire[31:0] addr_12596_7;

Selector_2 s12596_7(wires_3149_6[0], addr_3149_6, addr_positional[50387:50384], addr_12596_7);

wire[31:0] addr_12597_7;

Selector_2 s12597_7(wires_3149_6[1], addr_3149_6, addr_positional[50391:50388], addr_12597_7);

wire[31:0] addr_12598_7;

Selector_2 s12598_7(wires_3149_6[2], addr_3149_6, addr_positional[50395:50392], addr_12598_7);

wire[31:0] addr_12599_7;

Selector_2 s12599_7(wires_3149_6[3], addr_3149_6, addr_positional[50399:50396], addr_12599_7);

wire[31:0] addr_12600_7;

Selector_2 s12600_7(wires_3150_6[0], addr_3150_6, addr_positional[50403:50400], addr_12600_7);

wire[31:0] addr_12601_7;

Selector_2 s12601_7(wires_3150_6[1], addr_3150_6, addr_positional[50407:50404], addr_12601_7);

wire[31:0] addr_12602_7;

Selector_2 s12602_7(wires_3150_6[2], addr_3150_6, addr_positional[50411:50408], addr_12602_7);

wire[31:0] addr_12603_7;

Selector_2 s12603_7(wires_3150_6[3], addr_3150_6, addr_positional[50415:50412], addr_12603_7);

wire[31:0] addr_12604_7;

Selector_2 s12604_7(wires_3151_6[0], addr_3151_6, addr_positional[50419:50416], addr_12604_7);

wire[31:0] addr_12605_7;

Selector_2 s12605_7(wires_3151_6[1], addr_3151_6, addr_positional[50423:50420], addr_12605_7);

wire[31:0] addr_12606_7;

Selector_2 s12606_7(wires_3151_6[2], addr_3151_6, addr_positional[50427:50424], addr_12606_7);

wire[31:0] addr_12607_7;

Selector_2 s12607_7(wires_3151_6[3], addr_3151_6, addr_positional[50431:50428], addr_12607_7);

wire[31:0] addr_12608_7;

Selector_2 s12608_7(wires_3152_6[0], addr_3152_6, addr_positional[50435:50432], addr_12608_7);

wire[31:0] addr_12609_7;

Selector_2 s12609_7(wires_3152_6[1], addr_3152_6, addr_positional[50439:50436], addr_12609_7);

wire[31:0] addr_12610_7;

Selector_2 s12610_7(wires_3152_6[2], addr_3152_6, addr_positional[50443:50440], addr_12610_7);

wire[31:0] addr_12611_7;

Selector_2 s12611_7(wires_3152_6[3], addr_3152_6, addr_positional[50447:50444], addr_12611_7);

wire[31:0] addr_12612_7;

Selector_2 s12612_7(wires_3153_6[0], addr_3153_6, addr_positional[50451:50448], addr_12612_7);

wire[31:0] addr_12613_7;

Selector_2 s12613_7(wires_3153_6[1], addr_3153_6, addr_positional[50455:50452], addr_12613_7);

wire[31:0] addr_12614_7;

Selector_2 s12614_7(wires_3153_6[2], addr_3153_6, addr_positional[50459:50456], addr_12614_7);

wire[31:0] addr_12615_7;

Selector_2 s12615_7(wires_3153_6[3], addr_3153_6, addr_positional[50463:50460], addr_12615_7);

wire[31:0] addr_12616_7;

Selector_2 s12616_7(wires_3154_6[0], addr_3154_6, addr_positional[50467:50464], addr_12616_7);

wire[31:0] addr_12617_7;

Selector_2 s12617_7(wires_3154_6[1], addr_3154_6, addr_positional[50471:50468], addr_12617_7);

wire[31:0] addr_12618_7;

Selector_2 s12618_7(wires_3154_6[2], addr_3154_6, addr_positional[50475:50472], addr_12618_7);

wire[31:0] addr_12619_7;

Selector_2 s12619_7(wires_3154_6[3], addr_3154_6, addr_positional[50479:50476], addr_12619_7);

wire[31:0] addr_12620_7;

Selector_2 s12620_7(wires_3155_6[0], addr_3155_6, addr_positional[50483:50480], addr_12620_7);

wire[31:0] addr_12621_7;

Selector_2 s12621_7(wires_3155_6[1], addr_3155_6, addr_positional[50487:50484], addr_12621_7);

wire[31:0] addr_12622_7;

Selector_2 s12622_7(wires_3155_6[2], addr_3155_6, addr_positional[50491:50488], addr_12622_7);

wire[31:0] addr_12623_7;

Selector_2 s12623_7(wires_3155_6[3], addr_3155_6, addr_positional[50495:50492], addr_12623_7);

wire[31:0] addr_12624_7;

Selector_2 s12624_7(wires_3156_6[0], addr_3156_6, addr_positional[50499:50496], addr_12624_7);

wire[31:0] addr_12625_7;

Selector_2 s12625_7(wires_3156_6[1], addr_3156_6, addr_positional[50503:50500], addr_12625_7);

wire[31:0] addr_12626_7;

Selector_2 s12626_7(wires_3156_6[2], addr_3156_6, addr_positional[50507:50504], addr_12626_7);

wire[31:0] addr_12627_7;

Selector_2 s12627_7(wires_3156_6[3], addr_3156_6, addr_positional[50511:50508], addr_12627_7);

wire[31:0] addr_12628_7;

Selector_2 s12628_7(wires_3157_6[0], addr_3157_6, addr_positional[50515:50512], addr_12628_7);

wire[31:0] addr_12629_7;

Selector_2 s12629_7(wires_3157_6[1], addr_3157_6, addr_positional[50519:50516], addr_12629_7);

wire[31:0] addr_12630_7;

Selector_2 s12630_7(wires_3157_6[2], addr_3157_6, addr_positional[50523:50520], addr_12630_7);

wire[31:0] addr_12631_7;

Selector_2 s12631_7(wires_3157_6[3], addr_3157_6, addr_positional[50527:50524], addr_12631_7);

wire[31:0] addr_12632_7;

Selector_2 s12632_7(wires_3158_6[0], addr_3158_6, addr_positional[50531:50528], addr_12632_7);

wire[31:0] addr_12633_7;

Selector_2 s12633_7(wires_3158_6[1], addr_3158_6, addr_positional[50535:50532], addr_12633_7);

wire[31:0] addr_12634_7;

Selector_2 s12634_7(wires_3158_6[2], addr_3158_6, addr_positional[50539:50536], addr_12634_7);

wire[31:0] addr_12635_7;

Selector_2 s12635_7(wires_3158_6[3], addr_3158_6, addr_positional[50543:50540], addr_12635_7);

wire[31:0] addr_12636_7;

Selector_2 s12636_7(wires_3159_6[0], addr_3159_6, addr_positional[50547:50544], addr_12636_7);

wire[31:0] addr_12637_7;

Selector_2 s12637_7(wires_3159_6[1], addr_3159_6, addr_positional[50551:50548], addr_12637_7);

wire[31:0] addr_12638_7;

Selector_2 s12638_7(wires_3159_6[2], addr_3159_6, addr_positional[50555:50552], addr_12638_7);

wire[31:0] addr_12639_7;

Selector_2 s12639_7(wires_3159_6[3], addr_3159_6, addr_positional[50559:50556], addr_12639_7);

wire[31:0] addr_12640_7;

Selector_2 s12640_7(wires_3160_6[0], addr_3160_6, addr_positional[50563:50560], addr_12640_7);

wire[31:0] addr_12641_7;

Selector_2 s12641_7(wires_3160_6[1], addr_3160_6, addr_positional[50567:50564], addr_12641_7);

wire[31:0] addr_12642_7;

Selector_2 s12642_7(wires_3160_6[2], addr_3160_6, addr_positional[50571:50568], addr_12642_7);

wire[31:0] addr_12643_7;

Selector_2 s12643_7(wires_3160_6[3], addr_3160_6, addr_positional[50575:50572], addr_12643_7);

wire[31:0] addr_12644_7;

Selector_2 s12644_7(wires_3161_6[0], addr_3161_6, addr_positional[50579:50576], addr_12644_7);

wire[31:0] addr_12645_7;

Selector_2 s12645_7(wires_3161_6[1], addr_3161_6, addr_positional[50583:50580], addr_12645_7);

wire[31:0] addr_12646_7;

Selector_2 s12646_7(wires_3161_6[2], addr_3161_6, addr_positional[50587:50584], addr_12646_7);

wire[31:0] addr_12647_7;

Selector_2 s12647_7(wires_3161_6[3], addr_3161_6, addr_positional[50591:50588], addr_12647_7);

wire[31:0] addr_12648_7;

Selector_2 s12648_7(wires_3162_6[0], addr_3162_6, addr_positional[50595:50592], addr_12648_7);

wire[31:0] addr_12649_7;

Selector_2 s12649_7(wires_3162_6[1], addr_3162_6, addr_positional[50599:50596], addr_12649_7);

wire[31:0] addr_12650_7;

Selector_2 s12650_7(wires_3162_6[2], addr_3162_6, addr_positional[50603:50600], addr_12650_7);

wire[31:0] addr_12651_7;

Selector_2 s12651_7(wires_3162_6[3], addr_3162_6, addr_positional[50607:50604], addr_12651_7);

wire[31:0] addr_12652_7;

Selector_2 s12652_7(wires_3163_6[0], addr_3163_6, addr_positional[50611:50608], addr_12652_7);

wire[31:0] addr_12653_7;

Selector_2 s12653_7(wires_3163_6[1], addr_3163_6, addr_positional[50615:50612], addr_12653_7);

wire[31:0] addr_12654_7;

Selector_2 s12654_7(wires_3163_6[2], addr_3163_6, addr_positional[50619:50616], addr_12654_7);

wire[31:0] addr_12655_7;

Selector_2 s12655_7(wires_3163_6[3], addr_3163_6, addr_positional[50623:50620], addr_12655_7);

wire[31:0] addr_12656_7;

Selector_2 s12656_7(wires_3164_6[0], addr_3164_6, addr_positional[50627:50624], addr_12656_7);

wire[31:0] addr_12657_7;

Selector_2 s12657_7(wires_3164_6[1], addr_3164_6, addr_positional[50631:50628], addr_12657_7);

wire[31:0] addr_12658_7;

Selector_2 s12658_7(wires_3164_6[2], addr_3164_6, addr_positional[50635:50632], addr_12658_7);

wire[31:0] addr_12659_7;

Selector_2 s12659_7(wires_3164_6[3], addr_3164_6, addr_positional[50639:50636], addr_12659_7);

wire[31:0] addr_12660_7;

Selector_2 s12660_7(wires_3165_6[0], addr_3165_6, addr_positional[50643:50640], addr_12660_7);

wire[31:0] addr_12661_7;

Selector_2 s12661_7(wires_3165_6[1], addr_3165_6, addr_positional[50647:50644], addr_12661_7);

wire[31:0] addr_12662_7;

Selector_2 s12662_7(wires_3165_6[2], addr_3165_6, addr_positional[50651:50648], addr_12662_7);

wire[31:0] addr_12663_7;

Selector_2 s12663_7(wires_3165_6[3], addr_3165_6, addr_positional[50655:50652], addr_12663_7);

wire[31:0] addr_12664_7;

Selector_2 s12664_7(wires_3166_6[0], addr_3166_6, addr_positional[50659:50656], addr_12664_7);

wire[31:0] addr_12665_7;

Selector_2 s12665_7(wires_3166_6[1], addr_3166_6, addr_positional[50663:50660], addr_12665_7);

wire[31:0] addr_12666_7;

Selector_2 s12666_7(wires_3166_6[2], addr_3166_6, addr_positional[50667:50664], addr_12666_7);

wire[31:0] addr_12667_7;

Selector_2 s12667_7(wires_3166_6[3], addr_3166_6, addr_positional[50671:50668], addr_12667_7);

wire[31:0] addr_12668_7;

Selector_2 s12668_7(wires_3167_6[0], addr_3167_6, addr_positional[50675:50672], addr_12668_7);

wire[31:0] addr_12669_7;

Selector_2 s12669_7(wires_3167_6[1], addr_3167_6, addr_positional[50679:50676], addr_12669_7);

wire[31:0] addr_12670_7;

Selector_2 s12670_7(wires_3167_6[2], addr_3167_6, addr_positional[50683:50680], addr_12670_7);

wire[31:0] addr_12671_7;

Selector_2 s12671_7(wires_3167_6[3], addr_3167_6, addr_positional[50687:50684], addr_12671_7);

wire[31:0] addr_12672_7;

Selector_2 s12672_7(wires_3168_6[0], addr_3168_6, addr_positional[50691:50688], addr_12672_7);

wire[31:0] addr_12673_7;

Selector_2 s12673_7(wires_3168_6[1], addr_3168_6, addr_positional[50695:50692], addr_12673_7);

wire[31:0] addr_12674_7;

Selector_2 s12674_7(wires_3168_6[2], addr_3168_6, addr_positional[50699:50696], addr_12674_7);

wire[31:0] addr_12675_7;

Selector_2 s12675_7(wires_3168_6[3], addr_3168_6, addr_positional[50703:50700], addr_12675_7);

wire[31:0] addr_12676_7;

Selector_2 s12676_7(wires_3169_6[0], addr_3169_6, addr_positional[50707:50704], addr_12676_7);

wire[31:0] addr_12677_7;

Selector_2 s12677_7(wires_3169_6[1], addr_3169_6, addr_positional[50711:50708], addr_12677_7);

wire[31:0] addr_12678_7;

Selector_2 s12678_7(wires_3169_6[2], addr_3169_6, addr_positional[50715:50712], addr_12678_7);

wire[31:0] addr_12679_7;

Selector_2 s12679_7(wires_3169_6[3], addr_3169_6, addr_positional[50719:50716], addr_12679_7);

wire[31:0] addr_12680_7;

Selector_2 s12680_7(wires_3170_6[0], addr_3170_6, addr_positional[50723:50720], addr_12680_7);

wire[31:0] addr_12681_7;

Selector_2 s12681_7(wires_3170_6[1], addr_3170_6, addr_positional[50727:50724], addr_12681_7);

wire[31:0] addr_12682_7;

Selector_2 s12682_7(wires_3170_6[2], addr_3170_6, addr_positional[50731:50728], addr_12682_7);

wire[31:0] addr_12683_7;

Selector_2 s12683_7(wires_3170_6[3], addr_3170_6, addr_positional[50735:50732], addr_12683_7);

wire[31:0] addr_12684_7;

Selector_2 s12684_7(wires_3171_6[0], addr_3171_6, addr_positional[50739:50736], addr_12684_7);

wire[31:0] addr_12685_7;

Selector_2 s12685_7(wires_3171_6[1], addr_3171_6, addr_positional[50743:50740], addr_12685_7);

wire[31:0] addr_12686_7;

Selector_2 s12686_7(wires_3171_6[2], addr_3171_6, addr_positional[50747:50744], addr_12686_7);

wire[31:0] addr_12687_7;

Selector_2 s12687_7(wires_3171_6[3], addr_3171_6, addr_positional[50751:50748], addr_12687_7);

wire[31:0] addr_12688_7;

Selector_2 s12688_7(wires_3172_6[0], addr_3172_6, addr_positional[50755:50752], addr_12688_7);

wire[31:0] addr_12689_7;

Selector_2 s12689_7(wires_3172_6[1], addr_3172_6, addr_positional[50759:50756], addr_12689_7);

wire[31:0] addr_12690_7;

Selector_2 s12690_7(wires_3172_6[2], addr_3172_6, addr_positional[50763:50760], addr_12690_7);

wire[31:0] addr_12691_7;

Selector_2 s12691_7(wires_3172_6[3], addr_3172_6, addr_positional[50767:50764], addr_12691_7);

wire[31:0] addr_12692_7;

Selector_2 s12692_7(wires_3173_6[0], addr_3173_6, addr_positional[50771:50768], addr_12692_7);

wire[31:0] addr_12693_7;

Selector_2 s12693_7(wires_3173_6[1], addr_3173_6, addr_positional[50775:50772], addr_12693_7);

wire[31:0] addr_12694_7;

Selector_2 s12694_7(wires_3173_6[2], addr_3173_6, addr_positional[50779:50776], addr_12694_7);

wire[31:0] addr_12695_7;

Selector_2 s12695_7(wires_3173_6[3], addr_3173_6, addr_positional[50783:50780], addr_12695_7);

wire[31:0] addr_12696_7;

Selector_2 s12696_7(wires_3174_6[0], addr_3174_6, addr_positional[50787:50784], addr_12696_7);

wire[31:0] addr_12697_7;

Selector_2 s12697_7(wires_3174_6[1], addr_3174_6, addr_positional[50791:50788], addr_12697_7);

wire[31:0] addr_12698_7;

Selector_2 s12698_7(wires_3174_6[2], addr_3174_6, addr_positional[50795:50792], addr_12698_7);

wire[31:0] addr_12699_7;

Selector_2 s12699_7(wires_3174_6[3], addr_3174_6, addr_positional[50799:50796], addr_12699_7);

wire[31:0] addr_12700_7;

Selector_2 s12700_7(wires_3175_6[0], addr_3175_6, addr_positional[50803:50800], addr_12700_7);

wire[31:0] addr_12701_7;

Selector_2 s12701_7(wires_3175_6[1], addr_3175_6, addr_positional[50807:50804], addr_12701_7);

wire[31:0] addr_12702_7;

Selector_2 s12702_7(wires_3175_6[2], addr_3175_6, addr_positional[50811:50808], addr_12702_7);

wire[31:0] addr_12703_7;

Selector_2 s12703_7(wires_3175_6[3], addr_3175_6, addr_positional[50815:50812], addr_12703_7);

wire[31:0] addr_12704_7;

Selector_2 s12704_7(wires_3176_6[0], addr_3176_6, addr_positional[50819:50816], addr_12704_7);

wire[31:0] addr_12705_7;

Selector_2 s12705_7(wires_3176_6[1], addr_3176_6, addr_positional[50823:50820], addr_12705_7);

wire[31:0] addr_12706_7;

Selector_2 s12706_7(wires_3176_6[2], addr_3176_6, addr_positional[50827:50824], addr_12706_7);

wire[31:0] addr_12707_7;

Selector_2 s12707_7(wires_3176_6[3], addr_3176_6, addr_positional[50831:50828], addr_12707_7);

wire[31:0] addr_12708_7;

Selector_2 s12708_7(wires_3177_6[0], addr_3177_6, addr_positional[50835:50832], addr_12708_7);

wire[31:0] addr_12709_7;

Selector_2 s12709_7(wires_3177_6[1], addr_3177_6, addr_positional[50839:50836], addr_12709_7);

wire[31:0] addr_12710_7;

Selector_2 s12710_7(wires_3177_6[2], addr_3177_6, addr_positional[50843:50840], addr_12710_7);

wire[31:0] addr_12711_7;

Selector_2 s12711_7(wires_3177_6[3], addr_3177_6, addr_positional[50847:50844], addr_12711_7);

wire[31:0] addr_12712_7;

Selector_2 s12712_7(wires_3178_6[0], addr_3178_6, addr_positional[50851:50848], addr_12712_7);

wire[31:0] addr_12713_7;

Selector_2 s12713_7(wires_3178_6[1], addr_3178_6, addr_positional[50855:50852], addr_12713_7);

wire[31:0] addr_12714_7;

Selector_2 s12714_7(wires_3178_6[2], addr_3178_6, addr_positional[50859:50856], addr_12714_7);

wire[31:0] addr_12715_7;

Selector_2 s12715_7(wires_3178_6[3], addr_3178_6, addr_positional[50863:50860], addr_12715_7);

wire[31:0] addr_12716_7;

Selector_2 s12716_7(wires_3179_6[0], addr_3179_6, addr_positional[50867:50864], addr_12716_7);

wire[31:0] addr_12717_7;

Selector_2 s12717_7(wires_3179_6[1], addr_3179_6, addr_positional[50871:50868], addr_12717_7);

wire[31:0] addr_12718_7;

Selector_2 s12718_7(wires_3179_6[2], addr_3179_6, addr_positional[50875:50872], addr_12718_7);

wire[31:0] addr_12719_7;

Selector_2 s12719_7(wires_3179_6[3], addr_3179_6, addr_positional[50879:50876], addr_12719_7);

wire[31:0] addr_12720_7;

Selector_2 s12720_7(wires_3180_6[0], addr_3180_6, addr_positional[50883:50880], addr_12720_7);

wire[31:0] addr_12721_7;

Selector_2 s12721_7(wires_3180_6[1], addr_3180_6, addr_positional[50887:50884], addr_12721_7);

wire[31:0] addr_12722_7;

Selector_2 s12722_7(wires_3180_6[2], addr_3180_6, addr_positional[50891:50888], addr_12722_7);

wire[31:0] addr_12723_7;

Selector_2 s12723_7(wires_3180_6[3], addr_3180_6, addr_positional[50895:50892], addr_12723_7);

wire[31:0] addr_12724_7;

Selector_2 s12724_7(wires_3181_6[0], addr_3181_6, addr_positional[50899:50896], addr_12724_7);

wire[31:0] addr_12725_7;

Selector_2 s12725_7(wires_3181_6[1], addr_3181_6, addr_positional[50903:50900], addr_12725_7);

wire[31:0] addr_12726_7;

Selector_2 s12726_7(wires_3181_6[2], addr_3181_6, addr_positional[50907:50904], addr_12726_7);

wire[31:0] addr_12727_7;

Selector_2 s12727_7(wires_3181_6[3], addr_3181_6, addr_positional[50911:50908], addr_12727_7);

wire[31:0] addr_12728_7;

Selector_2 s12728_7(wires_3182_6[0], addr_3182_6, addr_positional[50915:50912], addr_12728_7);

wire[31:0] addr_12729_7;

Selector_2 s12729_7(wires_3182_6[1], addr_3182_6, addr_positional[50919:50916], addr_12729_7);

wire[31:0] addr_12730_7;

Selector_2 s12730_7(wires_3182_6[2], addr_3182_6, addr_positional[50923:50920], addr_12730_7);

wire[31:0] addr_12731_7;

Selector_2 s12731_7(wires_3182_6[3], addr_3182_6, addr_positional[50927:50924], addr_12731_7);

wire[31:0] addr_12732_7;

Selector_2 s12732_7(wires_3183_6[0], addr_3183_6, addr_positional[50931:50928], addr_12732_7);

wire[31:0] addr_12733_7;

Selector_2 s12733_7(wires_3183_6[1], addr_3183_6, addr_positional[50935:50932], addr_12733_7);

wire[31:0] addr_12734_7;

Selector_2 s12734_7(wires_3183_6[2], addr_3183_6, addr_positional[50939:50936], addr_12734_7);

wire[31:0] addr_12735_7;

Selector_2 s12735_7(wires_3183_6[3], addr_3183_6, addr_positional[50943:50940], addr_12735_7);

wire[31:0] addr_12736_7;

Selector_2 s12736_7(wires_3184_6[0], addr_3184_6, addr_positional[50947:50944], addr_12736_7);

wire[31:0] addr_12737_7;

Selector_2 s12737_7(wires_3184_6[1], addr_3184_6, addr_positional[50951:50948], addr_12737_7);

wire[31:0] addr_12738_7;

Selector_2 s12738_7(wires_3184_6[2], addr_3184_6, addr_positional[50955:50952], addr_12738_7);

wire[31:0] addr_12739_7;

Selector_2 s12739_7(wires_3184_6[3], addr_3184_6, addr_positional[50959:50956], addr_12739_7);

wire[31:0] addr_12740_7;

Selector_2 s12740_7(wires_3185_6[0], addr_3185_6, addr_positional[50963:50960], addr_12740_7);

wire[31:0] addr_12741_7;

Selector_2 s12741_7(wires_3185_6[1], addr_3185_6, addr_positional[50967:50964], addr_12741_7);

wire[31:0] addr_12742_7;

Selector_2 s12742_7(wires_3185_6[2], addr_3185_6, addr_positional[50971:50968], addr_12742_7);

wire[31:0] addr_12743_7;

Selector_2 s12743_7(wires_3185_6[3], addr_3185_6, addr_positional[50975:50972], addr_12743_7);

wire[31:0] addr_12744_7;

Selector_2 s12744_7(wires_3186_6[0], addr_3186_6, addr_positional[50979:50976], addr_12744_7);

wire[31:0] addr_12745_7;

Selector_2 s12745_7(wires_3186_6[1], addr_3186_6, addr_positional[50983:50980], addr_12745_7);

wire[31:0] addr_12746_7;

Selector_2 s12746_7(wires_3186_6[2], addr_3186_6, addr_positional[50987:50984], addr_12746_7);

wire[31:0] addr_12747_7;

Selector_2 s12747_7(wires_3186_6[3], addr_3186_6, addr_positional[50991:50988], addr_12747_7);

wire[31:0] addr_12748_7;

Selector_2 s12748_7(wires_3187_6[0], addr_3187_6, addr_positional[50995:50992], addr_12748_7);

wire[31:0] addr_12749_7;

Selector_2 s12749_7(wires_3187_6[1], addr_3187_6, addr_positional[50999:50996], addr_12749_7);

wire[31:0] addr_12750_7;

Selector_2 s12750_7(wires_3187_6[2], addr_3187_6, addr_positional[51003:51000], addr_12750_7);

wire[31:0] addr_12751_7;

Selector_2 s12751_7(wires_3187_6[3], addr_3187_6, addr_positional[51007:51004], addr_12751_7);

wire[31:0] addr_12752_7;

Selector_2 s12752_7(wires_3188_6[0], addr_3188_6, addr_positional[51011:51008], addr_12752_7);

wire[31:0] addr_12753_7;

Selector_2 s12753_7(wires_3188_6[1], addr_3188_6, addr_positional[51015:51012], addr_12753_7);

wire[31:0] addr_12754_7;

Selector_2 s12754_7(wires_3188_6[2], addr_3188_6, addr_positional[51019:51016], addr_12754_7);

wire[31:0] addr_12755_7;

Selector_2 s12755_7(wires_3188_6[3], addr_3188_6, addr_positional[51023:51020], addr_12755_7);

wire[31:0] addr_12756_7;

Selector_2 s12756_7(wires_3189_6[0], addr_3189_6, addr_positional[51027:51024], addr_12756_7);

wire[31:0] addr_12757_7;

Selector_2 s12757_7(wires_3189_6[1], addr_3189_6, addr_positional[51031:51028], addr_12757_7);

wire[31:0] addr_12758_7;

Selector_2 s12758_7(wires_3189_6[2], addr_3189_6, addr_positional[51035:51032], addr_12758_7);

wire[31:0] addr_12759_7;

Selector_2 s12759_7(wires_3189_6[3], addr_3189_6, addr_positional[51039:51036], addr_12759_7);

wire[31:0] addr_12760_7;

Selector_2 s12760_7(wires_3190_6[0], addr_3190_6, addr_positional[51043:51040], addr_12760_7);

wire[31:0] addr_12761_7;

Selector_2 s12761_7(wires_3190_6[1], addr_3190_6, addr_positional[51047:51044], addr_12761_7);

wire[31:0] addr_12762_7;

Selector_2 s12762_7(wires_3190_6[2], addr_3190_6, addr_positional[51051:51048], addr_12762_7);

wire[31:0] addr_12763_7;

Selector_2 s12763_7(wires_3190_6[3], addr_3190_6, addr_positional[51055:51052], addr_12763_7);

wire[31:0] addr_12764_7;

Selector_2 s12764_7(wires_3191_6[0], addr_3191_6, addr_positional[51059:51056], addr_12764_7);

wire[31:0] addr_12765_7;

Selector_2 s12765_7(wires_3191_6[1], addr_3191_6, addr_positional[51063:51060], addr_12765_7);

wire[31:0] addr_12766_7;

Selector_2 s12766_7(wires_3191_6[2], addr_3191_6, addr_positional[51067:51064], addr_12766_7);

wire[31:0] addr_12767_7;

Selector_2 s12767_7(wires_3191_6[3], addr_3191_6, addr_positional[51071:51068], addr_12767_7);

wire[31:0] addr_12768_7;

Selector_2 s12768_7(wires_3192_6[0], addr_3192_6, addr_positional[51075:51072], addr_12768_7);

wire[31:0] addr_12769_7;

Selector_2 s12769_7(wires_3192_6[1], addr_3192_6, addr_positional[51079:51076], addr_12769_7);

wire[31:0] addr_12770_7;

Selector_2 s12770_7(wires_3192_6[2], addr_3192_6, addr_positional[51083:51080], addr_12770_7);

wire[31:0] addr_12771_7;

Selector_2 s12771_7(wires_3192_6[3], addr_3192_6, addr_positional[51087:51084], addr_12771_7);

wire[31:0] addr_12772_7;

Selector_2 s12772_7(wires_3193_6[0], addr_3193_6, addr_positional[51091:51088], addr_12772_7);

wire[31:0] addr_12773_7;

Selector_2 s12773_7(wires_3193_6[1], addr_3193_6, addr_positional[51095:51092], addr_12773_7);

wire[31:0] addr_12774_7;

Selector_2 s12774_7(wires_3193_6[2], addr_3193_6, addr_positional[51099:51096], addr_12774_7);

wire[31:0] addr_12775_7;

Selector_2 s12775_7(wires_3193_6[3], addr_3193_6, addr_positional[51103:51100], addr_12775_7);

wire[31:0] addr_12776_7;

Selector_2 s12776_7(wires_3194_6[0], addr_3194_6, addr_positional[51107:51104], addr_12776_7);

wire[31:0] addr_12777_7;

Selector_2 s12777_7(wires_3194_6[1], addr_3194_6, addr_positional[51111:51108], addr_12777_7);

wire[31:0] addr_12778_7;

Selector_2 s12778_7(wires_3194_6[2], addr_3194_6, addr_positional[51115:51112], addr_12778_7);

wire[31:0] addr_12779_7;

Selector_2 s12779_7(wires_3194_6[3], addr_3194_6, addr_positional[51119:51116], addr_12779_7);

wire[31:0] addr_12780_7;

Selector_2 s12780_7(wires_3195_6[0], addr_3195_6, addr_positional[51123:51120], addr_12780_7);

wire[31:0] addr_12781_7;

Selector_2 s12781_7(wires_3195_6[1], addr_3195_6, addr_positional[51127:51124], addr_12781_7);

wire[31:0] addr_12782_7;

Selector_2 s12782_7(wires_3195_6[2], addr_3195_6, addr_positional[51131:51128], addr_12782_7);

wire[31:0] addr_12783_7;

Selector_2 s12783_7(wires_3195_6[3], addr_3195_6, addr_positional[51135:51132], addr_12783_7);

wire[31:0] addr_12784_7;

Selector_2 s12784_7(wires_3196_6[0], addr_3196_6, addr_positional[51139:51136], addr_12784_7);

wire[31:0] addr_12785_7;

Selector_2 s12785_7(wires_3196_6[1], addr_3196_6, addr_positional[51143:51140], addr_12785_7);

wire[31:0] addr_12786_7;

Selector_2 s12786_7(wires_3196_6[2], addr_3196_6, addr_positional[51147:51144], addr_12786_7);

wire[31:0] addr_12787_7;

Selector_2 s12787_7(wires_3196_6[3], addr_3196_6, addr_positional[51151:51148], addr_12787_7);

wire[31:0] addr_12788_7;

Selector_2 s12788_7(wires_3197_6[0], addr_3197_6, addr_positional[51155:51152], addr_12788_7);

wire[31:0] addr_12789_7;

Selector_2 s12789_7(wires_3197_6[1], addr_3197_6, addr_positional[51159:51156], addr_12789_7);

wire[31:0] addr_12790_7;

Selector_2 s12790_7(wires_3197_6[2], addr_3197_6, addr_positional[51163:51160], addr_12790_7);

wire[31:0] addr_12791_7;

Selector_2 s12791_7(wires_3197_6[3], addr_3197_6, addr_positional[51167:51164], addr_12791_7);

wire[31:0] addr_12792_7;

Selector_2 s12792_7(wires_3198_6[0], addr_3198_6, addr_positional[51171:51168], addr_12792_7);

wire[31:0] addr_12793_7;

Selector_2 s12793_7(wires_3198_6[1], addr_3198_6, addr_positional[51175:51172], addr_12793_7);

wire[31:0] addr_12794_7;

Selector_2 s12794_7(wires_3198_6[2], addr_3198_6, addr_positional[51179:51176], addr_12794_7);

wire[31:0] addr_12795_7;

Selector_2 s12795_7(wires_3198_6[3], addr_3198_6, addr_positional[51183:51180], addr_12795_7);

wire[31:0] addr_12796_7;

Selector_2 s12796_7(wires_3199_6[0], addr_3199_6, addr_positional[51187:51184], addr_12796_7);

wire[31:0] addr_12797_7;

Selector_2 s12797_7(wires_3199_6[1], addr_3199_6, addr_positional[51191:51188], addr_12797_7);

wire[31:0] addr_12798_7;

Selector_2 s12798_7(wires_3199_6[2], addr_3199_6, addr_positional[51195:51192], addr_12798_7);

wire[31:0] addr_12799_7;

Selector_2 s12799_7(wires_3199_6[3], addr_3199_6, addr_positional[51199:51196], addr_12799_7);

wire[31:0] addr_12800_7;

Selector_2 s12800_7(wires_3200_6[0], addr_3200_6, addr_positional[51203:51200], addr_12800_7);

wire[31:0] addr_12801_7;

Selector_2 s12801_7(wires_3200_6[1], addr_3200_6, addr_positional[51207:51204], addr_12801_7);

wire[31:0] addr_12802_7;

Selector_2 s12802_7(wires_3200_6[2], addr_3200_6, addr_positional[51211:51208], addr_12802_7);

wire[31:0] addr_12803_7;

Selector_2 s12803_7(wires_3200_6[3], addr_3200_6, addr_positional[51215:51212], addr_12803_7);

wire[31:0] addr_12804_7;

Selector_2 s12804_7(wires_3201_6[0], addr_3201_6, addr_positional[51219:51216], addr_12804_7);

wire[31:0] addr_12805_7;

Selector_2 s12805_7(wires_3201_6[1], addr_3201_6, addr_positional[51223:51220], addr_12805_7);

wire[31:0] addr_12806_7;

Selector_2 s12806_7(wires_3201_6[2], addr_3201_6, addr_positional[51227:51224], addr_12806_7);

wire[31:0] addr_12807_7;

Selector_2 s12807_7(wires_3201_6[3], addr_3201_6, addr_positional[51231:51228], addr_12807_7);

wire[31:0] addr_12808_7;

Selector_2 s12808_7(wires_3202_6[0], addr_3202_6, addr_positional[51235:51232], addr_12808_7);

wire[31:0] addr_12809_7;

Selector_2 s12809_7(wires_3202_6[1], addr_3202_6, addr_positional[51239:51236], addr_12809_7);

wire[31:0] addr_12810_7;

Selector_2 s12810_7(wires_3202_6[2], addr_3202_6, addr_positional[51243:51240], addr_12810_7);

wire[31:0] addr_12811_7;

Selector_2 s12811_7(wires_3202_6[3], addr_3202_6, addr_positional[51247:51244], addr_12811_7);

wire[31:0] addr_12812_7;

Selector_2 s12812_7(wires_3203_6[0], addr_3203_6, addr_positional[51251:51248], addr_12812_7);

wire[31:0] addr_12813_7;

Selector_2 s12813_7(wires_3203_6[1], addr_3203_6, addr_positional[51255:51252], addr_12813_7);

wire[31:0] addr_12814_7;

Selector_2 s12814_7(wires_3203_6[2], addr_3203_6, addr_positional[51259:51256], addr_12814_7);

wire[31:0] addr_12815_7;

Selector_2 s12815_7(wires_3203_6[3], addr_3203_6, addr_positional[51263:51260], addr_12815_7);

wire[31:0] addr_12816_7;

Selector_2 s12816_7(wires_3204_6[0], addr_3204_6, addr_positional[51267:51264], addr_12816_7);

wire[31:0] addr_12817_7;

Selector_2 s12817_7(wires_3204_6[1], addr_3204_6, addr_positional[51271:51268], addr_12817_7);

wire[31:0] addr_12818_7;

Selector_2 s12818_7(wires_3204_6[2], addr_3204_6, addr_positional[51275:51272], addr_12818_7);

wire[31:0] addr_12819_7;

Selector_2 s12819_7(wires_3204_6[3], addr_3204_6, addr_positional[51279:51276], addr_12819_7);

wire[31:0] addr_12820_7;

Selector_2 s12820_7(wires_3205_6[0], addr_3205_6, addr_positional[51283:51280], addr_12820_7);

wire[31:0] addr_12821_7;

Selector_2 s12821_7(wires_3205_6[1], addr_3205_6, addr_positional[51287:51284], addr_12821_7);

wire[31:0] addr_12822_7;

Selector_2 s12822_7(wires_3205_6[2], addr_3205_6, addr_positional[51291:51288], addr_12822_7);

wire[31:0] addr_12823_7;

Selector_2 s12823_7(wires_3205_6[3], addr_3205_6, addr_positional[51295:51292], addr_12823_7);

wire[31:0] addr_12824_7;

Selector_2 s12824_7(wires_3206_6[0], addr_3206_6, addr_positional[51299:51296], addr_12824_7);

wire[31:0] addr_12825_7;

Selector_2 s12825_7(wires_3206_6[1], addr_3206_6, addr_positional[51303:51300], addr_12825_7);

wire[31:0] addr_12826_7;

Selector_2 s12826_7(wires_3206_6[2], addr_3206_6, addr_positional[51307:51304], addr_12826_7);

wire[31:0] addr_12827_7;

Selector_2 s12827_7(wires_3206_6[3], addr_3206_6, addr_positional[51311:51308], addr_12827_7);

wire[31:0] addr_12828_7;

Selector_2 s12828_7(wires_3207_6[0], addr_3207_6, addr_positional[51315:51312], addr_12828_7);

wire[31:0] addr_12829_7;

Selector_2 s12829_7(wires_3207_6[1], addr_3207_6, addr_positional[51319:51316], addr_12829_7);

wire[31:0] addr_12830_7;

Selector_2 s12830_7(wires_3207_6[2], addr_3207_6, addr_positional[51323:51320], addr_12830_7);

wire[31:0] addr_12831_7;

Selector_2 s12831_7(wires_3207_6[3], addr_3207_6, addr_positional[51327:51324], addr_12831_7);

wire[31:0] addr_12832_7;

Selector_2 s12832_7(wires_3208_6[0], addr_3208_6, addr_positional[51331:51328], addr_12832_7);

wire[31:0] addr_12833_7;

Selector_2 s12833_7(wires_3208_6[1], addr_3208_6, addr_positional[51335:51332], addr_12833_7);

wire[31:0] addr_12834_7;

Selector_2 s12834_7(wires_3208_6[2], addr_3208_6, addr_positional[51339:51336], addr_12834_7);

wire[31:0] addr_12835_7;

Selector_2 s12835_7(wires_3208_6[3], addr_3208_6, addr_positional[51343:51340], addr_12835_7);

wire[31:0] addr_12836_7;

Selector_2 s12836_7(wires_3209_6[0], addr_3209_6, addr_positional[51347:51344], addr_12836_7);

wire[31:0] addr_12837_7;

Selector_2 s12837_7(wires_3209_6[1], addr_3209_6, addr_positional[51351:51348], addr_12837_7);

wire[31:0] addr_12838_7;

Selector_2 s12838_7(wires_3209_6[2], addr_3209_6, addr_positional[51355:51352], addr_12838_7);

wire[31:0] addr_12839_7;

Selector_2 s12839_7(wires_3209_6[3], addr_3209_6, addr_positional[51359:51356], addr_12839_7);

wire[31:0] addr_12840_7;

Selector_2 s12840_7(wires_3210_6[0], addr_3210_6, addr_positional[51363:51360], addr_12840_7);

wire[31:0] addr_12841_7;

Selector_2 s12841_7(wires_3210_6[1], addr_3210_6, addr_positional[51367:51364], addr_12841_7);

wire[31:0] addr_12842_7;

Selector_2 s12842_7(wires_3210_6[2], addr_3210_6, addr_positional[51371:51368], addr_12842_7);

wire[31:0] addr_12843_7;

Selector_2 s12843_7(wires_3210_6[3], addr_3210_6, addr_positional[51375:51372], addr_12843_7);

wire[31:0] addr_12844_7;

Selector_2 s12844_7(wires_3211_6[0], addr_3211_6, addr_positional[51379:51376], addr_12844_7);

wire[31:0] addr_12845_7;

Selector_2 s12845_7(wires_3211_6[1], addr_3211_6, addr_positional[51383:51380], addr_12845_7);

wire[31:0] addr_12846_7;

Selector_2 s12846_7(wires_3211_6[2], addr_3211_6, addr_positional[51387:51384], addr_12846_7);

wire[31:0] addr_12847_7;

Selector_2 s12847_7(wires_3211_6[3], addr_3211_6, addr_positional[51391:51388], addr_12847_7);

wire[31:0] addr_12848_7;

Selector_2 s12848_7(wires_3212_6[0], addr_3212_6, addr_positional[51395:51392], addr_12848_7);

wire[31:0] addr_12849_7;

Selector_2 s12849_7(wires_3212_6[1], addr_3212_6, addr_positional[51399:51396], addr_12849_7);

wire[31:0] addr_12850_7;

Selector_2 s12850_7(wires_3212_6[2], addr_3212_6, addr_positional[51403:51400], addr_12850_7);

wire[31:0] addr_12851_7;

Selector_2 s12851_7(wires_3212_6[3], addr_3212_6, addr_positional[51407:51404], addr_12851_7);

wire[31:0] addr_12852_7;

Selector_2 s12852_7(wires_3213_6[0], addr_3213_6, addr_positional[51411:51408], addr_12852_7);

wire[31:0] addr_12853_7;

Selector_2 s12853_7(wires_3213_6[1], addr_3213_6, addr_positional[51415:51412], addr_12853_7);

wire[31:0] addr_12854_7;

Selector_2 s12854_7(wires_3213_6[2], addr_3213_6, addr_positional[51419:51416], addr_12854_7);

wire[31:0] addr_12855_7;

Selector_2 s12855_7(wires_3213_6[3], addr_3213_6, addr_positional[51423:51420], addr_12855_7);

wire[31:0] addr_12856_7;

Selector_2 s12856_7(wires_3214_6[0], addr_3214_6, addr_positional[51427:51424], addr_12856_7);

wire[31:0] addr_12857_7;

Selector_2 s12857_7(wires_3214_6[1], addr_3214_6, addr_positional[51431:51428], addr_12857_7);

wire[31:0] addr_12858_7;

Selector_2 s12858_7(wires_3214_6[2], addr_3214_6, addr_positional[51435:51432], addr_12858_7);

wire[31:0] addr_12859_7;

Selector_2 s12859_7(wires_3214_6[3], addr_3214_6, addr_positional[51439:51436], addr_12859_7);

wire[31:0] addr_12860_7;

Selector_2 s12860_7(wires_3215_6[0], addr_3215_6, addr_positional[51443:51440], addr_12860_7);

wire[31:0] addr_12861_7;

Selector_2 s12861_7(wires_3215_6[1], addr_3215_6, addr_positional[51447:51444], addr_12861_7);

wire[31:0] addr_12862_7;

Selector_2 s12862_7(wires_3215_6[2], addr_3215_6, addr_positional[51451:51448], addr_12862_7);

wire[31:0] addr_12863_7;

Selector_2 s12863_7(wires_3215_6[3], addr_3215_6, addr_positional[51455:51452], addr_12863_7);

wire[31:0] addr_12864_7;

Selector_2 s12864_7(wires_3216_6[0], addr_3216_6, addr_positional[51459:51456], addr_12864_7);

wire[31:0] addr_12865_7;

Selector_2 s12865_7(wires_3216_6[1], addr_3216_6, addr_positional[51463:51460], addr_12865_7);

wire[31:0] addr_12866_7;

Selector_2 s12866_7(wires_3216_6[2], addr_3216_6, addr_positional[51467:51464], addr_12866_7);

wire[31:0] addr_12867_7;

Selector_2 s12867_7(wires_3216_6[3], addr_3216_6, addr_positional[51471:51468], addr_12867_7);

wire[31:0] addr_12868_7;

Selector_2 s12868_7(wires_3217_6[0], addr_3217_6, addr_positional[51475:51472], addr_12868_7);

wire[31:0] addr_12869_7;

Selector_2 s12869_7(wires_3217_6[1], addr_3217_6, addr_positional[51479:51476], addr_12869_7);

wire[31:0] addr_12870_7;

Selector_2 s12870_7(wires_3217_6[2], addr_3217_6, addr_positional[51483:51480], addr_12870_7);

wire[31:0] addr_12871_7;

Selector_2 s12871_7(wires_3217_6[3], addr_3217_6, addr_positional[51487:51484], addr_12871_7);

wire[31:0] addr_12872_7;

Selector_2 s12872_7(wires_3218_6[0], addr_3218_6, addr_positional[51491:51488], addr_12872_7);

wire[31:0] addr_12873_7;

Selector_2 s12873_7(wires_3218_6[1], addr_3218_6, addr_positional[51495:51492], addr_12873_7);

wire[31:0] addr_12874_7;

Selector_2 s12874_7(wires_3218_6[2], addr_3218_6, addr_positional[51499:51496], addr_12874_7);

wire[31:0] addr_12875_7;

Selector_2 s12875_7(wires_3218_6[3], addr_3218_6, addr_positional[51503:51500], addr_12875_7);

wire[31:0] addr_12876_7;

Selector_2 s12876_7(wires_3219_6[0], addr_3219_6, addr_positional[51507:51504], addr_12876_7);

wire[31:0] addr_12877_7;

Selector_2 s12877_7(wires_3219_6[1], addr_3219_6, addr_positional[51511:51508], addr_12877_7);

wire[31:0] addr_12878_7;

Selector_2 s12878_7(wires_3219_6[2], addr_3219_6, addr_positional[51515:51512], addr_12878_7);

wire[31:0] addr_12879_7;

Selector_2 s12879_7(wires_3219_6[3], addr_3219_6, addr_positional[51519:51516], addr_12879_7);

wire[31:0] addr_12880_7;

Selector_2 s12880_7(wires_3220_6[0], addr_3220_6, addr_positional[51523:51520], addr_12880_7);

wire[31:0] addr_12881_7;

Selector_2 s12881_7(wires_3220_6[1], addr_3220_6, addr_positional[51527:51524], addr_12881_7);

wire[31:0] addr_12882_7;

Selector_2 s12882_7(wires_3220_6[2], addr_3220_6, addr_positional[51531:51528], addr_12882_7);

wire[31:0] addr_12883_7;

Selector_2 s12883_7(wires_3220_6[3], addr_3220_6, addr_positional[51535:51532], addr_12883_7);

wire[31:0] addr_12884_7;

Selector_2 s12884_7(wires_3221_6[0], addr_3221_6, addr_positional[51539:51536], addr_12884_7);

wire[31:0] addr_12885_7;

Selector_2 s12885_7(wires_3221_6[1], addr_3221_6, addr_positional[51543:51540], addr_12885_7);

wire[31:0] addr_12886_7;

Selector_2 s12886_7(wires_3221_6[2], addr_3221_6, addr_positional[51547:51544], addr_12886_7);

wire[31:0] addr_12887_7;

Selector_2 s12887_7(wires_3221_6[3], addr_3221_6, addr_positional[51551:51548], addr_12887_7);

wire[31:0] addr_12888_7;

Selector_2 s12888_7(wires_3222_6[0], addr_3222_6, addr_positional[51555:51552], addr_12888_7);

wire[31:0] addr_12889_7;

Selector_2 s12889_7(wires_3222_6[1], addr_3222_6, addr_positional[51559:51556], addr_12889_7);

wire[31:0] addr_12890_7;

Selector_2 s12890_7(wires_3222_6[2], addr_3222_6, addr_positional[51563:51560], addr_12890_7);

wire[31:0] addr_12891_7;

Selector_2 s12891_7(wires_3222_6[3], addr_3222_6, addr_positional[51567:51564], addr_12891_7);

wire[31:0] addr_12892_7;

Selector_2 s12892_7(wires_3223_6[0], addr_3223_6, addr_positional[51571:51568], addr_12892_7);

wire[31:0] addr_12893_7;

Selector_2 s12893_7(wires_3223_6[1], addr_3223_6, addr_positional[51575:51572], addr_12893_7);

wire[31:0] addr_12894_7;

Selector_2 s12894_7(wires_3223_6[2], addr_3223_6, addr_positional[51579:51576], addr_12894_7);

wire[31:0] addr_12895_7;

Selector_2 s12895_7(wires_3223_6[3], addr_3223_6, addr_positional[51583:51580], addr_12895_7);

wire[31:0] addr_12896_7;

Selector_2 s12896_7(wires_3224_6[0], addr_3224_6, addr_positional[51587:51584], addr_12896_7);

wire[31:0] addr_12897_7;

Selector_2 s12897_7(wires_3224_6[1], addr_3224_6, addr_positional[51591:51588], addr_12897_7);

wire[31:0] addr_12898_7;

Selector_2 s12898_7(wires_3224_6[2], addr_3224_6, addr_positional[51595:51592], addr_12898_7);

wire[31:0] addr_12899_7;

Selector_2 s12899_7(wires_3224_6[3], addr_3224_6, addr_positional[51599:51596], addr_12899_7);

wire[31:0] addr_12900_7;

Selector_2 s12900_7(wires_3225_6[0], addr_3225_6, addr_positional[51603:51600], addr_12900_7);

wire[31:0] addr_12901_7;

Selector_2 s12901_7(wires_3225_6[1], addr_3225_6, addr_positional[51607:51604], addr_12901_7);

wire[31:0] addr_12902_7;

Selector_2 s12902_7(wires_3225_6[2], addr_3225_6, addr_positional[51611:51608], addr_12902_7);

wire[31:0] addr_12903_7;

Selector_2 s12903_7(wires_3225_6[3], addr_3225_6, addr_positional[51615:51612], addr_12903_7);

wire[31:0] addr_12904_7;

Selector_2 s12904_7(wires_3226_6[0], addr_3226_6, addr_positional[51619:51616], addr_12904_7);

wire[31:0] addr_12905_7;

Selector_2 s12905_7(wires_3226_6[1], addr_3226_6, addr_positional[51623:51620], addr_12905_7);

wire[31:0] addr_12906_7;

Selector_2 s12906_7(wires_3226_6[2], addr_3226_6, addr_positional[51627:51624], addr_12906_7);

wire[31:0] addr_12907_7;

Selector_2 s12907_7(wires_3226_6[3], addr_3226_6, addr_positional[51631:51628], addr_12907_7);

wire[31:0] addr_12908_7;

Selector_2 s12908_7(wires_3227_6[0], addr_3227_6, addr_positional[51635:51632], addr_12908_7);

wire[31:0] addr_12909_7;

Selector_2 s12909_7(wires_3227_6[1], addr_3227_6, addr_positional[51639:51636], addr_12909_7);

wire[31:0] addr_12910_7;

Selector_2 s12910_7(wires_3227_6[2], addr_3227_6, addr_positional[51643:51640], addr_12910_7);

wire[31:0] addr_12911_7;

Selector_2 s12911_7(wires_3227_6[3], addr_3227_6, addr_positional[51647:51644], addr_12911_7);

wire[31:0] addr_12912_7;

Selector_2 s12912_7(wires_3228_6[0], addr_3228_6, addr_positional[51651:51648], addr_12912_7);

wire[31:0] addr_12913_7;

Selector_2 s12913_7(wires_3228_6[1], addr_3228_6, addr_positional[51655:51652], addr_12913_7);

wire[31:0] addr_12914_7;

Selector_2 s12914_7(wires_3228_6[2], addr_3228_6, addr_positional[51659:51656], addr_12914_7);

wire[31:0] addr_12915_7;

Selector_2 s12915_7(wires_3228_6[3], addr_3228_6, addr_positional[51663:51660], addr_12915_7);

wire[31:0] addr_12916_7;

Selector_2 s12916_7(wires_3229_6[0], addr_3229_6, addr_positional[51667:51664], addr_12916_7);

wire[31:0] addr_12917_7;

Selector_2 s12917_7(wires_3229_6[1], addr_3229_6, addr_positional[51671:51668], addr_12917_7);

wire[31:0] addr_12918_7;

Selector_2 s12918_7(wires_3229_6[2], addr_3229_6, addr_positional[51675:51672], addr_12918_7);

wire[31:0] addr_12919_7;

Selector_2 s12919_7(wires_3229_6[3], addr_3229_6, addr_positional[51679:51676], addr_12919_7);

wire[31:0] addr_12920_7;

Selector_2 s12920_7(wires_3230_6[0], addr_3230_6, addr_positional[51683:51680], addr_12920_7);

wire[31:0] addr_12921_7;

Selector_2 s12921_7(wires_3230_6[1], addr_3230_6, addr_positional[51687:51684], addr_12921_7);

wire[31:0] addr_12922_7;

Selector_2 s12922_7(wires_3230_6[2], addr_3230_6, addr_positional[51691:51688], addr_12922_7);

wire[31:0] addr_12923_7;

Selector_2 s12923_7(wires_3230_6[3], addr_3230_6, addr_positional[51695:51692], addr_12923_7);

wire[31:0] addr_12924_7;

Selector_2 s12924_7(wires_3231_6[0], addr_3231_6, addr_positional[51699:51696], addr_12924_7);

wire[31:0] addr_12925_7;

Selector_2 s12925_7(wires_3231_6[1], addr_3231_6, addr_positional[51703:51700], addr_12925_7);

wire[31:0] addr_12926_7;

Selector_2 s12926_7(wires_3231_6[2], addr_3231_6, addr_positional[51707:51704], addr_12926_7);

wire[31:0] addr_12927_7;

Selector_2 s12927_7(wires_3231_6[3], addr_3231_6, addr_positional[51711:51708], addr_12927_7);

wire[31:0] addr_12928_7;

Selector_2 s12928_7(wires_3232_6[0], addr_3232_6, addr_positional[51715:51712], addr_12928_7);

wire[31:0] addr_12929_7;

Selector_2 s12929_7(wires_3232_6[1], addr_3232_6, addr_positional[51719:51716], addr_12929_7);

wire[31:0] addr_12930_7;

Selector_2 s12930_7(wires_3232_6[2], addr_3232_6, addr_positional[51723:51720], addr_12930_7);

wire[31:0] addr_12931_7;

Selector_2 s12931_7(wires_3232_6[3], addr_3232_6, addr_positional[51727:51724], addr_12931_7);

wire[31:0] addr_12932_7;

Selector_2 s12932_7(wires_3233_6[0], addr_3233_6, addr_positional[51731:51728], addr_12932_7);

wire[31:0] addr_12933_7;

Selector_2 s12933_7(wires_3233_6[1], addr_3233_6, addr_positional[51735:51732], addr_12933_7);

wire[31:0] addr_12934_7;

Selector_2 s12934_7(wires_3233_6[2], addr_3233_6, addr_positional[51739:51736], addr_12934_7);

wire[31:0] addr_12935_7;

Selector_2 s12935_7(wires_3233_6[3], addr_3233_6, addr_positional[51743:51740], addr_12935_7);

wire[31:0] addr_12936_7;

Selector_2 s12936_7(wires_3234_6[0], addr_3234_6, addr_positional[51747:51744], addr_12936_7);

wire[31:0] addr_12937_7;

Selector_2 s12937_7(wires_3234_6[1], addr_3234_6, addr_positional[51751:51748], addr_12937_7);

wire[31:0] addr_12938_7;

Selector_2 s12938_7(wires_3234_6[2], addr_3234_6, addr_positional[51755:51752], addr_12938_7);

wire[31:0] addr_12939_7;

Selector_2 s12939_7(wires_3234_6[3], addr_3234_6, addr_positional[51759:51756], addr_12939_7);

wire[31:0] addr_12940_7;

Selector_2 s12940_7(wires_3235_6[0], addr_3235_6, addr_positional[51763:51760], addr_12940_7);

wire[31:0] addr_12941_7;

Selector_2 s12941_7(wires_3235_6[1], addr_3235_6, addr_positional[51767:51764], addr_12941_7);

wire[31:0] addr_12942_7;

Selector_2 s12942_7(wires_3235_6[2], addr_3235_6, addr_positional[51771:51768], addr_12942_7);

wire[31:0] addr_12943_7;

Selector_2 s12943_7(wires_3235_6[3], addr_3235_6, addr_positional[51775:51772], addr_12943_7);

wire[31:0] addr_12944_7;

Selector_2 s12944_7(wires_3236_6[0], addr_3236_6, addr_positional[51779:51776], addr_12944_7);

wire[31:0] addr_12945_7;

Selector_2 s12945_7(wires_3236_6[1], addr_3236_6, addr_positional[51783:51780], addr_12945_7);

wire[31:0] addr_12946_7;

Selector_2 s12946_7(wires_3236_6[2], addr_3236_6, addr_positional[51787:51784], addr_12946_7);

wire[31:0] addr_12947_7;

Selector_2 s12947_7(wires_3236_6[3], addr_3236_6, addr_positional[51791:51788], addr_12947_7);

wire[31:0] addr_12948_7;

Selector_2 s12948_7(wires_3237_6[0], addr_3237_6, addr_positional[51795:51792], addr_12948_7);

wire[31:0] addr_12949_7;

Selector_2 s12949_7(wires_3237_6[1], addr_3237_6, addr_positional[51799:51796], addr_12949_7);

wire[31:0] addr_12950_7;

Selector_2 s12950_7(wires_3237_6[2], addr_3237_6, addr_positional[51803:51800], addr_12950_7);

wire[31:0] addr_12951_7;

Selector_2 s12951_7(wires_3237_6[3], addr_3237_6, addr_positional[51807:51804], addr_12951_7);

wire[31:0] addr_12952_7;

Selector_2 s12952_7(wires_3238_6[0], addr_3238_6, addr_positional[51811:51808], addr_12952_7);

wire[31:0] addr_12953_7;

Selector_2 s12953_7(wires_3238_6[1], addr_3238_6, addr_positional[51815:51812], addr_12953_7);

wire[31:0] addr_12954_7;

Selector_2 s12954_7(wires_3238_6[2], addr_3238_6, addr_positional[51819:51816], addr_12954_7);

wire[31:0] addr_12955_7;

Selector_2 s12955_7(wires_3238_6[3], addr_3238_6, addr_positional[51823:51820], addr_12955_7);

wire[31:0] addr_12956_7;

Selector_2 s12956_7(wires_3239_6[0], addr_3239_6, addr_positional[51827:51824], addr_12956_7);

wire[31:0] addr_12957_7;

Selector_2 s12957_7(wires_3239_6[1], addr_3239_6, addr_positional[51831:51828], addr_12957_7);

wire[31:0] addr_12958_7;

Selector_2 s12958_7(wires_3239_6[2], addr_3239_6, addr_positional[51835:51832], addr_12958_7);

wire[31:0] addr_12959_7;

Selector_2 s12959_7(wires_3239_6[3], addr_3239_6, addr_positional[51839:51836], addr_12959_7);

wire[31:0] addr_12960_7;

Selector_2 s12960_7(wires_3240_6[0], addr_3240_6, addr_positional[51843:51840], addr_12960_7);

wire[31:0] addr_12961_7;

Selector_2 s12961_7(wires_3240_6[1], addr_3240_6, addr_positional[51847:51844], addr_12961_7);

wire[31:0] addr_12962_7;

Selector_2 s12962_7(wires_3240_6[2], addr_3240_6, addr_positional[51851:51848], addr_12962_7);

wire[31:0] addr_12963_7;

Selector_2 s12963_7(wires_3240_6[3], addr_3240_6, addr_positional[51855:51852], addr_12963_7);

wire[31:0] addr_12964_7;

Selector_2 s12964_7(wires_3241_6[0], addr_3241_6, addr_positional[51859:51856], addr_12964_7);

wire[31:0] addr_12965_7;

Selector_2 s12965_7(wires_3241_6[1], addr_3241_6, addr_positional[51863:51860], addr_12965_7);

wire[31:0] addr_12966_7;

Selector_2 s12966_7(wires_3241_6[2], addr_3241_6, addr_positional[51867:51864], addr_12966_7);

wire[31:0] addr_12967_7;

Selector_2 s12967_7(wires_3241_6[3], addr_3241_6, addr_positional[51871:51868], addr_12967_7);

wire[31:0] addr_12968_7;

Selector_2 s12968_7(wires_3242_6[0], addr_3242_6, addr_positional[51875:51872], addr_12968_7);

wire[31:0] addr_12969_7;

Selector_2 s12969_7(wires_3242_6[1], addr_3242_6, addr_positional[51879:51876], addr_12969_7);

wire[31:0] addr_12970_7;

Selector_2 s12970_7(wires_3242_6[2], addr_3242_6, addr_positional[51883:51880], addr_12970_7);

wire[31:0] addr_12971_7;

Selector_2 s12971_7(wires_3242_6[3], addr_3242_6, addr_positional[51887:51884], addr_12971_7);

wire[31:0] addr_12972_7;

Selector_2 s12972_7(wires_3243_6[0], addr_3243_6, addr_positional[51891:51888], addr_12972_7);

wire[31:0] addr_12973_7;

Selector_2 s12973_7(wires_3243_6[1], addr_3243_6, addr_positional[51895:51892], addr_12973_7);

wire[31:0] addr_12974_7;

Selector_2 s12974_7(wires_3243_6[2], addr_3243_6, addr_positional[51899:51896], addr_12974_7);

wire[31:0] addr_12975_7;

Selector_2 s12975_7(wires_3243_6[3], addr_3243_6, addr_positional[51903:51900], addr_12975_7);

wire[31:0] addr_12976_7;

Selector_2 s12976_7(wires_3244_6[0], addr_3244_6, addr_positional[51907:51904], addr_12976_7);

wire[31:0] addr_12977_7;

Selector_2 s12977_7(wires_3244_6[1], addr_3244_6, addr_positional[51911:51908], addr_12977_7);

wire[31:0] addr_12978_7;

Selector_2 s12978_7(wires_3244_6[2], addr_3244_6, addr_positional[51915:51912], addr_12978_7);

wire[31:0] addr_12979_7;

Selector_2 s12979_7(wires_3244_6[3], addr_3244_6, addr_positional[51919:51916], addr_12979_7);

wire[31:0] addr_12980_7;

Selector_2 s12980_7(wires_3245_6[0], addr_3245_6, addr_positional[51923:51920], addr_12980_7);

wire[31:0] addr_12981_7;

Selector_2 s12981_7(wires_3245_6[1], addr_3245_6, addr_positional[51927:51924], addr_12981_7);

wire[31:0] addr_12982_7;

Selector_2 s12982_7(wires_3245_6[2], addr_3245_6, addr_positional[51931:51928], addr_12982_7);

wire[31:0] addr_12983_7;

Selector_2 s12983_7(wires_3245_6[3], addr_3245_6, addr_positional[51935:51932], addr_12983_7);

wire[31:0] addr_12984_7;

Selector_2 s12984_7(wires_3246_6[0], addr_3246_6, addr_positional[51939:51936], addr_12984_7);

wire[31:0] addr_12985_7;

Selector_2 s12985_7(wires_3246_6[1], addr_3246_6, addr_positional[51943:51940], addr_12985_7);

wire[31:0] addr_12986_7;

Selector_2 s12986_7(wires_3246_6[2], addr_3246_6, addr_positional[51947:51944], addr_12986_7);

wire[31:0] addr_12987_7;

Selector_2 s12987_7(wires_3246_6[3], addr_3246_6, addr_positional[51951:51948], addr_12987_7);

wire[31:0] addr_12988_7;

Selector_2 s12988_7(wires_3247_6[0], addr_3247_6, addr_positional[51955:51952], addr_12988_7);

wire[31:0] addr_12989_7;

Selector_2 s12989_7(wires_3247_6[1], addr_3247_6, addr_positional[51959:51956], addr_12989_7);

wire[31:0] addr_12990_7;

Selector_2 s12990_7(wires_3247_6[2], addr_3247_6, addr_positional[51963:51960], addr_12990_7);

wire[31:0] addr_12991_7;

Selector_2 s12991_7(wires_3247_6[3], addr_3247_6, addr_positional[51967:51964], addr_12991_7);

wire[31:0] addr_12992_7;

Selector_2 s12992_7(wires_3248_6[0], addr_3248_6, addr_positional[51971:51968], addr_12992_7);

wire[31:0] addr_12993_7;

Selector_2 s12993_7(wires_3248_6[1], addr_3248_6, addr_positional[51975:51972], addr_12993_7);

wire[31:0] addr_12994_7;

Selector_2 s12994_7(wires_3248_6[2], addr_3248_6, addr_positional[51979:51976], addr_12994_7);

wire[31:0] addr_12995_7;

Selector_2 s12995_7(wires_3248_6[3], addr_3248_6, addr_positional[51983:51980], addr_12995_7);

wire[31:0] addr_12996_7;

Selector_2 s12996_7(wires_3249_6[0], addr_3249_6, addr_positional[51987:51984], addr_12996_7);

wire[31:0] addr_12997_7;

Selector_2 s12997_7(wires_3249_6[1], addr_3249_6, addr_positional[51991:51988], addr_12997_7);

wire[31:0] addr_12998_7;

Selector_2 s12998_7(wires_3249_6[2], addr_3249_6, addr_positional[51995:51992], addr_12998_7);

wire[31:0] addr_12999_7;

Selector_2 s12999_7(wires_3249_6[3], addr_3249_6, addr_positional[51999:51996], addr_12999_7);

wire[31:0] addr_13000_7;

Selector_2 s13000_7(wires_3250_6[0], addr_3250_6, addr_positional[52003:52000], addr_13000_7);

wire[31:0] addr_13001_7;

Selector_2 s13001_7(wires_3250_6[1], addr_3250_6, addr_positional[52007:52004], addr_13001_7);

wire[31:0] addr_13002_7;

Selector_2 s13002_7(wires_3250_6[2], addr_3250_6, addr_positional[52011:52008], addr_13002_7);

wire[31:0] addr_13003_7;

Selector_2 s13003_7(wires_3250_6[3], addr_3250_6, addr_positional[52015:52012], addr_13003_7);

wire[31:0] addr_13004_7;

Selector_2 s13004_7(wires_3251_6[0], addr_3251_6, addr_positional[52019:52016], addr_13004_7);

wire[31:0] addr_13005_7;

Selector_2 s13005_7(wires_3251_6[1], addr_3251_6, addr_positional[52023:52020], addr_13005_7);

wire[31:0] addr_13006_7;

Selector_2 s13006_7(wires_3251_6[2], addr_3251_6, addr_positional[52027:52024], addr_13006_7);

wire[31:0] addr_13007_7;

Selector_2 s13007_7(wires_3251_6[3], addr_3251_6, addr_positional[52031:52028], addr_13007_7);

wire[31:0] addr_13008_7;

Selector_2 s13008_7(wires_3252_6[0], addr_3252_6, addr_positional[52035:52032], addr_13008_7);

wire[31:0] addr_13009_7;

Selector_2 s13009_7(wires_3252_6[1], addr_3252_6, addr_positional[52039:52036], addr_13009_7);

wire[31:0] addr_13010_7;

Selector_2 s13010_7(wires_3252_6[2], addr_3252_6, addr_positional[52043:52040], addr_13010_7);

wire[31:0] addr_13011_7;

Selector_2 s13011_7(wires_3252_6[3], addr_3252_6, addr_positional[52047:52044], addr_13011_7);

wire[31:0] addr_13012_7;

Selector_2 s13012_7(wires_3253_6[0], addr_3253_6, addr_positional[52051:52048], addr_13012_7);

wire[31:0] addr_13013_7;

Selector_2 s13013_7(wires_3253_6[1], addr_3253_6, addr_positional[52055:52052], addr_13013_7);

wire[31:0] addr_13014_7;

Selector_2 s13014_7(wires_3253_6[2], addr_3253_6, addr_positional[52059:52056], addr_13014_7);

wire[31:0] addr_13015_7;

Selector_2 s13015_7(wires_3253_6[3], addr_3253_6, addr_positional[52063:52060], addr_13015_7);

wire[31:0] addr_13016_7;

Selector_2 s13016_7(wires_3254_6[0], addr_3254_6, addr_positional[52067:52064], addr_13016_7);

wire[31:0] addr_13017_7;

Selector_2 s13017_7(wires_3254_6[1], addr_3254_6, addr_positional[52071:52068], addr_13017_7);

wire[31:0] addr_13018_7;

Selector_2 s13018_7(wires_3254_6[2], addr_3254_6, addr_positional[52075:52072], addr_13018_7);

wire[31:0] addr_13019_7;

Selector_2 s13019_7(wires_3254_6[3], addr_3254_6, addr_positional[52079:52076], addr_13019_7);

wire[31:0] addr_13020_7;

Selector_2 s13020_7(wires_3255_6[0], addr_3255_6, addr_positional[52083:52080], addr_13020_7);

wire[31:0] addr_13021_7;

Selector_2 s13021_7(wires_3255_6[1], addr_3255_6, addr_positional[52087:52084], addr_13021_7);

wire[31:0] addr_13022_7;

Selector_2 s13022_7(wires_3255_6[2], addr_3255_6, addr_positional[52091:52088], addr_13022_7);

wire[31:0] addr_13023_7;

Selector_2 s13023_7(wires_3255_6[3], addr_3255_6, addr_positional[52095:52092], addr_13023_7);

wire[31:0] addr_13024_7;

Selector_2 s13024_7(wires_3256_6[0], addr_3256_6, addr_positional[52099:52096], addr_13024_7);

wire[31:0] addr_13025_7;

Selector_2 s13025_7(wires_3256_6[1], addr_3256_6, addr_positional[52103:52100], addr_13025_7);

wire[31:0] addr_13026_7;

Selector_2 s13026_7(wires_3256_6[2], addr_3256_6, addr_positional[52107:52104], addr_13026_7);

wire[31:0] addr_13027_7;

Selector_2 s13027_7(wires_3256_6[3], addr_3256_6, addr_positional[52111:52108], addr_13027_7);

wire[31:0] addr_13028_7;

Selector_2 s13028_7(wires_3257_6[0], addr_3257_6, addr_positional[52115:52112], addr_13028_7);

wire[31:0] addr_13029_7;

Selector_2 s13029_7(wires_3257_6[1], addr_3257_6, addr_positional[52119:52116], addr_13029_7);

wire[31:0] addr_13030_7;

Selector_2 s13030_7(wires_3257_6[2], addr_3257_6, addr_positional[52123:52120], addr_13030_7);

wire[31:0] addr_13031_7;

Selector_2 s13031_7(wires_3257_6[3], addr_3257_6, addr_positional[52127:52124], addr_13031_7);

wire[31:0] addr_13032_7;

Selector_2 s13032_7(wires_3258_6[0], addr_3258_6, addr_positional[52131:52128], addr_13032_7);

wire[31:0] addr_13033_7;

Selector_2 s13033_7(wires_3258_6[1], addr_3258_6, addr_positional[52135:52132], addr_13033_7);

wire[31:0] addr_13034_7;

Selector_2 s13034_7(wires_3258_6[2], addr_3258_6, addr_positional[52139:52136], addr_13034_7);

wire[31:0] addr_13035_7;

Selector_2 s13035_7(wires_3258_6[3], addr_3258_6, addr_positional[52143:52140], addr_13035_7);

wire[31:0] addr_13036_7;

Selector_2 s13036_7(wires_3259_6[0], addr_3259_6, addr_positional[52147:52144], addr_13036_7);

wire[31:0] addr_13037_7;

Selector_2 s13037_7(wires_3259_6[1], addr_3259_6, addr_positional[52151:52148], addr_13037_7);

wire[31:0] addr_13038_7;

Selector_2 s13038_7(wires_3259_6[2], addr_3259_6, addr_positional[52155:52152], addr_13038_7);

wire[31:0] addr_13039_7;

Selector_2 s13039_7(wires_3259_6[3], addr_3259_6, addr_positional[52159:52156], addr_13039_7);

wire[31:0] addr_13040_7;

Selector_2 s13040_7(wires_3260_6[0], addr_3260_6, addr_positional[52163:52160], addr_13040_7);

wire[31:0] addr_13041_7;

Selector_2 s13041_7(wires_3260_6[1], addr_3260_6, addr_positional[52167:52164], addr_13041_7);

wire[31:0] addr_13042_7;

Selector_2 s13042_7(wires_3260_6[2], addr_3260_6, addr_positional[52171:52168], addr_13042_7);

wire[31:0] addr_13043_7;

Selector_2 s13043_7(wires_3260_6[3], addr_3260_6, addr_positional[52175:52172], addr_13043_7);

wire[31:0] addr_13044_7;

Selector_2 s13044_7(wires_3261_6[0], addr_3261_6, addr_positional[52179:52176], addr_13044_7);

wire[31:0] addr_13045_7;

Selector_2 s13045_7(wires_3261_6[1], addr_3261_6, addr_positional[52183:52180], addr_13045_7);

wire[31:0] addr_13046_7;

Selector_2 s13046_7(wires_3261_6[2], addr_3261_6, addr_positional[52187:52184], addr_13046_7);

wire[31:0] addr_13047_7;

Selector_2 s13047_7(wires_3261_6[3], addr_3261_6, addr_positional[52191:52188], addr_13047_7);

wire[31:0] addr_13048_7;

Selector_2 s13048_7(wires_3262_6[0], addr_3262_6, addr_positional[52195:52192], addr_13048_7);

wire[31:0] addr_13049_7;

Selector_2 s13049_7(wires_3262_6[1], addr_3262_6, addr_positional[52199:52196], addr_13049_7);

wire[31:0] addr_13050_7;

Selector_2 s13050_7(wires_3262_6[2], addr_3262_6, addr_positional[52203:52200], addr_13050_7);

wire[31:0] addr_13051_7;

Selector_2 s13051_7(wires_3262_6[3], addr_3262_6, addr_positional[52207:52204], addr_13051_7);

wire[31:0] addr_13052_7;

Selector_2 s13052_7(wires_3263_6[0], addr_3263_6, addr_positional[52211:52208], addr_13052_7);

wire[31:0] addr_13053_7;

Selector_2 s13053_7(wires_3263_6[1], addr_3263_6, addr_positional[52215:52212], addr_13053_7);

wire[31:0] addr_13054_7;

Selector_2 s13054_7(wires_3263_6[2], addr_3263_6, addr_positional[52219:52216], addr_13054_7);

wire[31:0] addr_13055_7;

Selector_2 s13055_7(wires_3263_6[3], addr_3263_6, addr_positional[52223:52220], addr_13055_7);

wire[31:0] addr_13056_7;

Selector_2 s13056_7(wires_3264_6[0], addr_3264_6, addr_positional[52227:52224], addr_13056_7);

wire[31:0] addr_13057_7;

Selector_2 s13057_7(wires_3264_6[1], addr_3264_6, addr_positional[52231:52228], addr_13057_7);

wire[31:0] addr_13058_7;

Selector_2 s13058_7(wires_3264_6[2], addr_3264_6, addr_positional[52235:52232], addr_13058_7);

wire[31:0] addr_13059_7;

Selector_2 s13059_7(wires_3264_6[3], addr_3264_6, addr_positional[52239:52236], addr_13059_7);

wire[31:0] addr_13060_7;

Selector_2 s13060_7(wires_3265_6[0], addr_3265_6, addr_positional[52243:52240], addr_13060_7);

wire[31:0] addr_13061_7;

Selector_2 s13061_7(wires_3265_6[1], addr_3265_6, addr_positional[52247:52244], addr_13061_7);

wire[31:0] addr_13062_7;

Selector_2 s13062_7(wires_3265_6[2], addr_3265_6, addr_positional[52251:52248], addr_13062_7);

wire[31:0] addr_13063_7;

Selector_2 s13063_7(wires_3265_6[3], addr_3265_6, addr_positional[52255:52252], addr_13063_7);

wire[31:0] addr_13064_7;

Selector_2 s13064_7(wires_3266_6[0], addr_3266_6, addr_positional[52259:52256], addr_13064_7);

wire[31:0] addr_13065_7;

Selector_2 s13065_7(wires_3266_6[1], addr_3266_6, addr_positional[52263:52260], addr_13065_7);

wire[31:0] addr_13066_7;

Selector_2 s13066_7(wires_3266_6[2], addr_3266_6, addr_positional[52267:52264], addr_13066_7);

wire[31:0] addr_13067_7;

Selector_2 s13067_7(wires_3266_6[3], addr_3266_6, addr_positional[52271:52268], addr_13067_7);

wire[31:0] addr_13068_7;

Selector_2 s13068_7(wires_3267_6[0], addr_3267_6, addr_positional[52275:52272], addr_13068_7);

wire[31:0] addr_13069_7;

Selector_2 s13069_7(wires_3267_6[1], addr_3267_6, addr_positional[52279:52276], addr_13069_7);

wire[31:0] addr_13070_7;

Selector_2 s13070_7(wires_3267_6[2], addr_3267_6, addr_positional[52283:52280], addr_13070_7);

wire[31:0] addr_13071_7;

Selector_2 s13071_7(wires_3267_6[3], addr_3267_6, addr_positional[52287:52284], addr_13071_7);

wire[31:0] addr_13072_7;

Selector_2 s13072_7(wires_3268_6[0], addr_3268_6, addr_positional[52291:52288], addr_13072_7);

wire[31:0] addr_13073_7;

Selector_2 s13073_7(wires_3268_6[1], addr_3268_6, addr_positional[52295:52292], addr_13073_7);

wire[31:0] addr_13074_7;

Selector_2 s13074_7(wires_3268_6[2], addr_3268_6, addr_positional[52299:52296], addr_13074_7);

wire[31:0] addr_13075_7;

Selector_2 s13075_7(wires_3268_6[3], addr_3268_6, addr_positional[52303:52300], addr_13075_7);

wire[31:0] addr_13076_7;

Selector_2 s13076_7(wires_3269_6[0], addr_3269_6, addr_positional[52307:52304], addr_13076_7);

wire[31:0] addr_13077_7;

Selector_2 s13077_7(wires_3269_6[1], addr_3269_6, addr_positional[52311:52308], addr_13077_7);

wire[31:0] addr_13078_7;

Selector_2 s13078_7(wires_3269_6[2], addr_3269_6, addr_positional[52315:52312], addr_13078_7);

wire[31:0] addr_13079_7;

Selector_2 s13079_7(wires_3269_6[3], addr_3269_6, addr_positional[52319:52316], addr_13079_7);

wire[31:0] addr_13080_7;

Selector_2 s13080_7(wires_3270_6[0], addr_3270_6, addr_positional[52323:52320], addr_13080_7);

wire[31:0] addr_13081_7;

Selector_2 s13081_7(wires_3270_6[1], addr_3270_6, addr_positional[52327:52324], addr_13081_7);

wire[31:0] addr_13082_7;

Selector_2 s13082_7(wires_3270_6[2], addr_3270_6, addr_positional[52331:52328], addr_13082_7);

wire[31:0] addr_13083_7;

Selector_2 s13083_7(wires_3270_6[3], addr_3270_6, addr_positional[52335:52332], addr_13083_7);

wire[31:0] addr_13084_7;

Selector_2 s13084_7(wires_3271_6[0], addr_3271_6, addr_positional[52339:52336], addr_13084_7);

wire[31:0] addr_13085_7;

Selector_2 s13085_7(wires_3271_6[1], addr_3271_6, addr_positional[52343:52340], addr_13085_7);

wire[31:0] addr_13086_7;

Selector_2 s13086_7(wires_3271_6[2], addr_3271_6, addr_positional[52347:52344], addr_13086_7);

wire[31:0] addr_13087_7;

Selector_2 s13087_7(wires_3271_6[3], addr_3271_6, addr_positional[52351:52348], addr_13087_7);

wire[31:0] addr_13088_7;

Selector_2 s13088_7(wires_3272_6[0], addr_3272_6, addr_positional[52355:52352], addr_13088_7);

wire[31:0] addr_13089_7;

Selector_2 s13089_7(wires_3272_6[1], addr_3272_6, addr_positional[52359:52356], addr_13089_7);

wire[31:0] addr_13090_7;

Selector_2 s13090_7(wires_3272_6[2], addr_3272_6, addr_positional[52363:52360], addr_13090_7);

wire[31:0] addr_13091_7;

Selector_2 s13091_7(wires_3272_6[3], addr_3272_6, addr_positional[52367:52364], addr_13091_7);

wire[31:0] addr_13092_7;

Selector_2 s13092_7(wires_3273_6[0], addr_3273_6, addr_positional[52371:52368], addr_13092_7);

wire[31:0] addr_13093_7;

Selector_2 s13093_7(wires_3273_6[1], addr_3273_6, addr_positional[52375:52372], addr_13093_7);

wire[31:0] addr_13094_7;

Selector_2 s13094_7(wires_3273_6[2], addr_3273_6, addr_positional[52379:52376], addr_13094_7);

wire[31:0] addr_13095_7;

Selector_2 s13095_7(wires_3273_6[3], addr_3273_6, addr_positional[52383:52380], addr_13095_7);

wire[31:0] addr_13096_7;

Selector_2 s13096_7(wires_3274_6[0], addr_3274_6, addr_positional[52387:52384], addr_13096_7);

wire[31:0] addr_13097_7;

Selector_2 s13097_7(wires_3274_6[1], addr_3274_6, addr_positional[52391:52388], addr_13097_7);

wire[31:0] addr_13098_7;

Selector_2 s13098_7(wires_3274_6[2], addr_3274_6, addr_positional[52395:52392], addr_13098_7);

wire[31:0] addr_13099_7;

Selector_2 s13099_7(wires_3274_6[3], addr_3274_6, addr_positional[52399:52396], addr_13099_7);

wire[31:0] addr_13100_7;

Selector_2 s13100_7(wires_3275_6[0], addr_3275_6, addr_positional[52403:52400], addr_13100_7);

wire[31:0] addr_13101_7;

Selector_2 s13101_7(wires_3275_6[1], addr_3275_6, addr_positional[52407:52404], addr_13101_7);

wire[31:0] addr_13102_7;

Selector_2 s13102_7(wires_3275_6[2], addr_3275_6, addr_positional[52411:52408], addr_13102_7);

wire[31:0] addr_13103_7;

Selector_2 s13103_7(wires_3275_6[3], addr_3275_6, addr_positional[52415:52412], addr_13103_7);

wire[31:0] addr_13104_7;

Selector_2 s13104_7(wires_3276_6[0], addr_3276_6, addr_positional[52419:52416], addr_13104_7);

wire[31:0] addr_13105_7;

Selector_2 s13105_7(wires_3276_6[1], addr_3276_6, addr_positional[52423:52420], addr_13105_7);

wire[31:0] addr_13106_7;

Selector_2 s13106_7(wires_3276_6[2], addr_3276_6, addr_positional[52427:52424], addr_13106_7);

wire[31:0] addr_13107_7;

Selector_2 s13107_7(wires_3276_6[3], addr_3276_6, addr_positional[52431:52428], addr_13107_7);

wire[31:0] addr_13108_7;

Selector_2 s13108_7(wires_3277_6[0], addr_3277_6, addr_positional[52435:52432], addr_13108_7);

wire[31:0] addr_13109_7;

Selector_2 s13109_7(wires_3277_6[1], addr_3277_6, addr_positional[52439:52436], addr_13109_7);

wire[31:0] addr_13110_7;

Selector_2 s13110_7(wires_3277_6[2], addr_3277_6, addr_positional[52443:52440], addr_13110_7);

wire[31:0] addr_13111_7;

Selector_2 s13111_7(wires_3277_6[3], addr_3277_6, addr_positional[52447:52444], addr_13111_7);

wire[31:0] addr_13112_7;

Selector_2 s13112_7(wires_3278_6[0], addr_3278_6, addr_positional[52451:52448], addr_13112_7);

wire[31:0] addr_13113_7;

Selector_2 s13113_7(wires_3278_6[1], addr_3278_6, addr_positional[52455:52452], addr_13113_7);

wire[31:0] addr_13114_7;

Selector_2 s13114_7(wires_3278_6[2], addr_3278_6, addr_positional[52459:52456], addr_13114_7);

wire[31:0] addr_13115_7;

Selector_2 s13115_7(wires_3278_6[3], addr_3278_6, addr_positional[52463:52460], addr_13115_7);

wire[31:0] addr_13116_7;

Selector_2 s13116_7(wires_3279_6[0], addr_3279_6, addr_positional[52467:52464], addr_13116_7);

wire[31:0] addr_13117_7;

Selector_2 s13117_7(wires_3279_6[1], addr_3279_6, addr_positional[52471:52468], addr_13117_7);

wire[31:0] addr_13118_7;

Selector_2 s13118_7(wires_3279_6[2], addr_3279_6, addr_positional[52475:52472], addr_13118_7);

wire[31:0] addr_13119_7;

Selector_2 s13119_7(wires_3279_6[3], addr_3279_6, addr_positional[52479:52476], addr_13119_7);

wire[31:0] addr_13120_7;

Selector_2 s13120_7(wires_3280_6[0], addr_3280_6, addr_positional[52483:52480], addr_13120_7);

wire[31:0] addr_13121_7;

Selector_2 s13121_7(wires_3280_6[1], addr_3280_6, addr_positional[52487:52484], addr_13121_7);

wire[31:0] addr_13122_7;

Selector_2 s13122_7(wires_3280_6[2], addr_3280_6, addr_positional[52491:52488], addr_13122_7);

wire[31:0] addr_13123_7;

Selector_2 s13123_7(wires_3280_6[3], addr_3280_6, addr_positional[52495:52492], addr_13123_7);

wire[31:0] addr_13124_7;

Selector_2 s13124_7(wires_3281_6[0], addr_3281_6, addr_positional[52499:52496], addr_13124_7);

wire[31:0] addr_13125_7;

Selector_2 s13125_7(wires_3281_6[1], addr_3281_6, addr_positional[52503:52500], addr_13125_7);

wire[31:0] addr_13126_7;

Selector_2 s13126_7(wires_3281_6[2], addr_3281_6, addr_positional[52507:52504], addr_13126_7);

wire[31:0] addr_13127_7;

Selector_2 s13127_7(wires_3281_6[3], addr_3281_6, addr_positional[52511:52508], addr_13127_7);

wire[31:0] addr_13128_7;

Selector_2 s13128_7(wires_3282_6[0], addr_3282_6, addr_positional[52515:52512], addr_13128_7);

wire[31:0] addr_13129_7;

Selector_2 s13129_7(wires_3282_6[1], addr_3282_6, addr_positional[52519:52516], addr_13129_7);

wire[31:0] addr_13130_7;

Selector_2 s13130_7(wires_3282_6[2], addr_3282_6, addr_positional[52523:52520], addr_13130_7);

wire[31:0] addr_13131_7;

Selector_2 s13131_7(wires_3282_6[3], addr_3282_6, addr_positional[52527:52524], addr_13131_7);

wire[31:0] addr_13132_7;

Selector_2 s13132_7(wires_3283_6[0], addr_3283_6, addr_positional[52531:52528], addr_13132_7);

wire[31:0] addr_13133_7;

Selector_2 s13133_7(wires_3283_6[1], addr_3283_6, addr_positional[52535:52532], addr_13133_7);

wire[31:0] addr_13134_7;

Selector_2 s13134_7(wires_3283_6[2], addr_3283_6, addr_positional[52539:52536], addr_13134_7);

wire[31:0] addr_13135_7;

Selector_2 s13135_7(wires_3283_6[3], addr_3283_6, addr_positional[52543:52540], addr_13135_7);

wire[31:0] addr_13136_7;

Selector_2 s13136_7(wires_3284_6[0], addr_3284_6, addr_positional[52547:52544], addr_13136_7);

wire[31:0] addr_13137_7;

Selector_2 s13137_7(wires_3284_6[1], addr_3284_6, addr_positional[52551:52548], addr_13137_7);

wire[31:0] addr_13138_7;

Selector_2 s13138_7(wires_3284_6[2], addr_3284_6, addr_positional[52555:52552], addr_13138_7);

wire[31:0] addr_13139_7;

Selector_2 s13139_7(wires_3284_6[3], addr_3284_6, addr_positional[52559:52556], addr_13139_7);

wire[31:0] addr_13140_7;

Selector_2 s13140_7(wires_3285_6[0], addr_3285_6, addr_positional[52563:52560], addr_13140_7);

wire[31:0] addr_13141_7;

Selector_2 s13141_7(wires_3285_6[1], addr_3285_6, addr_positional[52567:52564], addr_13141_7);

wire[31:0] addr_13142_7;

Selector_2 s13142_7(wires_3285_6[2], addr_3285_6, addr_positional[52571:52568], addr_13142_7);

wire[31:0] addr_13143_7;

Selector_2 s13143_7(wires_3285_6[3], addr_3285_6, addr_positional[52575:52572], addr_13143_7);

wire[31:0] addr_13144_7;

Selector_2 s13144_7(wires_3286_6[0], addr_3286_6, addr_positional[52579:52576], addr_13144_7);

wire[31:0] addr_13145_7;

Selector_2 s13145_7(wires_3286_6[1], addr_3286_6, addr_positional[52583:52580], addr_13145_7);

wire[31:0] addr_13146_7;

Selector_2 s13146_7(wires_3286_6[2], addr_3286_6, addr_positional[52587:52584], addr_13146_7);

wire[31:0] addr_13147_7;

Selector_2 s13147_7(wires_3286_6[3], addr_3286_6, addr_positional[52591:52588], addr_13147_7);

wire[31:0] addr_13148_7;

Selector_2 s13148_7(wires_3287_6[0], addr_3287_6, addr_positional[52595:52592], addr_13148_7);

wire[31:0] addr_13149_7;

Selector_2 s13149_7(wires_3287_6[1], addr_3287_6, addr_positional[52599:52596], addr_13149_7);

wire[31:0] addr_13150_7;

Selector_2 s13150_7(wires_3287_6[2], addr_3287_6, addr_positional[52603:52600], addr_13150_7);

wire[31:0] addr_13151_7;

Selector_2 s13151_7(wires_3287_6[3], addr_3287_6, addr_positional[52607:52604], addr_13151_7);

wire[31:0] addr_13152_7;

Selector_2 s13152_7(wires_3288_6[0], addr_3288_6, addr_positional[52611:52608], addr_13152_7);

wire[31:0] addr_13153_7;

Selector_2 s13153_7(wires_3288_6[1], addr_3288_6, addr_positional[52615:52612], addr_13153_7);

wire[31:0] addr_13154_7;

Selector_2 s13154_7(wires_3288_6[2], addr_3288_6, addr_positional[52619:52616], addr_13154_7);

wire[31:0] addr_13155_7;

Selector_2 s13155_7(wires_3288_6[3], addr_3288_6, addr_positional[52623:52620], addr_13155_7);

wire[31:0] addr_13156_7;

Selector_2 s13156_7(wires_3289_6[0], addr_3289_6, addr_positional[52627:52624], addr_13156_7);

wire[31:0] addr_13157_7;

Selector_2 s13157_7(wires_3289_6[1], addr_3289_6, addr_positional[52631:52628], addr_13157_7);

wire[31:0] addr_13158_7;

Selector_2 s13158_7(wires_3289_6[2], addr_3289_6, addr_positional[52635:52632], addr_13158_7);

wire[31:0] addr_13159_7;

Selector_2 s13159_7(wires_3289_6[3], addr_3289_6, addr_positional[52639:52636], addr_13159_7);

wire[31:0] addr_13160_7;

Selector_2 s13160_7(wires_3290_6[0], addr_3290_6, addr_positional[52643:52640], addr_13160_7);

wire[31:0] addr_13161_7;

Selector_2 s13161_7(wires_3290_6[1], addr_3290_6, addr_positional[52647:52644], addr_13161_7);

wire[31:0] addr_13162_7;

Selector_2 s13162_7(wires_3290_6[2], addr_3290_6, addr_positional[52651:52648], addr_13162_7);

wire[31:0] addr_13163_7;

Selector_2 s13163_7(wires_3290_6[3], addr_3290_6, addr_positional[52655:52652], addr_13163_7);

wire[31:0] addr_13164_7;

Selector_2 s13164_7(wires_3291_6[0], addr_3291_6, addr_positional[52659:52656], addr_13164_7);

wire[31:0] addr_13165_7;

Selector_2 s13165_7(wires_3291_6[1], addr_3291_6, addr_positional[52663:52660], addr_13165_7);

wire[31:0] addr_13166_7;

Selector_2 s13166_7(wires_3291_6[2], addr_3291_6, addr_positional[52667:52664], addr_13166_7);

wire[31:0] addr_13167_7;

Selector_2 s13167_7(wires_3291_6[3], addr_3291_6, addr_positional[52671:52668], addr_13167_7);

wire[31:0] addr_13168_7;

Selector_2 s13168_7(wires_3292_6[0], addr_3292_6, addr_positional[52675:52672], addr_13168_7);

wire[31:0] addr_13169_7;

Selector_2 s13169_7(wires_3292_6[1], addr_3292_6, addr_positional[52679:52676], addr_13169_7);

wire[31:0] addr_13170_7;

Selector_2 s13170_7(wires_3292_6[2], addr_3292_6, addr_positional[52683:52680], addr_13170_7);

wire[31:0] addr_13171_7;

Selector_2 s13171_7(wires_3292_6[3], addr_3292_6, addr_positional[52687:52684], addr_13171_7);

wire[31:0] addr_13172_7;

Selector_2 s13172_7(wires_3293_6[0], addr_3293_6, addr_positional[52691:52688], addr_13172_7);

wire[31:0] addr_13173_7;

Selector_2 s13173_7(wires_3293_6[1], addr_3293_6, addr_positional[52695:52692], addr_13173_7);

wire[31:0] addr_13174_7;

Selector_2 s13174_7(wires_3293_6[2], addr_3293_6, addr_positional[52699:52696], addr_13174_7);

wire[31:0] addr_13175_7;

Selector_2 s13175_7(wires_3293_6[3], addr_3293_6, addr_positional[52703:52700], addr_13175_7);

wire[31:0] addr_13176_7;

Selector_2 s13176_7(wires_3294_6[0], addr_3294_6, addr_positional[52707:52704], addr_13176_7);

wire[31:0] addr_13177_7;

Selector_2 s13177_7(wires_3294_6[1], addr_3294_6, addr_positional[52711:52708], addr_13177_7);

wire[31:0] addr_13178_7;

Selector_2 s13178_7(wires_3294_6[2], addr_3294_6, addr_positional[52715:52712], addr_13178_7);

wire[31:0] addr_13179_7;

Selector_2 s13179_7(wires_3294_6[3], addr_3294_6, addr_positional[52719:52716], addr_13179_7);

wire[31:0] addr_13180_7;

Selector_2 s13180_7(wires_3295_6[0], addr_3295_6, addr_positional[52723:52720], addr_13180_7);

wire[31:0] addr_13181_7;

Selector_2 s13181_7(wires_3295_6[1], addr_3295_6, addr_positional[52727:52724], addr_13181_7);

wire[31:0] addr_13182_7;

Selector_2 s13182_7(wires_3295_6[2], addr_3295_6, addr_positional[52731:52728], addr_13182_7);

wire[31:0] addr_13183_7;

Selector_2 s13183_7(wires_3295_6[3], addr_3295_6, addr_positional[52735:52732], addr_13183_7);

wire[31:0] addr_13184_7;

Selector_2 s13184_7(wires_3296_6[0], addr_3296_6, addr_positional[52739:52736], addr_13184_7);

wire[31:0] addr_13185_7;

Selector_2 s13185_7(wires_3296_6[1], addr_3296_6, addr_positional[52743:52740], addr_13185_7);

wire[31:0] addr_13186_7;

Selector_2 s13186_7(wires_3296_6[2], addr_3296_6, addr_positional[52747:52744], addr_13186_7);

wire[31:0] addr_13187_7;

Selector_2 s13187_7(wires_3296_6[3], addr_3296_6, addr_positional[52751:52748], addr_13187_7);

wire[31:0] addr_13188_7;

Selector_2 s13188_7(wires_3297_6[0], addr_3297_6, addr_positional[52755:52752], addr_13188_7);

wire[31:0] addr_13189_7;

Selector_2 s13189_7(wires_3297_6[1], addr_3297_6, addr_positional[52759:52756], addr_13189_7);

wire[31:0] addr_13190_7;

Selector_2 s13190_7(wires_3297_6[2], addr_3297_6, addr_positional[52763:52760], addr_13190_7);

wire[31:0] addr_13191_7;

Selector_2 s13191_7(wires_3297_6[3], addr_3297_6, addr_positional[52767:52764], addr_13191_7);

wire[31:0] addr_13192_7;

Selector_2 s13192_7(wires_3298_6[0], addr_3298_6, addr_positional[52771:52768], addr_13192_7);

wire[31:0] addr_13193_7;

Selector_2 s13193_7(wires_3298_6[1], addr_3298_6, addr_positional[52775:52772], addr_13193_7);

wire[31:0] addr_13194_7;

Selector_2 s13194_7(wires_3298_6[2], addr_3298_6, addr_positional[52779:52776], addr_13194_7);

wire[31:0] addr_13195_7;

Selector_2 s13195_7(wires_3298_6[3], addr_3298_6, addr_positional[52783:52780], addr_13195_7);

wire[31:0] addr_13196_7;

Selector_2 s13196_7(wires_3299_6[0], addr_3299_6, addr_positional[52787:52784], addr_13196_7);

wire[31:0] addr_13197_7;

Selector_2 s13197_7(wires_3299_6[1], addr_3299_6, addr_positional[52791:52788], addr_13197_7);

wire[31:0] addr_13198_7;

Selector_2 s13198_7(wires_3299_6[2], addr_3299_6, addr_positional[52795:52792], addr_13198_7);

wire[31:0] addr_13199_7;

Selector_2 s13199_7(wires_3299_6[3], addr_3299_6, addr_positional[52799:52796], addr_13199_7);

wire[31:0] addr_13200_7;

Selector_2 s13200_7(wires_3300_6[0], addr_3300_6, addr_positional[52803:52800], addr_13200_7);

wire[31:0] addr_13201_7;

Selector_2 s13201_7(wires_3300_6[1], addr_3300_6, addr_positional[52807:52804], addr_13201_7);

wire[31:0] addr_13202_7;

Selector_2 s13202_7(wires_3300_6[2], addr_3300_6, addr_positional[52811:52808], addr_13202_7);

wire[31:0] addr_13203_7;

Selector_2 s13203_7(wires_3300_6[3], addr_3300_6, addr_positional[52815:52812], addr_13203_7);

wire[31:0] addr_13204_7;

Selector_2 s13204_7(wires_3301_6[0], addr_3301_6, addr_positional[52819:52816], addr_13204_7);

wire[31:0] addr_13205_7;

Selector_2 s13205_7(wires_3301_6[1], addr_3301_6, addr_positional[52823:52820], addr_13205_7);

wire[31:0] addr_13206_7;

Selector_2 s13206_7(wires_3301_6[2], addr_3301_6, addr_positional[52827:52824], addr_13206_7);

wire[31:0] addr_13207_7;

Selector_2 s13207_7(wires_3301_6[3], addr_3301_6, addr_positional[52831:52828], addr_13207_7);

wire[31:0] addr_13208_7;

Selector_2 s13208_7(wires_3302_6[0], addr_3302_6, addr_positional[52835:52832], addr_13208_7);

wire[31:0] addr_13209_7;

Selector_2 s13209_7(wires_3302_6[1], addr_3302_6, addr_positional[52839:52836], addr_13209_7);

wire[31:0] addr_13210_7;

Selector_2 s13210_7(wires_3302_6[2], addr_3302_6, addr_positional[52843:52840], addr_13210_7);

wire[31:0] addr_13211_7;

Selector_2 s13211_7(wires_3302_6[3], addr_3302_6, addr_positional[52847:52844], addr_13211_7);

wire[31:0] addr_13212_7;

Selector_2 s13212_7(wires_3303_6[0], addr_3303_6, addr_positional[52851:52848], addr_13212_7);

wire[31:0] addr_13213_7;

Selector_2 s13213_7(wires_3303_6[1], addr_3303_6, addr_positional[52855:52852], addr_13213_7);

wire[31:0] addr_13214_7;

Selector_2 s13214_7(wires_3303_6[2], addr_3303_6, addr_positional[52859:52856], addr_13214_7);

wire[31:0] addr_13215_7;

Selector_2 s13215_7(wires_3303_6[3], addr_3303_6, addr_positional[52863:52860], addr_13215_7);

wire[31:0] addr_13216_7;

Selector_2 s13216_7(wires_3304_6[0], addr_3304_6, addr_positional[52867:52864], addr_13216_7);

wire[31:0] addr_13217_7;

Selector_2 s13217_7(wires_3304_6[1], addr_3304_6, addr_positional[52871:52868], addr_13217_7);

wire[31:0] addr_13218_7;

Selector_2 s13218_7(wires_3304_6[2], addr_3304_6, addr_positional[52875:52872], addr_13218_7);

wire[31:0] addr_13219_7;

Selector_2 s13219_7(wires_3304_6[3], addr_3304_6, addr_positional[52879:52876], addr_13219_7);

wire[31:0] addr_13220_7;

Selector_2 s13220_7(wires_3305_6[0], addr_3305_6, addr_positional[52883:52880], addr_13220_7);

wire[31:0] addr_13221_7;

Selector_2 s13221_7(wires_3305_6[1], addr_3305_6, addr_positional[52887:52884], addr_13221_7);

wire[31:0] addr_13222_7;

Selector_2 s13222_7(wires_3305_6[2], addr_3305_6, addr_positional[52891:52888], addr_13222_7);

wire[31:0] addr_13223_7;

Selector_2 s13223_7(wires_3305_6[3], addr_3305_6, addr_positional[52895:52892], addr_13223_7);

wire[31:0] addr_13224_7;

Selector_2 s13224_7(wires_3306_6[0], addr_3306_6, addr_positional[52899:52896], addr_13224_7);

wire[31:0] addr_13225_7;

Selector_2 s13225_7(wires_3306_6[1], addr_3306_6, addr_positional[52903:52900], addr_13225_7);

wire[31:0] addr_13226_7;

Selector_2 s13226_7(wires_3306_6[2], addr_3306_6, addr_positional[52907:52904], addr_13226_7);

wire[31:0] addr_13227_7;

Selector_2 s13227_7(wires_3306_6[3], addr_3306_6, addr_positional[52911:52908], addr_13227_7);

wire[31:0] addr_13228_7;

Selector_2 s13228_7(wires_3307_6[0], addr_3307_6, addr_positional[52915:52912], addr_13228_7);

wire[31:0] addr_13229_7;

Selector_2 s13229_7(wires_3307_6[1], addr_3307_6, addr_positional[52919:52916], addr_13229_7);

wire[31:0] addr_13230_7;

Selector_2 s13230_7(wires_3307_6[2], addr_3307_6, addr_positional[52923:52920], addr_13230_7);

wire[31:0] addr_13231_7;

Selector_2 s13231_7(wires_3307_6[3], addr_3307_6, addr_positional[52927:52924], addr_13231_7);

wire[31:0] addr_13232_7;

Selector_2 s13232_7(wires_3308_6[0], addr_3308_6, addr_positional[52931:52928], addr_13232_7);

wire[31:0] addr_13233_7;

Selector_2 s13233_7(wires_3308_6[1], addr_3308_6, addr_positional[52935:52932], addr_13233_7);

wire[31:0] addr_13234_7;

Selector_2 s13234_7(wires_3308_6[2], addr_3308_6, addr_positional[52939:52936], addr_13234_7);

wire[31:0] addr_13235_7;

Selector_2 s13235_7(wires_3308_6[3], addr_3308_6, addr_positional[52943:52940], addr_13235_7);

wire[31:0] addr_13236_7;

Selector_2 s13236_7(wires_3309_6[0], addr_3309_6, addr_positional[52947:52944], addr_13236_7);

wire[31:0] addr_13237_7;

Selector_2 s13237_7(wires_3309_6[1], addr_3309_6, addr_positional[52951:52948], addr_13237_7);

wire[31:0] addr_13238_7;

Selector_2 s13238_7(wires_3309_6[2], addr_3309_6, addr_positional[52955:52952], addr_13238_7);

wire[31:0] addr_13239_7;

Selector_2 s13239_7(wires_3309_6[3], addr_3309_6, addr_positional[52959:52956], addr_13239_7);

wire[31:0] addr_13240_7;

Selector_2 s13240_7(wires_3310_6[0], addr_3310_6, addr_positional[52963:52960], addr_13240_7);

wire[31:0] addr_13241_7;

Selector_2 s13241_7(wires_3310_6[1], addr_3310_6, addr_positional[52967:52964], addr_13241_7);

wire[31:0] addr_13242_7;

Selector_2 s13242_7(wires_3310_6[2], addr_3310_6, addr_positional[52971:52968], addr_13242_7);

wire[31:0] addr_13243_7;

Selector_2 s13243_7(wires_3310_6[3], addr_3310_6, addr_positional[52975:52972], addr_13243_7);

wire[31:0] addr_13244_7;

Selector_2 s13244_7(wires_3311_6[0], addr_3311_6, addr_positional[52979:52976], addr_13244_7);

wire[31:0] addr_13245_7;

Selector_2 s13245_7(wires_3311_6[1], addr_3311_6, addr_positional[52983:52980], addr_13245_7);

wire[31:0] addr_13246_7;

Selector_2 s13246_7(wires_3311_6[2], addr_3311_6, addr_positional[52987:52984], addr_13246_7);

wire[31:0] addr_13247_7;

Selector_2 s13247_7(wires_3311_6[3], addr_3311_6, addr_positional[52991:52988], addr_13247_7);

wire[31:0] addr_13248_7;

Selector_2 s13248_7(wires_3312_6[0], addr_3312_6, addr_positional[52995:52992], addr_13248_7);

wire[31:0] addr_13249_7;

Selector_2 s13249_7(wires_3312_6[1], addr_3312_6, addr_positional[52999:52996], addr_13249_7);

wire[31:0] addr_13250_7;

Selector_2 s13250_7(wires_3312_6[2], addr_3312_6, addr_positional[53003:53000], addr_13250_7);

wire[31:0] addr_13251_7;

Selector_2 s13251_7(wires_3312_6[3], addr_3312_6, addr_positional[53007:53004], addr_13251_7);

wire[31:0] addr_13252_7;

Selector_2 s13252_7(wires_3313_6[0], addr_3313_6, addr_positional[53011:53008], addr_13252_7);

wire[31:0] addr_13253_7;

Selector_2 s13253_7(wires_3313_6[1], addr_3313_6, addr_positional[53015:53012], addr_13253_7);

wire[31:0] addr_13254_7;

Selector_2 s13254_7(wires_3313_6[2], addr_3313_6, addr_positional[53019:53016], addr_13254_7);

wire[31:0] addr_13255_7;

Selector_2 s13255_7(wires_3313_6[3], addr_3313_6, addr_positional[53023:53020], addr_13255_7);

wire[31:0] addr_13256_7;

Selector_2 s13256_7(wires_3314_6[0], addr_3314_6, addr_positional[53027:53024], addr_13256_7);

wire[31:0] addr_13257_7;

Selector_2 s13257_7(wires_3314_6[1], addr_3314_6, addr_positional[53031:53028], addr_13257_7);

wire[31:0] addr_13258_7;

Selector_2 s13258_7(wires_3314_6[2], addr_3314_6, addr_positional[53035:53032], addr_13258_7);

wire[31:0] addr_13259_7;

Selector_2 s13259_7(wires_3314_6[3], addr_3314_6, addr_positional[53039:53036], addr_13259_7);

wire[31:0] addr_13260_7;

Selector_2 s13260_7(wires_3315_6[0], addr_3315_6, addr_positional[53043:53040], addr_13260_7);

wire[31:0] addr_13261_7;

Selector_2 s13261_7(wires_3315_6[1], addr_3315_6, addr_positional[53047:53044], addr_13261_7);

wire[31:0] addr_13262_7;

Selector_2 s13262_7(wires_3315_6[2], addr_3315_6, addr_positional[53051:53048], addr_13262_7);

wire[31:0] addr_13263_7;

Selector_2 s13263_7(wires_3315_6[3], addr_3315_6, addr_positional[53055:53052], addr_13263_7);

wire[31:0] addr_13264_7;

Selector_2 s13264_7(wires_3316_6[0], addr_3316_6, addr_positional[53059:53056], addr_13264_7);

wire[31:0] addr_13265_7;

Selector_2 s13265_7(wires_3316_6[1], addr_3316_6, addr_positional[53063:53060], addr_13265_7);

wire[31:0] addr_13266_7;

Selector_2 s13266_7(wires_3316_6[2], addr_3316_6, addr_positional[53067:53064], addr_13266_7);

wire[31:0] addr_13267_7;

Selector_2 s13267_7(wires_3316_6[3], addr_3316_6, addr_positional[53071:53068], addr_13267_7);

wire[31:0] addr_13268_7;

Selector_2 s13268_7(wires_3317_6[0], addr_3317_6, addr_positional[53075:53072], addr_13268_7);

wire[31:0] addr_13269_7;

Selector_2 s13269_7(wires_3317_6[1], addr_3317_6, addr_positional[53079:53076], addr_13269_7);

wire[31:0] addr_13270_7;

Selector_2 s13270_7(wires_3317_6[2], addr_3317_6, addr_positional[53083:53080], addr_13270_7);

wire[31:0] addr_13271_7;

Selector_2 s13271_7(wires_3317_6[3], addr_3317_6, addr_positional[53087:53084], addr_13271_7);

wire[31:0] addr_13272_7;

Selector_2 s13272_7(wires_3318_6[0], addr_3318_6, addr_positional[53091:53088], addr_13272_7);

wire[31:0] addr_13273_7;

Selector_2 s13273_7(wires_3318_6[1], addr_3318_6, addr_positional[53095:53092], addr_13273_7);

wire[31:0] addr_13274_7;

Selector_2 s13274_7(wires_3318_6[2], addr_3318_6, addr_positional[53099:53096], addr_13274_7);

wire[31:0] addr_13275_7;

Selector_2 s13275_7(wires_3318_6[3], addr_3318_6, addr_positional[53103:53100], addr_13275_7);

wire[31:0] addr_13276_7;

Selector_2 s13276_7(wires_3319_6[0], addr_3319_6, addr_positional[53107:53104], addr_13276_7);

wire[31:0] addr_13277_7;

Selector_2 s13277_7(wires_3319_6[1], addr_3319_6, addr_positional[53111:53108], addr_13277_7);

wire[31:0] addr_13278_7;

Selector_2 s13278_7(wires_3319_6[2], addr_3319_6, addr_positional[53115:53112], addr_13278_7);

wire[31:0] addr_13279_7;

Selector_2 s13279_7(wires_3319_6[3], addr_3319_6, addr_positional[53119:53116], addr_13279_7);

wire[31:0] addr_13280_7;

Selector_2 s13280_7(wires_3320_6[0], addr_3320_6, addr_positional[53123:53120], addr_13280_7);

wire[31:0] addr_13281_7;

Selector_2 s13281_7(wires_3320_6[1], addr_3320_6, addr_positional[53127:53124], addr_13281_7);

wire[31:0] addr_13282_7;

Selector_2 s13282_7(wires_3320_6[2], addr_3320_6, addr_positional[53131:53128], addr_13282_7);

wire[31:0] addr_13283_7;

Selector_2 s13283_7(wires_3320_6[3], addr_3320_6, addr_positional[53135:53132], addr_13283_7);

wire[31:0] addr_13284_7;

Selector_2 s13284_7(wires_3321_6[0], addr_3321_6, addr_positional[53139:53136], addr_13284_7);

wire[31:0] addr_13285_7;

Selector_2 s13285_7(wires_3321_6[1], addr_3321_6, addr_positional[53143:53140], addr_13285_7);

wire[31:0] addr_13286_7;

Selector_2 s13286_7(wires_3321_6[2], addr_3321_6, addr_positional[53147:53144], addr_13286_7);

wire[31:0] addr_13287_7;

Selector_2 s13287_7(wires_3321_6[3], addr_3321_6, addr_positional[53151:53148], addr_13287_7);

wire[31:0] addr_13288_7;

Selector_2 s13288_7(wires_3322_6[0], addr_3322_6, addr_positional[53155:53152], addr_13288_7);

wire[31:0] addr_13289_7;

Selector_2 s13289_7(wires_3322_6[1], addr_3322_6, addr_positional[53159:53156], addr_13289_7);

wire[31:0] addr_13290_7;

Selector_2 s13290_7(wires_3322_6[2], addr_3322_6, addr_positional[53163:53160], addr_13290_7);

wire[31:0] addr_13291_7;

Selector_2 s13291_7(wires_3322_6[3], addr_3322_6, addr_positional[53167:53164], addr_13291_7);

wire[31:0] addr_13292_7;

Selector_2 s13292_7(wires_3323_6[0], addr_3323_6, addr_positional[53171:53168], addr_13292_7);

wire[31:0] addr_13293_7;

Selector_2 s13293_7(wires_3323_6[1], addr_3323_6, addr_positional[53175:53172], addr_13293_7);

wire[31:0] addr_13294_7;

Selector_2 s13294_7(wires_3323_6[2], addr_3323_6, addr_positional[53179:53176], addr_13294_7);

wire[31:0] addr_13295_7;

Selector_2 s13295_7(wires_3323_6[3], addr_3323_6, addr_positional[53183:53180], addr_13295_7);

wire[31:0] addr_13296_7;

Selector_2 s13296_7(wires_3324_6[0], addr_3324_6, addr_positional[53187:53184], addr_13296_7);

wire[31:0] addr_13297_7;

Selector_2 s13297_7(wires_3324_6[1], addr_3324_6, addr_positional[53191:53188], addr_13297_7);

wire[31:0] addr_13298_7;

Selector_2 s13298_7(wires_3324_6[2], addr_3324_6, addr_positional[53195:53192], addr_13298_7);

wire[31:0] addr_13299_7;

Selector_2 s13299_7(wires_3324_6[3], addr_3324_6, addr_positional[53199:53196], addr_13299_7);

wire[31:0] addr_13300_7;

Selector_2 s13300_7(wires_3325_6[0], addr_3325_6, addr_positional[53203:53200], addr_13300_7);

wire[31:0] addr_13301_7;

Selector_2 s13301_7(wires_3325_6[1], addr_3325_6, addr_positional[53207:53204], addr_13301_7);

wire[31:0] addr_13302_7;

Selector_2 s13302_7(wires_3325_6[2], addr_3325_6, addr_positional[53211:53208], addr_13302_7);

wire[31:0] addr_13303_7;

Selector_2 s13303_7(wires_3325_6[3], addr_3325_6, addr_positional[53215:53212], addr_13303_7);

wire[31:0] addr_13304_7;

Selector_2 s13304_7(wires_3326_6[0], addr_3326_6, addr_positional[53219:53216], addr_13304_7);

wire[31:0] addr_13305_7;

Selector_2 s13305_7(wires_3326_6[1], addr_3326_6, addr_positional[53223:53220], addr_13305_7);

wire[31:0] addr_13306_7;

Selector_2 s13306_7(wires_3326_6[2], addr_3326_6, addr_positional[53227:53224], addr_13306_7);

wire[31:0] addr_13307_7;

Selector_2 s13307_7(wires_3326_6[3], addr_3326_6, addr_positional[53231:53228], addr_13307_7);

wire[31:0] addr_13308_7;

Selector_2 s13308_7(wires_3327_6[0], addr_3327_6, addr_positional[53235:53232], addr_13308_7);

wire[31:0] addr_13309_7;

Selector_2 s13309_7(wires_3327_6[1], addr_3327_6, addr_positional[53239:53236], addr_13309_7);

wire[31:0] addr_13310_7;

Selector_2 s13310_7(wires_3327_6[2], addr_3327_6, addr_positional[53243:53240], addr_13310_7);

wire[31:0] addr_13311_7;

Selector_2 s13311_7(wires_3327_6[3], addr_3327_6, addr_positional[53247:53244], addr_13311_7);

wire[31:0] addr_13312_7;

Selector_2 s13312_7(wires_3328_6[0], addr_3328_6, addr_positional[53251:53248], addr_13312_7);

wire[31:0] addr_13313_7;

Selector_2 s13313_7(wires_3328_6[1], addr_3328_6, addr_positional[53255:53252], addr_13313_7);

wire[31:0] addr_13314_7;

Selector_2 s13314_7(wires_3328_6[2], addr_3328_6, addr_positional[53259:53256], addr_13314_7);

wire[31:0] addr_13315_7;

Selector_2 s13315_7(wires_3328_6[3], addr_3328_6, addr_positional[53263:53260], addr_13315_7);

wire[31:0] addr_13316_7;

Selector_2 s13316_7(wires_3329_6[0], addr_3329_6, addr_positional[53267:53264], addr_13316_7);

wire[31:0] addr_13317_7;

Selector_2 s13317_7(wires_3329_6[1], addr_3329_6, addr_positional[53271:53268], addr_13317_7);

wire[31:0] addr_13318_7;

Selector_2 s13318_7(wires_3329_6[2], addr_3329_6, addr_positional[53275:53272], addr_13318_7);

wire[31:0] addr_13319_7;

Selector_2 s13319_7(wires_3329_6[3], addr_3329_6, addr_positional[53279:53276], addr_13319_7);

wire[31:0] addr_13320_7;

Selector_2 s13320_7(wires_3330_6[0], addr_3330_6, addr_positional[53283:53280], addr_13320_7);

wire[31:0] addr_13321_7;

Selector_2 s13321_7(wires_3330_6[1], addr_3330_6, addr_positional[53287:53284], addr_13321_7);

wire[31:0] addr_13322_7;

Selector_2 s13322_7(wires_3330_6[2], addr_3330_6, addr_positional[53291:53288], addr_13322_7);

wire[31:0] addr_13323_7;

Selector_2 s13323_7(wires_3330_6[3], addr_3330_6, addr_positional[53295:53292], addr_13323_7);

wire[31:0] addr_13324_7;

Selector_2 s13324_7(wires_3331_6[0], addr_3331_6, addr_positional[53299:53296], addr_13324_7);

wire[31:0] addr_13325_7;

Selector_2 s13325_7(wires_3331_6[1], addr_3331_6, addr_positional[53303:53300], addr_13325_7);

wire[31:0] addr_13326_7;

Selector_2 s13326_7(wires_3331_6[2], addr_3331_6, addr_positional[53307:53304], addr_13326_7);

wire[31:0] addr_13327_7;

Selector_2 s13327_7(wires_3331_6[3], addr_3331_6, addr_positional[53311:53308], addr_13327_7);

wire[31:0] addr_13328_7;

Selector_2 s13328_7(wires_3332_6[0], addr_3332_6, addr_positional[53315:53312], addr_13328_7);

wire[31:0] addr_13329_7;

Selector_2 s13329_7(wires_3332_6[1], addr_3332_6, addr_positional[53319:53316], addr_13329_7);

wire[31:0] addr_13330_7;

Selector_2 s13330_7(wires_3332_6[2], addr_3332_6, addr_positional[53323:53320], addr_13330_7);

wire[31:0] addr_13331_7;

Selector_2 s13331_7(wires_3332_6[3], addr_3332_6, addr_positional[53327:53324], addr_13331_7);

wire[31:0] addr_13332_7;

Selector_2 s13332_7(wires_3333_6[0], addr_3333_6, addr_positional[53331:53328], addr_13332_7);

wire[31:0] addr_13333_7;

Selector_2 s13333_7(wires_3333_6[1], addr_3333_6, addr_positional[53335:53332], addr_13333_7);

wire[31:0] addr_13334_7;

Selector_2 s13334_7(wires_3333_6[2], addr_3333_6, addr_positional[53339:53336], addr_13334_7);

wire[31:0] addr_13335_7;

Selector_2 s13335_7(wires_3333_6[3], addr_3333_6, addr_positional[53343:53340], addr_13335_7);

wire[31:0] addr_13336_7;

Selector_2 s13336_7(wires_3334_6[0], addr_3334_6, addr_positional[53347:53344], addr_13336_7);

wire[31:0] addr_13337_7;

Selector_2 s13337_7(wires_3334_6[1], addr_3334_6, addr_positional[53351:53348], addr_13337_7);

wire[31:0] addr_13338_7;

Selector_2 s13338_7(wires_3334_6[2], addr_3334_6, addr_positional[53355:53352], addr_13338_7);

wire[31:0] addr_13339_7;

Selector_2 s13339_7(wires_3334_6[3], addr_3334_6, addr_positional[53359:53356], addr_13339_7);

wire[31:0] addr_13340_7;

Selector_2 s13340_7(wires_3335_6[0], addr_3335_6, addr_positional[53363:53360], addr_13340_7);

wire[31:0] addr_13341_7;

Selector_2 s13341_7(wires_3335_6[1], addr_3335_6, addr_positional[53367:53364], addr_13341_7);

wire[31:0] addr_13342_7;

Selector_2 s13342_7(wires_3335_6[2], addr_3335_6, addr_positional[53371:53368], addr_13342_7);

wire[31:0] addr_13343_7;

Selector_2 s13343_7(wires_3335_6[3], addr_3335_6, addr_positional[53375:53372], addr_13343_7);

wire[31:0] addr_13344_7;

Selector_2 s13344_7(wires_3336_6[0], addr_3336_6, addr_positional[53379:53376], addr_13344_7);

wire[31:0] addr_13345_7;

Selector_2 s13345_7(wires_3336_6[1], addr_3336_6, addr_positional[53383:53380], addr_13345_7);

wire[31:0] addr_13346_7;

Selector_2 s13346_7(wires_3336_6[2], addr_3336_6, addr_positional[53387:53384], addr_13346_7);

wire[31:0] addr_13347_7;

Selector_2 s13347_7(wires_3336_6[3], addr_3336_6, addr_positional[53391:53388], addr_13347_7);

wire[31:0] addr_13348_7;

Selector_2 s13348_7(wires_3337_6[0], addr_3337_6, addr_positional[53395:53392], addr_13348_7);

wire[31:0] addr_13349_7;

Selector_2 s13349_7(wires_3337_6[1], addr_3337_6, addr_positional[53399:53396], addr_13349_7);

wire[31:0] addr_13350_7;

Selector_2 s13350_7(wires_3337_6[2], addr_3337_6, addr_positional[53403:53400], addr_13350_7);

wire[31:0] addr_13351_7;

Selector_2 s13351_7(wires_3337_6[3], addr_3337_6, addr_positional[53407:53404], addr_13351_7);

wire[31:0] addr_13352_7;

Selector_2 s13352_7(wires_3338_6[0], addr_3338_6, addr_positional[53411:53408], addr_13352_7);

wire[31:0] addr_13353_7;

Selector_2 s13353_7(wires_3338_6[1], addr_3338_6, addr_positional[53415:53412], addr_13353_7);

wire[31:0] addr_13354_7;

Selector_2 s13354_7(wires_3338_6[2], addr_3338_6, addr_positional[53419:53416], addr_13354_7);

wire[31:0] addr_13355_7;

Selector_2 s13355_7(wires_3338_6[3], addr_3338_6, addr_positional[53423:53420], addr_13355_7);

wire[31:0] addr_13356_7;

Selector_2 s13356_7(wires_3339_6[0], addr_3339_6, addr_positional[53427:53424], addr_13356_7);

wire[31:0] addr_13357_7;

Selector_2 s13357_7(wires_3339_6[1], addr_3339_6, addr_positional[53431:53428], addr_13357_7);

wire[31:0] addr_13358_7;

Selector_2 s13358_7(wires_3339_6[2], addr_3339_6, addr_positional[53435:53432], addr_13358_7);

wire[31:0] addr_13359_7;

Selector_2 s13359_7(wires_3339_6[3], addr_3339_6, addr_positional[53439:53436], addr_13359_7);

wire[31:0] addr_13360_7;

Selector_2 s13360_7(wires_3340_6[0], addr_3340_6, addr_positional[53443:53440], addr_13360_7);

wire[31:0] addr_13361_7;

Selector_2 s13361_7(wires_3340_6[1], addr_3340_6, addr_positional[53447:53444], addr_13361_7);

wire[31:0] addr_13362_7;

Selector_2 s13362_7(wires_3340_6[2], addr_3340_6, addr_positional[53451:53448], addr_13362_7);

wire[31:0] addr_13363_7;

Selector_2 s13363_7(wires_3340_6[3], addr_3340_6, addr_positional[53455:53452], addr_13363_7);

wire[31:0] addr_13364_7;

Selector_2 s13364_7(wires_3341_6[0], addr_3341_6, addr_positional[53459:53456], addr_13364_7);

wire[31:0] addr_13365_7;

Selector_2 s13365_7(wires_3341_6[1], addr_3341_6, addr_positional[53463:53460], addr_13365_7);

wire[31:0] addr_13366_7;

Selector_2 s13366_7(wires_3341_6[2], addr_3341_6, addr_positional[53467:53464], addr_13366_7);

wire[31:0] addr_13367_7;

Selector_2 s13367_7(wires_3341_6[3], addr_3341_6, addr_positional[53471:53468], addr_13367_7);

wire[31:0] addr_13368_7;

Selector_2 s13368_7(wires_3342_6[0], addr_3342_6, addr_positional[53475:53472], addr_13368_7);

wire[31:0] addr_13369_7;

Selector_2 s13369_7(wires_3342_6[1], addr_3342_6, addr_positional[53479:53476], addr_13369_7);

wire[31:0] addr_13370_7;

Selector_2 s13370_7(wires_3342_6[2], addr_3342_6, addr_positional[53483:53480], addr_13370_7);

wire[31:0] addr_13371_7;

Selector_2 s13371_7(wires_3342_6[3], addr_3342_6, addr_positional[53487:53484], addr_13371_7);

wire[31:0] addr_13372_7;

Selector_2 s13372_7(wires_3343_6[0], addr_3343_6, addr_positional[53491:53488], addr_13372_7);

wire[31:0] addr_13373_7;

Selector_2 s13373_7(wires_3343_6[1], addr_3343_6, addr_positional[53495:53492], addr_13373_7);

wire[31:0] addr_13374_7;

Selector_2 s13374_7(wires_3343_6[2], addr_3343_6, addr_positional[53499:53496], addr_13374_7);

wire[31:0] addr_13375_7;

Selector_2 s13375_7(wires_3343_6[3], addr_3343_6, addr_positional[53503:53500], addr_13375_7);

wire[31:0] addr_13376_7;

Selector_2 s13376_7(wires_3344_6[0], addr_3344_6, addr_positional[53507:53504], addr_13376_7);

wire[31:0] addr_13377_7;

Selector_2 s13377_7(wires_3344_6[1], addr_3344_6, addr_positional[53511:53508], addr_13377_7);

wire[31:0] addr_13378_7;

Selector_2 s13378_7(wires_3344_6[2], addr_3344_6, addr_positional[53515:53512], addr_13378_7);

wire[31:0] addr_13379_7;

Selector_2 s13379_7(wires_3344_6[3], addr_3344_6, addr_positional[53519:53516], addr_13379_7);

wire[31:0] addr_13380_7;

Selector_2 s13380_7(wires_3345_6[0], addr_3345_6, addr_positional[53523:53520], addr_13380_7);

wire[31:0] addr_13381_7;

Selector_2 s13381_7(wires_3345_6[1], addr_3345_6, addr_positional[53527:53524], addr_13381_7);

wire[31:0] addr_13382_7;

Selector_2 s13382_7(wires_3345_6[2], addr_3345_6, addr_positional[53531:53528], addr_13382_7);

wire[31:0] addr_13383_7;

Selector_2 s13383_7(wires_3345_6[3], addr_3345_6, addr_positional[53535:53532], addr_13383_7);

wire[31:0] addr_13384_7;

Selector_2 s13384_7(wires_3346_6[0], addr_3346_6, addr_positional[53539:53536], addr_13384_7);

wire[31:0] addr_13385_7;

Selector_2 s13385_7(wires_3346_6[1], addr_3346_6, addr_positional[53543:53540], addr_13385_7);

wire[31:0] addr_13386_7;

Selector_2 s13386_7(wires_3346_6[2], addr_3346_6, addr_positional[53547:53544], addr_13386_7);

wire[31:0] addr_13387_7;

Selector_2 s13387_7(wires_3346_6[3], addr_3346_6, addr_positional[53551:53548], addr_13387_7);

wire[31:0] addr_13388_7;

Selector_2 s13388_7(wires_3347_6[0], addr_3347_6, addr_positional[53555:53552], addr_13388_7);

wire[31:0] addr_13389_7;

Selector_2 s13389_7(wires_3347_6[1], addr_3347_6, addr_positional[53559:53556], addr_13389_7);

wire[31:0] addr_13390_7;

Selector_2 s13390_7(wires_3347_6[2], addr_3347_6, addr_positional[53563:53560], addr_13390_7);

wire[31:0] addr_13391_7;

Selector_2 s13391_7(wires_3347_6[3], addr_3347_6, addr_positional[53567:53564], addr_13391_7);

wire[31:0] addr_13392_7;

Selector_2 s13392_7(wires_3348_6[0], addr_3348_6, addr_positional[53571:53568], addr_13392_7);

wire[31:0] addr_13393_7;

Selector_2 s13393_7(wires_3348_6[1], addr_3348_6, addr_positional[53575:53572], addr_13393_7);

wire[31:0] addr_13394_7;

Selector_2 s13394_7(wires_3348_6[2], addr_3348_6, addr_positional[53579:53576], addr_13394_7);

wire[31:0] addr_13395_7;

Selector_2 s13395_7(wires_3348_6[3], addr_3348_6, addr_positional[53583:53580], addr_13395_7);

wire[31:0] addr_13396_7;

Selector_2 s13396_7(wires_3349_6[0], addr_3349_6, addr_positional[53587:53584], addr_13396_7);

wire[31:0] addr_13397_7;

Selector_2 s13397_7(wires_3349_6[1], addr_3349_6, addr_positional[53591:53588], addr_13397_7);

wire[31:0] addr_13398_7;

Selector_2 s13398_7(wires_3349_6[2], addr_3349_6, addr_positional[53595:53592], addr_13398_7);

wire[31:0] addr_13399_7;

Selector_2 s13399_7(wires_3349_6[3], addr_3349_6, addr_positional[53599:53596], addr_13399_7);

wire[31:0] addr_13400_7;

Selector_2 s13400_7(wires_3350_6[0], addr_3350_6, addr_positional[53603:53600], addr_13400_7);

wire[31:0] addr_13401_7;

Selector_2 s13401_7(wires_3350_6[1], addr_3350_6, addr_positional[53607:53604], addr_13401_7);

wire[31:0] addr_13402_7;

Selector_2 s13402_7(wires_3350_6[2], addr_3350_6, addr_positional[53611:53608], addr_13402_7);

wire[31:0] addr_13403_7;

Selector_2 s13403_7(wires_3350_6[3], addr_3350_6, addr_positional[53615:53612], addr_13403_7);

wire[31:0] addr_13404_7;

Selector_2 s13404_7(wires_3351_6[0], addr_3351_6, addr_positional[53619:53616], addr_13404_7);

wire[31:0] addr_13405_7;

Selector_2 s13405_7(wires_3351_6[1], addr_3351_6, addr_positional[53623:53620], addr_13405_7);

wire[31:0] addr_13406_7;

Selector_2 s13406_7(wires_3351_6[2], addr_3351_6, addr_positional[53627:53624], addr_13406_7);

wire[31:0] addr_13407_7;

Selector_2 s13407_7(wires_3351_6[3], addr_3351_6, addr_positional[53631:53628], addr_13407_7);

wire[31:0] addr_13408_7;

Selector_2 s13408_7(wires_3352_6[0], addr_3352_6, addr_positional[53635:53632], addr_13408_7);

wire[31:0] addr_13409_7;

Selector_2 s13409_7(wires_3352_6[1], addr_3352_6, addr_positional[53639:53636], addr_13409_7);

wire[31:0] addr_13410_7;

Selector_2 s13410_7(wires_3352_6[2], addr_3352_6, addr_positional[53643:53640], addr_13410_7);

wire[31:0] addr_13411_7;

Selector_2 s13411_7(wires_3352_6[3], addr_3352_6, addr_positional[53647:53644], addr_13411_7);

wire[31:0] addr_13412_7;

Selector_2 s13412_7(wires_3353_6[0], addr_3353_6, addr_positional[53651:53648], addr_13412_7);

wire[31:0] addr_13413_7;

Selector_2 s13413_7(wires_3353_6[1], addr_3353_6, addr_positional[53655:53652], addr_13413_7);

wire[31:0] addr_13414_7;

Selector_2 s13414_7(wires_3353_6[2], addr_3353_6, addr_positional[53659:53656], addr_13414_7);

wire[31:0] addr_13415_7;

Selector_2 s13415_7(wires_3353_6[3], addr_3353_6, addr_positional[53663:53660], addr_13415_7);

wire[31:0] addr_13416_7;

Selector_2 s13416_7(wires_3354_6[0], addr_3354_6, addr_positional[53667:53664], addr_13416_7);

wire[31:0] addr_13417_7;

Selector_2 s13417_7(wires_3354_6[1], addr_3354_6, addr_positional[53671:53668], addr_13417_7);

wire[31:0] addr_13418_7;

Selector_2 s13418_7(wires_3354_6[2], addr_3354_6, addr_positional[53675:53672], addr_13418_7);

wire[31:0] addr_13419_7;

Selector_2 s13419_7(wires_3354_6[3], addr_3354_6, addr_positional[53679:53676], addr_13419_7);

wire[31:0] addr_13420_7;

Selector_2 s13420_7(wires_3355_6[0], addr_3355_6, addr_positional[53683:53680], addr_13420_7);

wire[31:0] addr_13421_7;

Selector_2 s13421_7(wires_3355_6[1], addr_3355_6, addr_positional[53687:53684], addr_13421_7);

wire[31:0] addr_13422_7;

Selector_2 s13422_7(wires_3355_6[2], addr_3355_6, addr_positional[53691:53688], addr_13422_7);

wire[31:0] addr_13423_7;

Selector_2 s13423_7(wires_3355_6[3], addr_3355_6, addr_positional[53695:53692], addr_13423_7);

wire[31:0] addr_13424_7;

Selector_2 s13424_7(wires_3356_6[0], addr_3356_6, addr_positional[53699:53696], addr_13424_7);

wire[31:0] addr_13425_7;

Selector_2 s13425_7(wires_3356_6[1], addr_3356_6, addr_positional[53703:53700], addr_13425_7);

wire[31:0] addr_13426_7;

Selector_2 s13426_7(wires_3356_6[2], addr_3356_6, addr_positional[53707:53704], addr_13426_7);

wire[31:0] addr_13427_7;

Selector_2 s13427_7(wires_3356_6[3], addr_3356_6, addr_positional[53711:53708], addr_13427_7);

wire[31:0] addr_13428_7;

Selector_2 s13428_7(wires_3357_6[0], addr_3357_6, addr_positional[53715:53712], addr_13428_7);

wire[31:0] addr_13429_7;

Selector_2 s13429_7(wires_3357_6[1], addr_3357_6, addr_positional[53719:53716], addr_13429_7);

wire[31:0] addr_13430_7;

Selector_2 s13430_7(wires_3357_6[2], addr_3357_6, addr_positional[53723:53720], addr_13430_7);

wire[31:0] addr_13431_7;

Selector_2 s13431_7(wires_3357_6[3], addr_3357_6, addr_positional[53727:53724], addr_13431_7);

wire[31:0] addr_13432_7;

Selector_2 s13432_7(wires_3358_6[0], addr_3358_6, addr_positional[53731:53728], addr_13432_7);

wire[31:0] addr_13433_7;

Selector_2 s13433_7(wires_3358_6[1], addr_3358_6, addr_positional[53735:53732], addr_13433_7);

wire[31:0] addr_13434_7;

Selector_2 s13434_7(wires_3358_6[2], addr_3358_6, addr_positional[53739:53736], addr_13434_7);

wire[31:0] addr_13435_7;

Selector_2 s13435_7(wires_3358_6[3], addr_3358_6, addr_positional[53743:53740], addr_13435_7);

wire[31:0] addr_13436_7;

Selector_2 s13436_7(wires_3359_6[0], addr_3359_6, addr_positional[53747:53744], addr_13436_7);

wire[31:0] addr_13437_7;

Selector_2 s13437_7(wires_3359_6[1], addr_3359_6, addr_positional[53751:53748], addr_13437_7);

wire[31:0] addr_13438_7;

Selector_2 s13438_7(wires_3359_6[2], addr_3359_6, addr_positional[53755:53752], addr_13438_7);

wire[31:0] addr_13439_7;

Selector_2 s13439_7(wires_3359_6[3], addr_3359_6, addr_positional[53759:53756], addr_13439_7);

wire[31:0] addr_13440_7;

Selector_2 s13440_7(wires_3360_6[0], addr_3360_6, addr_positional[53763:53760], addr_13440_7);

wire[31:0] addr_13441_7;

Selector_2 s13441_7(wires_3360_6[1], addr_3360_6, addr_positional[53767:53764], addr_13441_7);

wire[31:0] addr_13442_7;

Selector_2 s13442_7(wires_3360_6[2], addr_3360_6, addr_positional[53771:53768], addr_13442_7);

wire[31:0] addr_13443_7;

Selector_2 s13443_7(wires_3360_6[3], addr_3360_6, addr_positional[53775:53772], addr_13443_7);

wire[31:0] addr_13444_7;

Selector_2 s13444_7(wires_3361_6[0], addr_3361_6, addr_positional[53779:53776], addr_13444_7);

wire[31:0] addr_13445_7;

Selector_2 s13445_7(wires_3361_6[1], addr_3361_6, addr_positional[53783:53780], addr_13445_7);

wire[31:0] addr_13446_7;

Selector_2 s13446_7(wires_3361_6[2], addr_3361_6, addr_positional[53787:53784], addr_13446_7);

wire[31:0] addr_13447_7;

Selector_2 s13447_7(wires_3361_6[3], addr_3361_6, addr_positional[53791:53788], addr_13447_7);

wire[31:0] addr_13448_7;

Selector_2 s13448_7(wires_3362_6[0], addr_3362_6, addr_positional[53795:53792], addr_13448_7);

wire[31:0] addr_13449_7;

Selector_2 s13449_7(wires_3362_6[1], addr_3362_6, addr_positional[53799:53796], addr_13449_7);

wire[31:0] addr_13450_7;

Selector_2 s13450_7(wires_3362_6[2], addr_3362_6, addr_positional[53803:53800], addr_13450_7);

wire[31:0] addr_13451_7;

Selector_2 s13451_7(wires_3362_6[3], addr_3362_6, addr_positional[53807:53804], addr_13451_7);

wire[31:0] addr_13452_7;

Selector_2 s13452_7(wires_3363_6[0], addr_3363_6, addr_positional[53811:53808], addr_13452_7);

wire[31:0] addr_13453_7;

Selector_2 s13453_7(wires_3363_6[1], addr_3363_6, addr_positional[53815:53812], addr_13453_7);

wire[31:0] addr_13454_7;

Selector_2 s13454_7(wires_3363_6[2], addr_3363_6, addr_positional[53819:53816], addr_13454_7);

wire[31:0] addr_13455_7;

Selector_2 s13455_7(wires_3363_6[3], addr_3363_6, addr_positional[53823:53820], addr_13455_7);

wire[31:0] addr_13456_7;

Selector_2 s13456_7(wires_3364_6[0], addr_3364_6, addr_positional[53827:53824], addr_13456_7);

wire[31:0] addr_13457_7;

Selector_2 s13457_7(wires_3364_6[1], addr_3364_6, addr_positional[53831:53828], addr_13457_7);

wire[31:0] addr_13458_7;

Selector_2 s13458_7(wires_3364_6[2], addr_3364_6, addr_positional[53835:53832], addr_13458_7);

wire[31:0] addr_13459_7;

Selector_2 s13459_7(wires_3364_6[3], addr_3364_6, addr_positional[53839:53836], addr_13459_7);

wire[31:0] addr_13460_7;

Selector_2 s13460_7(wires_3365_6[0], addr_3365_6, addr_positional[53843:53840], addr_13460_7);

wire[31:0] addr_13461_7;

Selector_2 s13461_7(wires_3365_6[1], addr_3365_6, addr_positional[53847:53844], addr_13461_7);

wire[31:0] addr_13462_7;

Selector_2 s13462_7(wires_3365_6[2], addr_3365_6, addr_positional[53851:53848], addr_13462_7);

wire[31:0] addr_13463_7;

Selector_2 s13463_7(wires_3365_6[3], addr_3365_6, addr_positional[53855:53852], addr_13463_7);

wire[31:0] addr_13464_7;

Selector_2 s13464_7(wires_3366_6[0], addr_3366_6, addr_positional[53859:53856], addr_13464_7);

wire[31:0] addr_13465_7;

Selector_2 s13465_7(wires_3366_6[1], addr_3366_6, addr_positional[53863:53860], addr_13465_7);

wire[31:0] addr_13466_7;

Selector_2 s13466_7(wires_3366_6[2], addr_3366_6, addr_positional[53867:53864], addr_13466_7);

wire[31:0] addr_13467_7;

Selector_2 s13467_7(wires_3366_6[3], addr_3366_6, addr_positional[53871:53868], addr_13467_7);

wire[31:0] addr_13468_7;

Selector_2 s13468_7(wires_3367_6[0], addr_3367_6, addr_positional[53875:53872], addr_13468_7);

wire[31:0] addr_13469_7;

Selector_2 s13469_7(wires_3367_6[1], addr_3367_6, addr_positional[53879:53876], addr_13469_7);

wire[31:0] addr_13470_7;

Selector_2 s13470_7(wires_3367_6[2], addr_3367_6, addr_positional[53883:53880], addr_13470_7);

wire[31:0] addr_13471_7;

Selector_2 s13471_7(wires_3367_6[3], addr_3367_6, addr_positional[53887:53884], addr_13471_7);

wire[31:0] addr_13472_7;

Selector_2 s13472_7(wires_3368_6[0], addr_3368_6, addr_positional[53891:53888], addr_13472_7);

wire[31:0] addr_13473_7;

Selector_2 s13473_7(wires_3368_6[1], addr_3368_6, addr_positional[53895:53892], addr_13473_7);

wire[31:0] addr_13474_7;

Selector_2 s13474_7(wires_3368_6[2], addr_3368_6, addr_positional[53899:53896], addr_13474_7);

wire[31:0] addr_13475_7;

Selector_2 s13475_7(wires_3368_6[3], addr_3368_6, addr_positional[53903:53900], addr_13475_7);

wire[31:0] addr_13476_7;

Selector_2 s13476_7(wires_3369_6[0], addr_3369_6, addr_positional[53907:53904], addr_13476_7);

wire[31:0] addr_13477_7;

Selector_2 s13477_7(wires_3369_6[1], addr_3369_6, addr_positional[53911:53908], addr_13477_7);

wire[31:0] addr_13478_7;

Selector_2 s13478_7(wires_3369_6[2], addr_3369_6, addr_positional[53915:53912], addr_13478_7);

wire[31:0] addr_13479_7;

Selector_2 s13479_7(wires_3369_6[3], addr_3369_6, addr_positional[53919:53916], addr_13479_7);

wire[31:0] addr_13480_7;

Selector_2 s13480_7(wires_3370_6[0], addr_3370_6, addr_positional[53923:53920], addr_13480_7);

wire[31:0] addr_13481_7;

Selector_2 s13481_7(wires_3370_6[1], addr_3370_6, addr_positional[53927:53924], addr_13481_7);

wire[31:0] addr_13482_7;

Selector_2 s13482_7(wires_3370_6[2], addr_3370_6, addr_positional[53931:53928], addr_13482_7);

wire[31:0] addr_13483_7;

Selector_2 s13483_7(wires_3370_6[3], addr_3370_6, addr_positional[53935:53932], addr_13483_7);

wire[31:0] addr_13484_7;

Selector_2 s13484_7(wires_3371_6[0], addr_3371_6, addr_positional[53939:53936], addr_13484_7);

wire[31:0] addr_13485_7;

Selector_2 s13485_7(wires_3371_6[1], addr_3371_6, addr_positional[53943:53940], addr_13485_7);

wire[31:0] addr_13486_7;

Selector_2 s13486_7(wires_3371_6[2], addr_3371_6, addr_positional[53947:53944], addr_13486_7);

wire[31:0] addr_13487_7;

Selector_2 s13487_7(wires_3371_6[3], addr_3371_6, addr_positional[53951:53948], addr_13487_7);

wire[31:0] addr_13488_7;

Selector_2 s13488_7(wires_3372_6[0], addr_3372_6, addr_positional[53955:53952], addr_13488_7);

wire[31:0] addr_13489_7;

Selector_2 s13489_7(wires_3372_6[1], addr_3372_6, addr_positional[53959:53956], addr_13489_7);

wire[31:0] addr_13490_7;

Selector_2 s13490_7(wires_3372_6[2], addr_3372_6, addr_positional[53963:53960], addr_13490_7);

wire[31:0] addr_13491_7;

Selector_2 s13491_7(wires_3372_6[3], addr_3372_6, addr_positional[53967:53964], addr_13491_7);

wire[31:0] addr_13492_7;

Selector_2 s13492_7(wires_3373_6[0], addr_3373_6, addr_positional[53971:53968], addr_13492_7);

wire[31:0] addr_13493_7;

Selector_2 s13493_7(wires_3373_6[1], addr_3373_6, addr_positional[53975:53972], addr_13493_7);

wire[31:0] addr_13494_7;

Selector_2 s13494_7(wires_3373_6[2], addr_3373_6, addr_positional[53979:53976], addr_13494_7);

wire[31:0] addr_13495_7;

Selector_2 s13495_7(wires_3373_6[3], addr_3373_6, addr_positional[53983:53980], addr_13495_7);

wire[31:0] addr_13496_7;

Selector_2 s13496_7(wires_3374_6[0], addr_3374_6, addr_positional[53987:53984], addr_13496_7);

wire[31:0] addr_13497_7;

Selector_2 s13497_7(wires_3374_6[1], addr_3374_6, addr_positional[53991:53988], addr_13497_7);

wire[31:0] addr_13498_7;

Selector_2 s13498_7(wires_3374_6[2], addr_3374_6, addr_positional[53995:53992], addr_13498_7);

wire[31:0] addr_13499_7;

Selector_2 s13499_7(wires_3374_6[3], addr_3374_6, addr_positional[53999:53996], addr_13499_7);

wire[31:0] addr_13500_7;

Selector_2 s13500_7(wires_3375_6[0], addr_3375_6, addr_positional[54003:54000], addr_13500_7);

wire[31:0] addr_13501_7;

Selector_2 s13501_7(wires_3375_6[1], addr_3375_6, addr_positional[54007:54004], addr_13501_7);

wire[31:0] addr_13502_7;

Selector_2 s13502_7(wires_3375_6[2], addr_3375_6, addr_positional[54011:54008], addr_13502_7);

wire[31:0] addr_13503_7;

Selector_2 s13503_7(wires_3375_6[3], addr_3375_6, addr_positional[54015:54012], addr_13503_7);

wire[31:0] addr_13504_7;

Selector_2 s13504_7(wires_3376_6[0], addr_3376_6, addr_positional[54019:54016], addr_13504_7);

wire[31:0] addr_13505_7;

Selector_2 s13505_7(wires_3376_6[1], addr_3376_6, addr_positional[54023:54020], addr_13505_7);

wire[31:0] addr_13506_7;

Selector_2 s13506_7(wires_3376_6[2], addr_3376_6, addr_positional[54027:54024], addr_13506_7);

wire[31:0] addr_13507_7;

Selector_2 s13507_7(wires_3376_6[3], addr_3376_6, addr_positional[54031:54028], addr_13507_7);

wire[31:0] addr_13508_7;

Selector_2 s13508_7(wires_3377_6[0], addr_3377_6, addr_positional[54035:54032], addr_13508_7);

wire[31:0] addr_13509_7;

Selector_2 s13509_7(wires_3377_6[1], addr_3377_6, addr_positional[54039:54036], addr_13509_7);

wire[31:0] addr_13510_7;

Selector_2 s13510_7(wires_3377_6[2], addr_3377_6, addr_positional[54043:54040], addr_13510_7);

wire[31:0] addr_13511_7;

Selector_2 s13511_7(wires_3377_6[3], addr_3377_6, addr_positional[54047:54044], addr_13511_7);

wire[31:0] addr_13512_7;

Selector_2 s13512_7(wires_3378_6[0], addr_3378_6, addr_positional[54051:54048], addr_13512_7);

wire[31:0] addr_13513_7;

Selector_2 s13513_7(wires_3378_6[1], addr_3378_6, addr_positional[54055:54052], addr_13513_7);

wire[31:0] addr_13514_7;

Selector_2 s13514_7(wires_3378_6[2], addr_3378_6, addr_positional[54059:54056], addr_13514_7);

wire[31:0] addr_13515_7;

Selector_2 s13515_7(wires_3378_6[3], addr_3378_6, addr_positional[54063:54060], addr_13515_7);

wire[31:0] addr_13516_7;

Selector_2 s13516_7(wires_3379_6[0], addr_3379_6, addr_positional[54067:54064], addr_13516_7);

wire[31:0] addr_13517_7;

Selector_2 s13517_7(wires_3379_6[1], addr_3379_6, addr_positional[54071:54068], addr_13517_7);

wire[31:0] addr_13518_7;

Selector_2 s13518_7(wires_3379_6[2], addr_3379_6, addr_positional[54075:54072], addr_13518_7);

wire[31:0] addr_13519_7;

Selector_2 s13519_7(wires_3379_6[3], addr_3379_6, addr_positional[54079:54076], addr_13519_7);

wire[31:0] addr_13520_7;

Selector_2 s13520_7(wires_3380_6[0], addr_3380_6, addr_positional[54083:54080], addr_13520_7);

wire[31:0] addr_13521_7;

Selector_2 s13521_7(wires_3380_6[1], addr_3380_6, addr_positional[54087:54084], addr_13521_7);

wire[31:0] addr_13522_7;

Selector_2 s13522_7(wires_3380_6[2], addr_3380_6, addr_positional[54091:54088], addr_13522_7);

wire[31:0] addr_13523_7;

Selector_2 s13523_7(wires_3380_6[3], addr_3380_6, addr_positional[54095:54092], addr_13523_7);

wire[31:0] addr_13524_7;

Selector_2 s13524_7(wires_3381_6[0], addr_3381_6, addr_positional[54099:54096], addr_13524_7);

wire[31:0] addr_13525_7;

Selector_2 s13525_7(wires_3381_6[1], addr_3381_6, addr_positional[54103:54100], addr_13525_7);

wire[31:0] addr_13526_7;

Selector_2 s13526_7(wires_3381_6[2], addr_3381_6, addr_positional[54107:54104], addr_13526_7);

wire[31:0] addr_13527_7;

Selector_2 s13527_7(wires_3381_6[3], addr_3381_6, addr_positional[54111:54108], addr_13527_7);

wire[31:0] addr_13528_7;

Selector_2 s13528_7(wires_3382_6[0], addr_3382_6, addr_positional[54115:54112], addr_13528_7);

wire[31:0] addr_13529_7;

Selector_2 s13529_7(wires_3382_6[1], addr_3382_6, addr_positional[54119:54116], addr_13529_7);

wire[31:0] addr_13530_7;

Selector_2 s13530_7(wires_3382_6[2], addr_3382_6, addr_positional[54123:54120], addr_13530_7);

wire[31:0] addr_13531_7;

Selector_2 s13531_7(wires_3382_6[3], addr_3382_6, addr_positional[54127:54124], addr_13531_7);

wire[31:0] addr_13532_7;

Selector_2 s13532_7(wires_3383_6[0], addr_3383_6, addr_positional[54131:54128], addr_13532_7);

wire[31:0] addr_13533_7;

Selector_2 s13533_7(wires_3383_6[1], addr_3383_6, addr_positional[54135:54132], addr_13533_7);

wire[31:0] addr_13534_7;

Selector_2 s13534_7(wires_3383_6[2], addr_3383_6, addr_positional[54139:54136], addr_13534_7);

wire[31:0] addr_13535_7;

Selector_2 s13535_7(wires_3383_6[3], addr_3383_6, addr_positional[54143:54140], addr_13535_7);

wire[31:0] addr_13536_7;

Selector_2 s13536_7(wires_3384_6[0], addr_3384_6, addr_positional[54147:54144], addr_13536_7);

wire[31:0] addr_13537_7;

Selector_2 s13537_7(wires_3384_6[1], addr_3384_6, addr_positional[54151:54148], addr_13537_7);

wire[31:0] addr_13538_7;

Selector_2 s13538_7(wires_3384_6[2], addr_3384_6, addr_positional[54155:54152], addr_13538_7);

wire[31:0] addr_13539_7;

Selector_2 s13539_7(wires_3384_6[3], addr_3384_6, addr_positional[54159:54156], addr_13539_7);

wire[31:0] addr_13540_7;

Selector_2 s13540_7(wires_3385_6[0], addr_3385_6, addr_positional[54163:54160], addr_13540_7);

wire[31:0] addr_13541_7;

Selector_2 s13541_7(wires_3385_6[1], addr_3385_6, addr_positional[54167:54164], addr_13541_7);

wire[31:0] addr_13542_7;

Selector_2 s13542_7(wires_3385_6[2], addr_3385_6, addr_positional[54171:54168], addr_13542_7);

wire[31:0] addr_13543_7;

Selector_2 s13543_7(wires_3385_6[3], addr_3385_6, addr_positional[54175:54172], addr_13543_7);

wire[31:0] addr_13544_7;

Selector_2 s13544_7(wires_3386_6[0], addr_3386_6, addr_positional[54179:54176], addr_13544_7);

wire[31:0] addr_13545_7;

Selector_2 s13545_7(wires_3386_6[1], addr_3386_6, addr_positional[54183:54180], addr_13545_7);

wire[31:0] addr_13546_7;

Selector_2 s13546_7(wires_3386_6[2], addr_3386_6, addr_positional[54187:54184], addr_13546_7);

wire[31:0] addr_13547_7;

Selector_2 s13547_7(wires_3386_6[3], addr_3386_6, addr_positional[54191:54188], addr_13547_7);

wire[31:0] addr_13548_7;

Selector_2 s13548_7(wires_3387_6[0], addr_3387_6, addr_positional[54195:54192], addr_13548_7);

wire[31:0] addr_13549_7;

Selector_2 s13549_7(wires_3387_6[1], addr_3387_6, addr_positional[54199:54196], addr_13549_7);

wire[31:0] addr_13550_7;

Selector_2 s13550_7(wires_3387_6[2], addr_3387_6, addr_positional[54203:54200], addr_13550_7);

wire[31:0] addr_13551_7;

Selector_2 s13551_7(wires_3387_6[3], addr_3387_6, addr_positional[54207:54204], addr_13551_7);

wire[31:0] addr_13552_7;

Selector_2 s13552_7(wires_3388_6[0], addr_3388_6, addr_positional[54211:54208], addr_13552_7);

wire[31:0] addr_13553_7;

Selector_2 s13553_7(wires_3388_6[1], addr_3388_6, addr_positional[54215:54212], addr_13553_7);

wire[31:0] addr_13554_7;

Selector_2 s13554_7(wires_3388_6[2], addr_3388_6, addr_positional[54219:54216], addr_13554_7);

wire[31:0] addr_13555_7;

Selector_2 s13555_7(wires_3388_6[3], addr_3388_6, addr_positional[54223:54220], addr_13555_7);

wire[31:0] addr_13556_7;

Selector_2 s13556_7(wires_3389_6[0], addr_3389_6, addr_positional[54227:54224], addr_13556_7);

wire[31:0] addr_13557_7;

Selector_2 s13557_7(wires_3389_6[1], addr_3389_6, addr_positional[54231:54228], addr_13557_7);

wire[31:0] addr_13558_7;

Selector_2 s13558_7(wires_3389_6[2], addr_3389_6, addr_positional[54235:54232], addr_13558_7);

wire[31:0] addr_13559_7;

Selector_2 s13559_7(wires_3389_6[3], addr_3389_6, addr_positional[54239:54236], addr_13559_7);

wire[31:0] addr_13560_7;

Selector_2 s13560_7(wires_3390_6[0], addr_3390_6, addr_positional[54243:54240], addr_13560_7);

wire[31:0] addr_13561_7;

Selector_2 s13561_7(wires_3390_6[1], addr_3390_6, addr_positional[54247:54244], addr_13561_7);

wire[31:0] addr_13562_7;

Selector_2 s13562_7(wires_3390_6[2], addr_3390_6, addr_positional[54251:54248], addr_13562_7);

wire[31:0] addr_13563_7;

Selector_2 s13563_7(wires_3390_6[3], addr_3390_6, addr_positional[54255:54252], addr_13563_7);

wire[31:0] addr_13564_7;

Selector_2 s13564_7(wires_3391_6[0], addr_3391_6, addr_positional[54259:54256], addr_13564_7);

wire[31:0] addr_13565_7;

Selector_2 s13565_7(wires_3391_6[1], addr_3391_6, addr_positional[54263:54260], addr_13565_7);

wire[31:0] addr_13566_7;

Selector_2 s13566_7(wires_3391_6[2], addr_3391_6, addr_positional[54267:54264], addr_13566_7);

wire[31:0] addr_13567_7;

Selector_2 s13567_7(wires_3391_6[3], addr_3391_6, addr_positional[54271:54268], addr_13567_7);

wire[31:0] addr_13568_7;

Selector_2 s13568_7(wires_3392_6[0], addr_3392_6, addr_positional[54275:54272], addr_13568_7);

wire[31:0] addr_13569_7;

Selector_2 s13569_7(wires_3392_6[1], addr_3392_6, addr_positional[54279:54276], addr_13569_7);

wire[31:0] addr_13570_7;

Selector_2 s13570_7(wires_3392_6[2], addr_3392_6, addr_positional[54283:54280], addr_13570_7);

wire[31:0] addr_13571_7;

Selector_2 s13571_7(wires_3392_6[3], addr_3392_6, addr_positional[54287:54284], addr_13571_7);

wire[31:0] addr_13572_7;

Selector_2 s13572_7(wires_3393_6[0], addr_3393_6, addr_positional[54291:54288], addr_13572_7);

wire[31:0] addr_13573_7;

Selector_2 s13573_7(wires_3393_6[1], addr_3393_6, addr_positional[54295:54292], addr_13573_7);

wire[31:0] addr_13574_7;

Selector_2 s13574_7(wires_3393_6[2], addr_3393_6, addr_positional[54299:54296], addr_13574_7);

wire[31:0] addr_13575_7;

Selector_2 s13575_7(wires_3393_6[3], addr_3393_6, addr_positional[54303:54300], addr_13575_7);

wire[31:0] addr_13576_7;

Selector_2 s13576_7(wires_3394_6[0], addr_3394_6, addr_positional[54307:54304], addr_13576_7);

wire[31:0] addr_13577_7;

Selector_2 s13577_7(wires_3394_6[1], addr_3394_6, addr_positional[54311:54308], addr_13577_7);

wire[31:0] addr_13578_7;

Selector_2 s13578_7(wires_3394_6[2], addr_3394_6, addr_positional[54315:54312], addr_13578_7);

wire[31:0] addr_13579_7;

Selector_2 s13579_7(wires_3394_6[3], addr_3394_6, addr_positional[54319:54316], addr_13579_7);

wire[31:0] addr_13580_7;

Selector_2 s13580_7(wires_3395_6[0], addr_3395_6, addr_positional[54323:54320], addr_13580_7);

wire[31:0] addr_13581_7;

Selector_2 s13581_7(wires_3395_6[1], addr_3395_6, addr_positional[54327:54324], addr_13581_7);

wire[31:0] addr_13582_7;

Selector_2 s13582_7(wires_3395_6[2], addr_3395_6, addr_positional[54331:54328], addr_13582_7);

wire[31:0] addr_13583_7;

Selector_2 s13583_7(wires_3395_6[3], addr_3395_6, addr_positional[54335:54332], addr_13583_7);

wire[31:0] addr_13584_7;

Selector_2 s13584_7(wires_3396_6[0], addr_3396_6, addr_positional[54339:54336], addr_13584_7);

wire[31:0] addr_13585_7;

Selector_2 s13585_7(wires_3396_6[1], addr_3396_6, addr_positional[54343:54340], addr_13585_7);

wire[31:0] addr_13586_7;

Selector_2 s13586_7(wires_3396_6[2], addr_3396_6, addr_positional[54347:54344], addr_13586_7);

wire[31:0] addr_13587_7;

Selector_2 s13587_7(wires_3396_6[3], addr_3396_6, addr_positional[54351:54348], addr_13587_7);

wire[31:0] addr_13588_7;

Selector_2 s13588_7(wires_3397_6[0], addr_3397_6, addr_positional[54355:54352], addr_13588_7);

wire[31:0] addr_13589_7;

Selector_2 s13589_7(wires_3397_6[1], addr_3397_6, addr_positional[54359:54356], addr_13589_7);

wire[31:0] addr_13590_7;

Selector_2 s13590_7(wires_3397_6[2], addr_3397_6, addr_positional[54363:54360], addr_13590_7);

wire[31:0] addr_13591_7;

Selector_2 s13591_7(wires_3397_6[3], addr_3397_6, addr_positional[54367:54364], addr_13591_7);

wire[31:0] addr_13592_7;

Selector_2 s13592_7(wires_3398_6[0], addr_3398_6, addr_positional[54371:54368], addr_13592_7);

wire[31:0] addr_13593_7;

Selector_2 s13593_7(wires_3398_6[1], addr_3398_6, addr_positional[54375:54372], addr_13593_7);

wire[31:0] addr_13594_7;

Selector_2 s13594_7(wires_3398_6[2], addr_3398_6, addr_positional[54379:54376], addr_13594_7);

wire[31:0] addr_13595_7;

Selector_2 s13595_7(wires_3398_6[3], addr_3398_6, addr_positional[54383:54380], addr_13595_7);

wire[31:0] addr_13596_7;

Selector_2 s13596_7(wires_3399_6[0], addr_3399_6, addr_positional[54387:54384], addr_13596_7);

wire[31:0] addr_13597_7;

Selector_2 s13597_7(wires_3399_6[1], addr_3399_6, addr_positional[54391:54388], addr_13597_7);

wire[31:0] addr_13598_7;

Selector_2 s13598_7(wires_3399_6[2], addr_3399_6, addr_positional[54395:54392], addr_13598_7);

wire[31:0] addr_13599_7;

Selector_2 s13599_7(wires_3399_6[3], addr_3399_6, addr_positional[54399:54396], addr_13599_7);

wire[31:0] addr_13600_7;

Selector_2 s13600_7(wires_3400_6[0], addr_3400_6, addr_positional[54403:54400], addr_13600_7);

wire[31:0] addr_13601_7;

Selector_2 s13601_7(wires_3400_6[1], addr_3400_6, addr_positional[54407:54404], addr_13601_7);

wire[31:0] addr_13602_7;

Selector_2 s13602_7(wires_3400_6[2], addr_3400_6, addr_positional[54411:54408], addr_13602_7);

wire[31:0] addr_13603_7;

Selector_2 s13603_7(wires_3400_6[3], addr_3400_6, addr_positional[54415:54412], addr_13603_7);

wire[31:0] addr_13604_7;

Selector_2 s13604_7(wires_3401_6[0], addr_3401_6, addr_positional[54419:54416], addr_13604_7);

wire[31:0] addr_13605_7;

Selector_2 s13605_7(wires_3401_6[1], addr_3401_6, addr_positional[54423:54420], addr_13605_7);

wire[31:0] addr_13606_7;

Selector_2 s13606_7(wires_3401_6[2], addr_3401_6, addr_positional[54427:54424], addr_13606_7);

wire[31:0] addr_13607_7;

Selector_2 s13607_7(wires_3401_6[3], addr_3401_6, addr_positional[54431:54428], addr_13607_7);

wire[31:0] addr_13608_7;

Selector_2 s13608_7(wires_3402_6[0], addr_3402_6, addr_positional[54435:54432], addr_13608_7);

wire[31:0] addr_13609_7;

Selector_2 s13609_7(wires_3402_6[1], addr_3402_6, addr_positional[54439:54436], addr_13609_7);

wire[31:0] addr_13610_7;

Selector_2 s13610_7(wires_3402_6[2], addr_3402_6, addr_positional[54443:54440], addr_13610_7);

wire[31:0] addr_13611_7;

Selector_2 s13611_7(wires_3402_6[3], addr_3402_6, addr_positional[54447:54444], addr_13611_7);

wire[31:0] addr_13612_7;

Selector_2 s13612_7(wires_3403_6[0], addr_3403_6, addr_positional[54451:54448], addr_13612_7);

wire[31:0] addr_13613_7;

Selector_2 s13613_7(wires_3403_6[1], addr_3403_6, addr_positional[54455:54452], addr_13613_7);

wire[31:0] addr_13614_7;

Selector_2 s13614_7(wires_3403_6[2], addr_3403_6, addr_positional[54459:54456], addr_13614_7);

wire[31:0] addr_13615_7;

Selector_2 s13615_7(wires_3403_6[3], addr_3403_6, addr_positional[54463:54460], addr_13615_7);

wire[31:0] addr_13616_7;

Selector_2 s13616_7(wires_3404_6[0], addr_3404_6, addr_positional[54467:54464], addr_13616_7);

wire[31:0] addr_13617_7;

Selector_2 s13617_7(wires_3404_6[1], addr_3404_6, addr_positional[54471:54468], addr_13617_7);

wire[31:0] addr_13618_7;

Selector_2 s13618_7(wires_3404_6[2], addr_3404_6, addr_positional[54475:54472], addr_13618_7);

wire[31:0] addr_13619_7;

Selector_2 s13619_7(wires_3404_6[3], addr_3404_6, addr_positional[54479:54476], addr_13619_7);

wire[31:0] addr_13620_7;

Selector_2 s13620_7(wires_3405_6[0], addr_3405_6, addr_positional[54483:54480], addr_13620_7);

wire[31:0] addr_13621_7;

Selector_2 s13621_7(wires_3405_6[1], addr_3405_6, addr_positional[54487:54484], addr_13621_7);

wire[31:0] addr_13622_7;

Selector_2 s13622_7(wires_3405_6[2], addr_3405_6, addr_positional[54491:54488], addr_13622_7);

wire[31:0] addr_13623_7;

Selector_2 s13623_7(wires_3405_6[3], addr_3405_6, addr_positional[54495:54492], addr_13623_7);

wire[31:0] addr_13624_7;

Selector_2 s13624_7(wires_3406_6[0], addr_3406_6, addr_positional[54499:54496], addr_13624_7);

wire[31:0] addr_13625_7;

Selector_2 s13625_7(wires_3406_6[1], addr_3406_6, addr_positional[54503:54500], addr_13625_7);

wire[31:0] addr_13626_7;

Selector_2 s13626_7(wires_3406_6[2], addr_3406_6, addr_positional[54507:54504], addr_13626_7);

wire[31:0] addr_13627_7;

Selector_2 s13627_7(wires_3406_6[3], addr_3406_6, addr_positional[54511:54508], addr_13627_7);

wire[31:0] addr_13628_7;

Selector_2 s13628_7(wires_3407_6[0], addr_3407_6, addr_positional[54515:54512], addr_13628_7);

wire[31:0] addr_13629_7;

Selector_2 s13629_7(wires_3407_6[1], addr_3407_6, addr_positional[54519:54516], addr_13629_7);

wire[31:0] addr_13630_7;

Selector_2 s13630_7(wires_3407_6[2], addr_3407_6, addr_positional[54523:54520], addr_13630_7);

wire[31:0] addr_13631_7;

Selector_2 s13631_7(wires_3407_6[3], addr_3407_6, addr_positional[54527:54524], addr_13631_7);

wire[31:0] addr_13632_7;

Selector_2 s13632_7(wires_3408_6[0], addr_3408_6, addr_positional[54531:54528], addr_13632_7);

wire[31:0] addr_13633_7;

Selector_2 s13633_7(wires_3408_6[1], addr_3408_6, addr_positional[54535:54532], addr_13633_7);

wire[31:0] addr_13634_7;

Selector_2 s13634_7(wires_3408_6[2], addr_3408_6, addr_positional[54539:54536], addr_13634_7);

wire[31:0] addr_13635_7;

Selector_2 s13635_7(wires_3408_6[3], addr_3408_6, addr_positional[54543:54540], addr_13635_7);

wire[31:0] addr_13636_7;

Selector_2 s13636_7(wires_3409_6[0], addr_3409_6, addr_positional[54547:54544], addr_13636_7);

wire[31:0] addr_13637_7;

Selector_2 s13637_7(wires_3409_6[1], addr_3409_6, addr_positional[54551:54548], addr_13637_7);

wire[31:0] addr_13638_7;

Selector_2 s13638_7(wires_3409_6[2], addr_3409_6, addr_positional[54555:54552], addr_13638_7);

wire[31:0] addr_13639_7;

Selector_2 s13639_7(wires_3409_6[3], addr_3409_6, addr_positional[54559:54556], addr_13639_7);

wire[31:0] addr_13640_7;

Selector_2 s13640_7(wires_3410_6[0], addr_3410_6, addr_positional[54563:54560], addr_13640_7);

wire[31:0] addr_13641_7;

Selector_2 s13641_7(wires_3410_6[1], addr_3410_6, addr_positional[54567:54564], addr_13641_7);

wire[31:0] addr_13642_7;

Selector_2 s13642_7(wires_3410_6[2], addr_3410_6, addr_positional[54571:54568], addr_13642_7);

wire[31:0] addr_13643_7;

Selector_2 s13643_7(wires_3410_6[3], addr_3410_6, addr_positional[54575:54572], addr_13643_7);

wire[31:0] addr_13644_7;

Selector_2 s13644_7(wires_3411_6[0], addr_3411_6, addr_positional[54579:54576], addr_13644_7);

wire[31:0] addr_13645_7;

Selector_2 s13645_7(wires_3411_6[1], addr_3411_6, addr_positional[54583:54580], addr_13645_7);

wire[31:0] addr_13646_7;

Selector_2 s13646_7(wires_3411_6[2], addr_3411_6, addr_positional[54587:54584], addr_13646_7);

wire[31:0] addr_13647_7;

Selector_2 s13647_7(wires_3411_6[3], addr_3411_6, addr_positional[54591:54588], addr_13647_7);

wire[31:0] addr_13648_7;

Selector_2 s13648_7(wires_3412_6[0], addr_3412_6, addr_positional[54595:54592], addr_13648_7);

wire[31:0] addr_13649_7;

Selector_2 s13649_7(wires_3412_6[1], addr_3412_6, addr_positional[54599:54596], addr_13649_7);

wire[31:0] addr_13650_7;

Selector_2 s13650_7(wires_3412_6[2], addr_3412_6, addr_positional[54603:54600], addr_13650_7);

wire[31:0] addr_13651_7;

Selector_2 s13651_7(wires_3412_6[3], addr_3412_6, addr_positional[54607:54604], addr_13651_7);

wire[31:0] addr_13652_7;

Selector_2 s13652_7(wires_3413_6[0], addr_3413_6, addr_positional[54611:54608], addr_13652_7);

wire[31:0] addr_13653_7;

Selector_2 s13653_7(wires_3413_6[1], addr_3413_6, addr_positional[54615:54612], addr_13653_7);

wire[31:0] addr_13654_7;

Selector_2 s13654_7(wires_3413_6[2], addr_3413_6, addr_positional[54619:54616], addr_13654_7);

wire[31:0] addr_13655_7;

Selector_2 s13655_7(wires_3413_6[3], addr_3413_6, addr_positional[54623:54620], addr_13655_7);

wire[31:0] addr_13656_7;

Selector_2 s13656_7(wires_3414_6[0], addr_3414_6, addr_positional[54627:54624], addr_13656_7);

wire[31:0] addr_13657_7;

Selector_2 s13657_7(wires_3414_6[1], addr_3414_6, addr_positional[54631:54628], addr_13657_7);

wire[31:0] addr_13658_7;

Selector_2 s13658_7(wires_3414_6[2], addr_3414_6, addr_positional[54635:54632], addr_13658_7);

wire[31:0] addr_13659_7;

Selector_2 s13659_7(wires_3414_6[3], addr_3414_6, addr_positional[54639:54636], addr_13659_7);

wire[31:0] addr_13660_7;

Selector_2 s13660_7(wires_3415_6[0], addr_3415_6, addr_positional[54643:54640], addr_13660_7);

wire[31:0] addr_13661_7;

Selector_2 s13661_7(wires_3415_6[1], addr_3415_6, addr_positional[54647:54644], addr_13661_7);

wire[31:0] addr_13662_7;

Selector_2 s13662_7(wires_3415_6[2], addr_3415_6, addr_positional[54651:54648], addr_13662_7);

wire[31:0] addr_13663_7;

Selector_2 s13663_7(wires_3415_6[3], addr_3415_6, addr_positional[54655:54652], addr_13663_7);

wire[31:0] addr_13664_7;

Selector_2 s13664_7(wires_3416_6[0], addr_3416_6, addr_positional[54659:54656], addr_13664_7);

wire[31:0] addr_13665_7;

Selector_2 s13665_7(wires_3416_6[1], addr_3416_6, addr_positional[54663:54660], addr_13665_7);

wire[31:0] addr_13666_7;

Selector_2 s13666_7(wires_3416_6[2], addr_3416_6, addr_positional[54667:54664], addr_13666_7);

wire[31:0] addr_13667_7;

Selector_2 s13667_7(wires_3416_6[3], addr_3416_6, addr_positional[54671:54668], addr_13667_7);

wire[31:0] addr_13668_7;

Selector_2 s13668_7(wires_3417_6[0], addr_3417_6, addr_positional[54675:54672], addr_13668_7);

wire[31:0] addr_13669_7;

Selector_2 s13669_7(wires_3417_6[1], addr_3417_6, addr_positional[54679:54676], addr_13669_7);

wire[31:0] addr_13670_7;

Selector_2 s13670_7(wires_3417_6[2], addr_3417_6, addr_positional[54683:54680], addr_13670_7);

wire[31:0] addr_13671_7;

Selector_2 s13671_7(wires_3417_6[3], addr_3417_6, addr_positional[54687:54684], addr_13671_7);

wire[31:0] addr_13672_7;

Selector_2 s13672_7(wires_3418_6[0], addr_3418_6, addr_positional[54691:54688], addr_13672_7);

wire[31:0] addr_13673_7;

Selector_2 s13673_7(wires_3418_6[1], addr_3418_6, addr_positional[54695:54692], addr_13673_7);

wire[31:0] addr_13674_7;

Selector_2 s13674_7(wires_3418_6[2], addr_3418_6, addr_positional[54699:54696], addr_13674_7);

wire[31:0] addr_13675_7;

Selector_2 s13675_7(wires_3418_6[3], addr_3418_6, addr_positional[54703:54700], addr_13675_7);

wire[31:0] addr_13676_7;

Selector_2 s13676_7(wires_3419_6[0], addr_3419_6, addr_positional[54707:54704], addr_13676_7);

wire[31:0] addr_13677_7;

Selector_2 s13677_7(wires_3419_6[1], addr_3419_6, addr_positional[54711:54708], addr_13677_7);

wire[31:0] addr_13678_7;

Selector_2 s13678_7(wires_3419_6[2], addr_3419_6, addr_positional[54715:54712], addr_13678_7);

wire[31:0] addr_13679_7;

Selector_2 s13679_7(wires_3419_6[3], addr_3419_6, addr_positional[54719:54716], addr_13679_7);

wire[31:0] addr_13680_7;

Selector_2 s13680_7(wires_3420_6[0], addr_3420_6, addr_positional[54723:54720], addr_13680_7);

wire[31:0] addr_13681_7;

Selector_2 s13681_7(wires_3420_6[1], addr_3420_6, addr_positional[54727:54724], addr_13681_7);

wire[31:0] addr_13682_7;

Selector_2 s13682_7(wires_3420_6[2], addr_3420_6, addr_positional[54731:54728], addr_13682_7);

wire[31:0] addr_13683_7;

Selector_2 s13683_7(wires_3420_6[3], addr_3420_6, addr_positional[54735:54732], addr_13683_7);

wire[31:0] addr_13684_7;

Selector_2 s13684_7(wires_3421_6[0], addr_3421_6, addr_positional[54739:54736], addr_13684_7);

wire[31:0] addr_13685_7;

Selector_2 s13685_7(wires_3421_6[1], addr_3421_6, addr_positional[54743:54740], addr_13685_7);

wire[31:0] addr_13686_7;

Selector_2 s13686_7(wires_3421_6[2], addr_3421_6, addr_positional[54747:54744], addr_13686_7);

wire[31:0] addr_13687_7;

Selector_2 s13687_7(wires_3421_6[3], addr_3421_6, addr_positional[54751:54748], addr_13687_7);

wire[31:0] addr_13688_7;

Selector_2 s13688_7(wires_3422_6[0], addr_3422_6, addr_positional[54755:54752], addr_13688_7);

wire[31:0] addr_13689_7;

Selector_2 s13689_7(wires_3422_6[1], addr_3422_6, addr_positional[54759:54756], addr_13689_7);

wire[31:0] addr_13690_7;

Selector_2 s13690_7(wires_3422_6[2], addr_3422_6, addr_positional[54763:54760], addr_13690_7);

wire[31:0] addr_13691_7;

Selector_2 s13691_7(wires_3422_6[3], addr_3422_6, addr_positional[54767:54764], addr_13691_7);

wire[31:0] addr_13692_7;

Selector_2 s13692_7(wires_3423_6[0], addr_3423_6, addr_positional[54771:54768], addr_13692_7);

wire[31:0] addr_13693_7;

Selector_2 s13693_7(wires_3423_6[1], addr_3423_6, addr_positional[54775:54772], addr_13693_7);

wire[31:0] addr_13694_7;

Selector_2 s13694_7(wires_3423_6[2], addr_3423_6, addr_positional[54779:54776], addr_13694_7);

wire[31:0] addr_13695_7;

Selector_2 s13695_7(wires_3423_6[3], addr_3423_6, addr_positional[54783:54780], addr_13695_7);

wire[31:0] addr_13696_7;

Selector_2 s13696_7(wires_3424_6[0], addr_3424_6, addr_positional[54787:54784], addr_13696_7);

wire[31:0] addr_13697_7;

Selector_2 s13697_7(wires_3424_6[1], addr_3424_6, addr_positional[54791:54788], addr_13697_7);

wire[31:0] addr_13698_7;

Selector_2 s13698_7(wires_3424_6[2], addr_3424_6, addr_positional[54795:54792], addr_13698_7);

wire[31:0] addr_13699_7;

Selector_2 s13699_7(wires_3424_6[3], addr_3424_6, addr_positional[54799:54796], addr_13699_7);

wire[31:0] addr_13700_7;

Selector_2 s13700_7(wires_3425_6[0], addr_3425_6, addr_positional[54803:54800], addr_13700_7);

wire[31:0] addr_13701_7;

Selector_2 s13701_7(wires_3425_6[1], addr_3425_6, addr_positional[54807:54804], addr_13701_7);

wire[31:0] addr_13702_7;

Selector_2 s13702_7(wires_3425_6[2], addr_3425_6, addr_positional[54811:54808], addr_13702_7);

wire[31:0] addr_13703_7;

Selector_2 s13703_7(wires_3425_6[3], addr_3425_6, addr_positional[54815:54812], addr_13703_7);

wire[31:0] addr_13704_7;

Selector_2 s13704_7(wires_3426_6[0], addr_3426_6, addr_positional[54819:54816], addr_13704_7);

wire[31:0] addr_13705_7;

Selector_2 s13705_7(wires_3426_6[1], addr_3426_6, addr_positional[54823:54820], addr_13705_7);

wire[31:0] addr_13706_7;

Selector_2 s13706_7(wires_3426_6[2], addr_3426_6, addr_positional[54827:54824], addr_13706_7);

wire[31:0] addr_13707_7;

Selector_2 s13707_7(wires_3426_6[3], addr_3426_6, addr_positional[54831:54828], addr_13707_7);

wire[31:0] addr_13708_7;

Selector_2 s13708_7(wires_3427_6[0], addr_3427_6, addr_positional[54835:54832], addr_13708_7);

wire[31:0] addr_13709_7;

Selector_2 s13709_7(wires_3427_6[1], addr_3427_6, addr_positional[54839:54836], addr_13709_7);

wire[31:0] addr_13710_7;

Selector_2 s13710_7(wires_3427_6[2], addr_3427_6, addr_positional[54843:54840], addr_13710_7);

wire[31:0] addr_13711_7;

Selector_2 s13711_7(wires_3427_6[3], addr_3427_6, addr_positional[54847:54844], addr_13711_7);

wire[31:0] addr_13712_7;

Selector_2 s13712_7(wires_3428_6[0], addr_3428_6, addr_positional[54851:54848], addr_13712_7);

wire[31:0] addr_13713_7;

Selector_2 s13713_7(wires_3428_6[1], addr_3428_6, addr_positional[54855:54852], addr_13713_7);

wire[31:0] addr_13714_7;

Selector_2 s13714_7(wires_3428_6[2], addr_3428_6, addr_positional[54859:54856], addr_13714_7);

wire[31:0] addr_13715_7;

Selector_2 s13715_7(wires_3428_6[3], addr_3428_6, addr_positional[54863:54860], addr_13715_7);

wire[31:0] addr_13716_7;

Selector_2 s13716_7(wires_3429_6[0], addr_3429_6, addr_positional[54867:54864], addr_13716_7);

wire[31:0] addr_13717_7;

Selector_2 s13717_7(wires_3429_6[1], addr_3429_6, addr_positional[54871:54868], addr_13717_7);

wire[31:0] addr_13718_7;

Selector_2 s13718_7(wires_3429_6[2], addr_3429_6, addr_positional[54875:54872], addr_13718_7);

wire[31:0] addr_13719_7;

Selector_2 s13719_7(wires_3429_6[3], addr_3429_6, addr_positional[54879:54876], addr_13719_7);

wire[31:0] addr_13720_7;

Selector_2 s13720_7(wires_3430_6[0], addr_3430_6, addr_positional[54883:54880], addr_13720_7);

wire[31:0] addr_13721_7;

Selector_2 s13721_7(wires_3430_6[1], addr_3430_6, addr_positional[54887:54884], addr_13721_7);

wire[31:0] addr_13722_7;

Selector_2 s13722_7(wires_3430_6[2], addr_3430_6, addr_positional[54891:54888], addr_13722_7);

wire[31:0] addr_13723_7;

Selector_2 s13723_7(wires_3430_6[3], addr_3430_6, addr_positional[54895:54892], addr_13723_7);

wire[31:0] addr_13724_7;

Selector_2 s13724_7(wires_3431_6[0], addr_3431_6, addr_positional[54899:54896], addr_13724_7);

wire[31:0] addr_13725_7;

Selector_2 s13725_7(wires_3431_6[1], addr_3431_6, addr_positional[54903:54900], addr_13725_7);

wire[31:0] addr_13726_7;

Selector_2 s13726_7(wires_3431_6[2], addr_3431_6, addr_positional[54907:54904], addr_13726_7);

wire[31:0] addr_13727_7;

Selector_2 s13727_7(wires_3431_6[3], addr_3431_6, addr_positional[54911:54908], addr_13727_7);

wire[31:0] addr_13728_7;

Selector_2 s13728_7(wires_3432_6[0], addr_3432_6, addr_positional[54915:54912], addr_13728_7);

wire[31:0] addr_13729_7;

Selector_2 s13729_7(wires_3432_6[1], addr_3432_6, addr_positional[54919:54916], addr_13729_7);

wire[31:0] addr_13730_7;

Selector_2 s13730_7(wires_3432_6[2], addr_3432_6, addr_positional[54923:54920], addr_13730_7);

wire[31:0] addr_13731_7;

Selector_2 s13731_7(wires_3432_6[3], addr_3432_6, addr_positional[54927:54924], addr_13731_7);

wire[31:0] addr_13732_7;

Selector_2 s13732_7(wires_3433_6[0], addr_3433_6, addr_positional[54931:54928], addr_13732_7);

wire[31:0] addr_13733_7;

Selector_2 s13733_7(wires_3433_6[1], addr_3433_6, addr_positional[54935:54932], addr_13733_7);

wire[31:0] addr_13734_7;

Selector_2 s13734_7(wires_3433_6[2], addr_3433_6, addr_positional[54939:54936], addr_13734_7);

wire[31:0] addr_13735_7;

Selector_2 s13735_7(wires_3433_6[3], addr_3433_6, addr_positional[54943:54940], addr_13735_7);

wire[31:0] addr_13736_7;

Selector_2 s13736_7(wires_3434_6[0], addr_3434_6, addr_positional[54947:54944], addr_13736_7);

wire[31:0] addr_13737_7;

Selector_2 s13737_7(wires_3434_6[1], addr_3434_6, addr_positional[54951:54948], addr_13737_7);

wire[31:0] addr_13738_7;

Selector_2 s13738_7(wires_3434_6[2], addr_3434_6, addr_positional[54955:54952], addr_13738_7);

wire[31:0] addr_13739_7;

Selector_2 s13739_7(wires_3434_6[3], addr_3434_6, addr_positional[54959:54956], addr_13739_7);

wire[31:0] addr_13740_7;

Selector_2 s13740_7(wires_3435_6[0], addr_3435_6, addr_positional[54963:54960], addr_13740_7);

wire[31:0] addr_13741_7;

Selector_2 s13741_7(wires_3435_6[1], addr_3435_6, addr_positional[54967:54964], addr_13741_7);

wire[31:0] addr_13742_7;

Selector_2 s13742_7(wires_3435_6[2], addr_3435_6, addr_positional[54971:54968], addr_13742_7);

wire[31:0] addr_13743_7;

Selector_2 s13743_7(wires_3435_6[3], addr_3435_6, addr_positional[54975:54972], addr_13743_7);

wire[31:0] addr_13744_7;

Selector_2 s13744_7(wires_3436_6[0], addr_3436_6, addr_positional[54979:54976], addr_13744_7);

wire[31:0] addr_13745_7;

Selector_2 s13745_7(wires_3436_6[1], addr_3436_6, addr_positional[54983:54980], addr_13745_7);

wire[31:0] addr_13746_7;

Selector_2 s13746_7(wires_3436_6[2], addr_3436_6, addr_positional[54987:54984], addr_13746_7);

wire[31:0] addr_13747_7;

Selector_2 s13747_7(wires_3436_6[3], addr_3436_6, addr_positional[54991:54988], addr_13747_7);

wire[31:0] addr_13748_7;

Selector_2 s13748_7(wires_3437_6[0], addr_3437_6, addr_positional[54995:54992], addr_13748_7);

wire[31:0] addr_13749_7;

Selector_2 s13749_7(wires_3437_6[1], addr_3437_6, addr_positional[54999:54996], addr_13749_7);

wire[31:0] addr_13750_7;

Selector_2 s13750_7(wires_3437_6[2], addr_3437_6, addr_positional[55003:55000], addr_13750_7);

wire[31:0] addr_13751_7;

Selector_2 s13751_7(wires_3437_6[3], addr_3437_6, addr_positional[55007:55004], addr_13751_7);

wire[31:0] addr_13752_7;

Selector_2 s13752_7(wires_3438_6[0], addr_3438_6, addr_positional[55011:55008], addr_13752_7);

wire[31:0] addr_13753_7;

Selector_2 s13753_7(wires_3438_6[1], addr_3438_6, addr_positional[55015:55012], addr_13753_7);

wire[31:0] addr_13754_7;

Selector_2 s13754_7(wires_3438_6[2], addr_3438_6, addr_positional[55019:55016], addr_13754_7);

wire[31:0] addr_13755_7;

Selector_2 s13755_7(wires_3438_6[3], addr_3438_6, addr_positional[55023:55020], addr_13755_7);

wire[31:0] addr_13756_7;

Selector_2 s13756_7(wires_3439_6[0], addr_3439_6, addr_positional[55027:55024], addr_13756_7);

wire[31:0] addr_13757_7;

Selector_2 s13757_7(wires_3439_6[1], addr_3439_6, addr_positional[55031:55028], addr_13757_7);

wire[31:0] addr_13758_7;

Selector_2 s13758_7(wires_3439_6[2], addr_3439_6, addr_positional[55035:55032], addr_13758_7);

wire[31:0] addr_13759_7;

Selector_2 s13759_7(wires_3439_6[3], addr_3439_6, addr_positional[55039:55036], addr_13759_7);

wire[31:0] addr_13760_7;

Selector_2 s13760_7(wires_3440_6[0], addr_3440_6, addr_positional[55043:55040], addr_13760_7);

wire[31:0] addr_13761_7;

Selector_2 s13761_7(wires_3440_6[1], addr_3440_6, addr_positional[55047:55044], addr_13761_7);

wire[31:0] addr_13762_7;

Selector_2 s13762_7(wires_3440_6[2], addr_3440_6, addr_positional[55051:55048], addr_13762_7);

wire[31:0] addr_13763_7;

Selector_2 s13763_7(wires_3440_6[3], addr_3440_6, addr_positional[55055:55052], addr_13763_7);

wire[31:0] addr_13764_7;

Selector_2 s13764_7(wires_3441_6[0], addr_3441_6, addr_positional[55059:55056], addr_13764_7);

wire[31:0] addr_13765_7;

Selector_2 s13765_7(wires_3441_6[1], addr_3441_6, addr_positional[55063:55060], addr_13765_7);

wire[31:0] addr_13766_7;

Selector_2 s13766_7(wires_3441_6[2], addr_3441_6, addr_positional[55067:55064], addr_13766_7);

wire[31:0] addr_13767_7;

Selector_2 s13767_7(wires_3441_6[3], addr_3441_6, addr_positional[55071:55068], addr_13767_7);

wire[31:0] addr_13768_7;

Selector_2 s13768_7(wires_3442_6[0], addr_3442_6, addr_positional[55075:55072], addr_13768_7);

wire[31:0] addr_13769_7;

Selector_2 s13769_7(wires_3442_6[1], addr_3442_6, addr_positional[55079:55076], addr_13769_7);

wire[31:0] addr_13770_7;

Selector_2 s13770_7(wires_3442_6[2], addr_3442_6, addr_positional[55083:55080], addr_13770_7);

wire[31:0] addr_13771_7;

Selector_2 s13771_7(wires_3442_6[3], addr_3442_6, addr_positional[55087:55084], addr_13771_7);

wire[31:0] addr_13772_7;

Selector_2 s13772_7(wires_3443_6[0], addr_3443_6, addr_positional[55091:55088], addr_13772_7);

wire[31:0] addr_13773_7;

Selector_2 s13773_7(wires_3443_6[1], addr_3443_6, addr_positional[55095:55092], addr_13773_7);

wire[31:0] addr_13774_7;

Selector_2 s13774_7(wires_3443_6[2], addr_3443_6, addr_positional[55099:55096], addr_13774_7);

wire[31:0] addr_13775_7;

Selector_2 s13775_7(wires_3443_6[3], addr_3443_6, addr_positional[55103:55100], addr_13775_7);

wire[31:0] addr_13776_7;

Selector_2 s13776_7(wires_3444_6[0], addr_3444_6, addr_positional[55107:55104], addr_13776_7);

wire[31:0] addr_13777_7;

Selector_2 s13777_7(wires_3444_6[1], addr_3444_6, addr_positional[55111:55108], addr_13777_7);

wire[31:0] addr_13778_7;

Selector_2 s13778_7(wires_3444_6[2], addr_3444_6, addr_positional[55115:55112], addr_13778_7);

wire[31:0] addr_13779_7;

Selector_2 s13779_7(wires_3444_6[3], addr_3444_6, addr_positional[55119:55116], addr_13779_7);

wire[31:0] addr_13780_7;

Selector_2 s13780_7(wires_3445_6[0], addr_3445_6, addr_positional[55123:55120], addr_13780_7);

wire[31:0] addr_13781_7;

Selector_2 s13781_7(wires_3445_6[1], addr_3445_6, addr_positional[55127:55124], addr_13781_7);

wire[31:0] addr_13782_7;

Selector_2 s13782_7(wires_3445_6[2], addr_3445_6, addr_positional[55131:55128], addr_13782_7);

wire[31:0] addr_13783_7;

Selector_2 s13783_7(wires_3445_6[3], addr_3445_6, addr_positional[55135:55132], addr_13783_7);

wire[31:0] addr_13784_7;

Selector_2 s13784_7(wires_3446_6[0], addr_3446_6, addr_positional[55139:55136], addr_13784_7);

wire[31:0] addr_13785_7;

Selector_2 s13785_7(wires_3446_6[1], addr_3446_6, addr_positional[55143:55140], addr_13785_7);

wire[31:0] addr_13786_7;

Selector_2 s13786_7(wires_3446_6[2], addr_3446_6, addr_positional[55147:55144], addr_13786_7);

wire[31:0] addr_13787_7;

Selector_2 s13787_7(wires_3446_6[3], addr_3446_6, addr_positional[55151:55148], addr_13787_7);

wire[31:0] addr_13788_7;

Selector_2 s13788_7(wires_3447_6[0], addr_3447_6, addr_positional[55155:55152], addr_13788_7);

wire[31:0] addr_13789_7;

Selector_2 s13789_7(wires_3447_6[1], addr_3447_6, addr_positional[55159:55156], addr_13789_7);

wire[31:0] addr_13790_7;

Selector_2 s13790_7(wires_3447_6[2], addr_3447_6, addr_positional[55163:55160], addr_13790_7);

wire[31:0] addr_13791_7;

Selector_2 s13791_7(wires_3447_6[3], addr_3447_6, addr_positional[55167:55164], addr_13791_7);

wire[31:0] addr_13792_7;

Selector_2 s13792_7(wires_3448_6[0], addr_3448_6, addr_positional[55171:55168], addr_13792_7);

wire[31:0] addr_13793_7;

Selector_2 s13793_7(wires_3448_6[1], addr_3448_6, addr_positional[55175:55172], addr_13793_7);

wire[31:0] addr_13794_7;

Selector_2 s13794_7(wires_3448_6[2], addr_3448_6, addr_positional[55179:55176], addr_13794_7);

wire[31:0] addr_13795_7;

Selector_2 s13795_7(wires_3448_6[3], addr_3448_6, addr_positional[55183:55180], addr_13795_7);

wire[31:0] addr_13796_7;

Selector_2 s13796_7(wires_3449_6[0], addr_3449_6, addr_positional[55187:55184], addr_13796_7);

wire[31:0] addr_13797_7;

Selector_2 s13797_7(wires_3449_6[1], addr_3449_6, addr_positional[55191:55188], addr_13797_7);

wire[31:0] addr_13798_7;

Selector_2 s13798_7(wires_3449_6[2], addr_3449_6, addr_positional[55195:55192], addr_13798_7);

wire[31:0] addr_13799_7;

Selector_2 s13799_7(wires_3449_6[3], addr_3449_6, addr_positional[55199:55196], addr_13799_7);

wire[31:0] addr_13800_7;

Selector_2 s13800_7(wires_3450_6[0], addr_3450_6, addr_positional[55203:55200], addr_13800_7);

wire[31:0] addr_13801_7;

Selector_2 s13801_7(wires_3450_6[1], addr_3450_6, addr_positional[55207:55204], addr_13801_7);

wire[31:0] addr_13802_7;

Selector_2 s13802_7(wires_3450_6[2], addr_3450_6, addr_positional[55211:55208], addr_13802_7);

wire[31:0] addr_13803_7;

Selector_2 s13803_7(wires_3450_6[3], addr_3450_6, addr_positional[55215:55212], addr_13803_7);

wire[31:0] addr_13804_7;

Selector_2 s13804_7(wires_3451_6[0], addr_3451_6, addr_positional[55219:55216], addr_13804_7);

wire[31:0] addr_13805_7;

Selector_2 s13805_7(wires_3451_6[1], addr_3451_6, addr_positional[55223:55220], addr_13805_7);

wire[31:0] addr_13806_7;

Selector_2 s13806_7(wires_3451_6[2], addr_3451_6, addr_positional[55227:55224], addr_13806_7);

wire[31:0] addr_13807_7;

Selector_2 s13807_7(wires_3451_6[3], addr_3451_6, addr_positional[55231:55228], addr_13807_7);

wire[31:0] addr_13808_7;

Selector_2 s13808_7(wires_3452_6[0], addr_3452_6, addr_positional[55235:55232], addr_13808_7);

wire[31:0] addr_13809_7;

Selector_2 s13809_7(wires_3452_6[1], addr_3452_6, addr_positional[55239:55236], addr_13809_7);

wire[31:0] addr_13810_7;

Selector_2 s13810_7(wires_3452_6[2], addr_3452_6, addr_positional[55243:55240], addr_13810_7);

wire[31:0] addr_13811_7;

Selector_2 s13811_7(wires_3452_6[3], addr_3452_6, addr_positional[55247:55244], addr_13811_7);

wire[31:0] addr_13812_7;

Selector_2 s13812_7(wires_3453_6[0], addr_3453_6, addr_positional[55251:55248], addr_13812_7);

wire[31:0] addr_13813_7;

Selector_2 s13813_7(wires_3453_6[1], addr_3453_6, addr_positional[55255:55252], addr_13813_7);

wire[31:0] addr_13814_7;

Selector_2 s13814_7(wires_3453_6[2], addr_3453_6, addr_positional[55259:55256], addr_13814_7);

wire[31:0] addr_13815_7;

Selector_2 s13815_7(wires_3453_6[3], addr_3453_6, addr_positional[55263:55260], addr_13815_7);

wire[31:0] addr_13816_7;

Selector_2 s13816_7(wires_3454_6[0], addr_3454_6, addr_positional[55267:55264], addr_13816_7);

wire[31:0] addr_13817_7;

Selector_2 s13817_7(wires_3454_6[1], addr_3454_6, addr_positional[55271:55268], addr_13817_7);

wire[31:0] addr_13818_7;

Selector_2 s13818_7(wires_3454_6[2], addr_3454_6, addr_positional[55275:55272], addr_13818_7);

wire[31:0] addr_13819_7;

Selector_2 s13819_7(wires_3454_6[3], addr_3454_6, addr_positional[55279:55276], addr_13819_7);

wire[31:0] addr_13820_7;

Selector_2 s13820_7(wires_3455_6[0], addr_3455_6, addr_positional[55283:55280], addr_13820_7);

wire[31:0] addr_13821_7;

Selector_2 s13821_7(wires_3455_6[1], addr_3455_6, addr_positional[55287:55284], addr_13821_7);

wire[31:0] addr_13822_7;

Selector_2 s13822_7(wires_3455_6[2], addr_3455_6, addr_positional[55291:55288], addr_13822_7);

wire[31:0] addr_13823_7;

Selector_2 s13823_7(wires_3455_6[3], addr_3455_6, addr_positional[55295:55292], addr_13823_7);

wire[31:0] addr_13824_7;

Selector_2 s13824_7(wires_3456_6[0], addr_3456_6, addr_positional[55299:55296], addr_13824_7);

wire[31:0] addr_13825_7;

Selector_2 s13825_7(wires_3456_6[1], addr_3456_6, addr_positional[55303:55300], addr_13825_7);

wire[31:0] addr_13826_7;

Selector_2 s13826_7(wires_3456_6[2], addr_3456_6, addr_positional[55307:55304], addr_13826_7);

wire[31:0] addr_13827_7;

Selector_2 s13827_7(wires_3456_6[3], addr_3456_6, addr_positional[55311:55308], addr_13827_7);

wire[31:0] addr_13828_7;

Selector_2 s13828_7(wires_3457_6[0], addr_3457_6, addr_positional[55315:55312], addr_13828_7);

wire[31:0] addr_13829_7;

Selector_2 s13829_7(wires_3457_6[1], addr_3457_6, addr_positional[55319:55316], addr_13829_7);

wire[31:0] addr_13830_7;

Selector_2 s13830_7(wires_3457_6[2], addr_3457_6, addr_positional[55323:55320], addr_13830_7);

wire[31:0] addr_13831_7;

Selector_2 s13831_7(wires_3457_6[3], addr_3457_6, addr_positional[55327:55324], addr_13831_7);

wire[31:0] addr_13832_7;

Selector_2 s13832_7(wires_3458_6[0], addr_3458_6, addr_positional[55331:55328], addr_13832_7);

wire[31:0] addr_13833_7;

Selector_2 s13833_7(wires_3458_6[1], addr_3458_6, addr_positional[55335:55332], addr_13833_7);

wire[31:0] addr_13834_7;

Selector_2 s13834_7(wires_3458_6[2], addr_3458_6, addr_positional[55339:55336], addr_13834_7);

wire[31:0] addr_13835_7;

Selector_2 s13835_7(wires_3458_6[3], addr_3458_6, addr_positional[55343:55340], addr_13835_7);

wire[31:0] addr_13836_7;

Selector_2 s13836_7(wires_3459_6[0], addr_3459_6, addr_positional[55347:55344], addr_13836_7);

wire[31:0] addr_13837_7;

Selector_2 s13837_7(wires_3459_6[1], addr_3459_6, addr_positional[55351:55348], addr_13837_7);

wire[31:0] addr_13838_7;

Selector_2 s13838_7(wires_3459_6[2], addr_3459_6, addr_positional[55355:55352], addr_13838_7);

wire[31:0] addr_13839_7;

Selector_2 s13839_7(wires_3459_6[3], addr_3459_6, addr_positional[55359:55356], addr_13839_7);

wire[31:0] addr_13840_7;

Selector_2 s13840_7(wires_3460_6[0], addr_3460_6, addr_positional[55363:55360], addr_13840_7);

wire[31:0] addr_13841_7;

Selector_2 s13841_7(wires_3460_6[1], addr_3460_6, addr_positional[55367:55364], addr_13841_7);

wire[31:0] addr_13842_7;

Selector_2 s13842_7(wires_3460_6[2], addr_3460_6, addr_positional[55371:55368], addr_13842_7);

wire[31:0] addr_13843_7;

Selector_2 s13843_7(wires_3460_6[3], addr_3460_6, addr_positional[55375:55372], addr_13843_7);

wire[31:0] addr_13844_7;

Selector_2 s13844_7(wires_3461_6[0], addr_3461_6, addr_positional[55379:55376], addr_13844_7);

wire[31:0] addr_13845_7;

Selector_2 s13845_7(wires_3461_6[1], addr_3461_6, addr_positional[55383:55380], addr_13845_7);

wire[31:0] addr_13846_7;

Selector_2 s13846_7(wires_3461_6[2], addr_3461_6, addr_positional[55387:55384], addr_13846_7);

wire[31:0] addr_13847_7;

Selector_2 s13847_7(wires_3461_6[3], addr_3461_6, addr_positional[55391:55388], addr_13847_7);

wire[31:0] addr_13848_7;

Selector_2 s13848_7(wires_3462_6[0], addr_3462_6, addr_positional[55395:55392], addr_13848_7);

wire[31:0] addr_13849_7;

Selector_2 s13849_7(wires_3462_6[1], addr_3462_6, addr_positional[55399:55396], addr_13849_7);

wire[31:0] addr_13850_7;

Selector_2 s13850_7(wires_3462_6[2], addr_3462_6, addr_positional[55403:55400], addr_13850_7);

wire[31:0] addr_13851_7;

Selector_2 s13851_7(wires_3462_6[3], addr_3462_6, addr_positional[55407:55404], addr_13851_7);

wire[31:0] addr_13852_7;

Selector_2 s13852_7(wires_3463_6[0], addr_3463_6, addr_positional[55411:55408], addr_13852_7);

wire[31:0] addr_13853_7;

Selector_2 s13853_7(wires_3463_6[1], addr_3463_6, addr_positional[55415:55412], addr_13853_7);

wire[31:0] addr_13854_7;

Selector_2 s13854_7(wires_3463_6[2], addr_3463_6, addr_positional[55419:55416], addr_13854_7);

wire[31:0] addr_13855_7;

Selector_2 s13855_7(wires_3463_6[3], addr_3463_6, addr_positional[55423:55420], addr_13855_7);

wire[31:0] addr_13856_7;

Selector_2 s13856_7(wires_3464_6[0], addr_3464_6, addr_positional[55427:55424], addr_13856_7);

wire[31:0] addr_13857_7;

Selector_2 s13857_7(wires_3464_6[1], addr_3464_6, addr_positional[55431:55428], addr_13857_7);

wire[31:0] addr_13858_7;

Selector_2 s13858_7(wires_3464_6[2], addr_3464_6, addr_positional[55435:55432], addr_13858_7);

wire[31:0] addr_13859_7;

Selector_2 s13859_7(wires_3464_6[3], addr_3464_6, addr_positional[55439:55436], addr_13859_7);

wire[31:0] addr_13860_7;

Selector_2 s13860_7(wires_3465_6[0], addr_3465_6, addr_positional[55443:55440], addr_13860_7);

wire[31:0] addr_13861_7;

Selector_2 s13861_7(wires_3465_6[1], addr_3465_6, addr_positional[55447:55444], addr_13861_7);

wire[31:0] addr_13862_7;

Selector_2 s13862_7(wires_3465_6[2], addr_3465_6, addr_positional[55451:55448], addr_13862_7);

wire[31:0] addr_13863_7;

Selector_2 s13863_7(wires_3465_6[3], addr_3465_6, addr_positional[55455:55452], addr_13863_7);

wire[31:0] addr_13864_7;

Selector_2 s13864_7(wires_3466_6[0], addr_3466_6, addr_positional[55459:55456], addr_13864_7);

wire[31:0] addr_13865_7;

Selector_2 s13865_7(wires_3466_6[1], addr_3466_6, addr_positional[55463:55460], addr_13865_7);

wire[31:0] addr_13866_7;

Selector_2 s13866_7(wires_3466_6[2], addr_3466_6, addr_positional[55467:55464], addr_13866_7);

wire[31:0] addr_13867_7;

Selector_2 s13867_7(wires_3466_6[3], addr_3466_6, addr_positional[55471:55468], addr_13867_7);

wire[31:0] addr_13868_7;

Selector_2 s13868_7(wires_3467_6[0], addr_3467_6, addr_positional[55475:55472], addr_13868_7);

wire[31:0] addr_13869_7;

Selector_2 s13869_7(wires_3467_6[1], addr_3467_6, addr_positional[55479:55476], addr_13869_7);

wire[31:0] addr_13870_7;

Selector_2 s13870_7(wires_3467_6[2], addr_3467_6, addr_positional[55483:55480], addr_13870_7);

wire[31:0] addr_13871_7;

Selector_2 s13871_7(wires_3467_6[3], addr_3467_6, addr_positional[55487:55484], addr_13871_7);

wire[31:0] addr_13872_7;

Selector_2 s13872_7(wires_3468_6[0], addr_3468_6, addr_positional[55491:55488], addr_13872_7);

wire[31:0] addr_13873_7;

Selector_2 s13873_7(wires_3468_6[1], addr_3468_6, addr_positional[55495:55492], addr_13873_7);

wire[31:0] addr_13874_7;

Selector_2 s13874_7(wires_3468_6[2], addr_3468_6, addr_positional[55499:55496], addr_13874_7);

wire[31:0] addr_13875_7;

Selector_2 s13875_7(wires_3468_6[3], addr_3468_6, addr_positional[55503:55500], addr_13875_7);

wire[31:0] addr_13876_7;

Selector_2 s13876_7(wires_3469_6[0], addr_3469_6, addr_positional[55507:55504], addr_13876_7);

wire[31:0] addr_13877_7;

Selector_2 s13877_7(wires_3469_6[1], addr_3469_6, addr_positional[55511:55508], addr_13877_7);

wire[31:0] addr_13878_7;

Selector_2 s13878_7(wires_3469_6[2], addr_3469_6, addr_positional[55515:55512], addr_13878_7);

wire[31:0] addr_13879_7;

Selector_2 s13879_7(wires_3469_6[3], addr_3469_6, addr_positional[55519:55516], addr_13879_7);

wire[31:0] addr_13880_7;

Selector_2 s13880_7(wires_3470_6[0], addr_3470_6, addr_positional[55523:55520], addr_13880_7);

wire[31:0] addr_13881_7;

Selector_2 s13881_7(wires_3470_6[1], addr_3470_6, addr_positional[55527:55524], addr_13881_7);

wire[31:0] addr_13882_7;

Selector_2 s13882_7(wires_3470_6[2], addr_3470_6, addr_positional[55531:55528], addr_13882_7);

wire[31:0] addr_13883_7;

Selector_2 s13883_7(wires_3470_6[3], addr_3470_6, addr_positional[55535:55532], addr_13883_7);

wire[31:0] addr_13884_7;

Selector_2 s13884_7(wires_3471_6[0], addr_3471_6, addr_positional[55539:55536], addr_13884_7);

wire[31:0] addr_13885_7;

Selector_2 s13885_7(wires_3471_6[1], addr_3471_6, addr_positional[55543:55540], addr_13885_7);

wire[31:0] addr_13886_7;

Selector_2 s13886_7(wires_3471_6[2], addr_3471_6, addr_positional[55547:55544], addr_13886_7);

wire[31:0] addr_13887_7;

Selector_2 s13887_7(wires_3471_6[3], addr_3471_6, addr_positional[55551:55548], addr_13887_7);

wire[31:0] addr_13888_7;

Selector_2 s13888_7(wires_3472_6[0], addr_3472_6, addr_positional[55555:55552], addr_13888_7);

wire[31:0] addr_13889_7;

Selector_2 s13889_7(wires_3472_6[1], addr_3472_6, addr_positional[55559:55556], addr_13889_7);

wire[31:0] addr_13890_7;

Selector_2 s13890_7(wires_3472_6[2], addr_3472_6, addr_positional[55563:55560], addr_13890_7);

wire[31:0] addr_13891_7;

Selector_2 s13891_7(wires_3472_6[3], addr_3472_6, addr_positional[55567:55564], addr_13891_7);

wire[31:0] addr_13892_7;

Selector_2 s13892_7(wires_3473_6[0], addr_3473_6, addr_positional[55571:55568], addr_13892_7);

wire[31:0] addr_13893_7;

Selector_2 s13893_7(wires_3473_6[1], addr_3473_6, addr_positional[55575:55572], addr_13893_7);

wire[31:0] addr_13894_7;

Selector_2 s13894_7(wires_3473_6[2], addr_3473_6, addr_positional[55579:55576], addr_13894_7);

wire[31:0] addr_13895_7;

Selector_2 s13895_7(wires_3473_6[3], addr_3473_6, addr_positional[55583:55580], addr_13895_7);

wire[31:0] addr_13896_7;

Selector_2 s13896_7(wires_3474_6[0], addr_3474_6, addr_positional[55587:55584], addr_13896_7);

wire[31:0] addr_13897_7;

Selector_2 s13897_7(wires_3474_6[1], addr_3474_6, addr_positional[55591:55588], addr_13897_7);

wire[31:0] addr_13898_7;

Selector_2 s13898_7(wires_3474_6[2], addr_3474_6, addr_positional[55595:55592], addr_13898_7);

wire[31:0] addr_13899_7;

Selector_2 s13899_7(wires_3474_6[3], addr_3474_6, addr_positional[55599:55596], addr_13899_7);

wire[31:0] addr_13900_7;

Selector_2 s13900_7(wires_3475_6[0], addr_3475_6, addr_positional[55603:55600], addr_13900_7);

wire[31:0] addr_13901_7;

Selector_2 s13901_7(wires_3475_6[1], addr_3475_6, addr_positional[55607:55604], addr_13901_7);

wire[31:0] addr_13902_7;

Selector_2 s13902_7(wires_3475_6[2], addr_3475_6, addr_positional[55611:55608], addr_13902_7);

wire[31:0] addr_13903_7;

Selector_2 s13903_7(wires_3475_6[3], addr_3475_6, addr_positional[55615:55612], addr_13903_7);

wire[31:0] addr_13904_7;

Selector_2 s13904_7(wires_3476_6[0], addr_3476_6, addr_positional[55619:55616], addr_13904_7);

wire[31:0] addr_13905_7;

Selector_2 s13905_7(wires_3476_6[1], addr_3476_6, addr_positional[55623:55620], addr_13905_7);

wire[31:0] addr_13906_7;

Selector_2 s13906_7(wires_3476_6[2], addr_3476_6, addr_positional[55627:55624], addr_13906_7);

wire[31:0] addr_13907_7;

Selector_2 s13907_7(wires_3476_6[3], addr_3476_6, addr_positional[55631:55628], addr_13907_7);

wire[31:0] addr_13908_7;

Selector_2 s13908_7(wires_3477_6[0], addr_3477_6, addr_positional[55635:55632], addr_13908_7);

wire[31:0] addr_13909_7;

Selector_2 s13909_7(wires_3477_6[1], addr_3477_6, addr_positional[55639:55636], addr_13909_7);

wire[31:0] addr_13910_7;

Selector_2 s13910_7(wires_3477_6[2], addr_3477_6, addr_positional[55643:55640], addr_13910_7);

wire[31:0] addr_13911_7;

Selector_2 s13911_7(wires_3477_6[3], addr_3477_6, addr_positional[55647:55644], addr_13911_7);

wire[31:0] addr_13912_7;

Selector_2 s13912_7(wires_3478_6[0], addr_3478_6, addr_positional[55651:55648], addr_13912_7);

wire[31:0] addr_13913_7;

Selector_2 s13913_7(wires_3478_6[1], addr_3478_6, addr_positional[55655:55652], addr_13913_7);

wire[31:0] addr_13914_7;

Selector_2 s13914_7(wires_3478_6[2], addr_3478_6, addr_positional[55659:55656], addr_13914_7);

wire[31:0] addr_13915_7;

Selector_2 s13915_7(wires_3478_6[3], addr_3478_6, addr_positional[55663:55660], addr_13915_7);

wire[31:0] addr_13916_7;

Selector_2 s13916_7(wires_3479_6[0], addr_3479_6, addr_positional[55667:55664], addr_13916_7);

wire[31:0] addr_13917_7;

Selector_2 s13917_7(wires_3479_6[1], addr_3479_6, addr_positional[55671:55668], addr_13917_7);

wire[31:0] addr_13918_7;

Selector_2 s13918_7(wires_3479_6[2], addr_3479_6, addr_positional[55675:55672], addr_13918_7);

wire[31:0] addr_13919_7;

Selector_2 s13919_7(wires_3479_6[3], addr_3479_6, addr_positional[55679:55676], addr_13919_7);

wire[31:0] addr_13920_7;

Selector_2 s13920_7(wires_3480_6[0], addr_3480_6, addr_positional[55683:55680], addr_13920_7);

wire[31:0] addr_13921_7;

Selector_2 s13921_7(wires_3480_6[1], addr_3480_6, addr_positional[55687:55684], addr_13921_7);

wire[31:0] addr_13922_7;

Selector_2 s13922_7(wires_3480_6[2], addr_3480_6, addr_positional[55691:55688], addr_13922_7);

wire[31:0] addr_13923_7;

Selector_2 s13923_7(wires_3480_6[3], addr_3480_6, addr_positional[55695:55692], addr_13923_7);

wire[31:0] addr_13924_7;

Selector_2 s13924_7(wires_3481_6[0], addr_3481_6, addr_positional[55699:55696], addr_13924_7);

wire[31:0] addr_13925_7;

Selector_2 s13925_7(wires_3481_6[1], addr_3481_6, addr_positional[55703:55700], addr_13925_7);

wire[31:0] addr_13926_7;

Selector_2 s13926_7(wires_3481_6[2], addr_3481_6, addr_positional[55707:55704], addr_13926_7);

wire[31:0] addr_13927_7;

Selector_2 s13927_7(wires_3481_6[3], addr_3481_6, addr_positional[55711:55708], addr_13927_7);

wire[31:0] addr_13928_7;

Selector_2 s13928_7(wires_3482_6[0], addr_3482_6, addr_positional[55715:55712], addr_13928_7);

wire[31:0] addr_13929_7;

Selector_2 s13929_7(wires_3482_6[1], addr_3482_6, addr_positional[55719:55716], addr_13929_7);

wire[31:0] addr_13930_7;

Selector_2 s13930_7(wires_3482_6[2], addr_3482_6, addr_positional[55723:55720], addr_13930_7);

wire[31:0] addr_13931_7;

Selector_2 s13931_7(wires_3482_6[3], addr_3482_6, addr_positional[55727:55724], addr_13931_7);

wire[31:0] addr_13932_7;

Selector_2 s13932_7(wires_3483_6[0], addr_3483_6, addr_positional[55731:55728], addr_13932_7);

wire[31:0] addr_13933_7;

Selector_2 s13933_7(wires_3483_6[1], addr_3483_6, addr_positional[55735:55732], addr_13933_7);

wire[31:0] addr_13934_7;

Selector_2 s13934_7(wires_3483_6[2], addr_3483_6, addr_positional[55739:55736], addr_13934_7);

wire[31:0] addr_13935_7;

Selector_2 s13935_7(wires_3483_6[3], addr_3483_6, addr_positional[55743:55740], addr_13935_7);

wire[31:0] addr_13936_7;

Selector_2 s13936_7(wires_3484_6[0], addr_3484_6, addr_positional[55747:55744], addr_13936_7);

wire[31:0] addr_13937_7;

Selector_2 s13937_7(wires_3484_6[1], addr_3484_6, addr_positional[55751:55748], addr_13937_7);

wire[31:0] addr_13938_7;

Selector_2 s13938_7(wires_3484_6[2], addr_3484_6, addr_positional[55755:55752], addr_13938_7);

wire[31:0] addr_13939_7;

Selector_2 s13939_7(wires_3484_6[3], addr_3484_6, addr_positional[55759:55756], addr_13939_7);

wire[31:0] addr_13940_7;

Selector_2 s13940_7(wires_3485_6[0], addr_3485_6, addr_positional[55763:55760], addr_13940_7);

wire[31:0] addr_13941_7;

Selector_2 s13941_7(wires_3485_6[1], addr_3485_6, addr_positional[55767:55764], addr_13941_7);

wire[31:0] addr_13942_7;

Selector_2 s13942_7(wires_3485_6[2], addr_3485_6, addr_positional[55771:55768], addr_13942_7);

wire[31:0] addr_13943_7;

Selector_2 s13943_7(wires_3485_6[3], addr_3485_6, addr_positional[55775:55772], addr_13943_7);

wire[31:0] addr_13944_7;

Selector_2 s13944_7(wires_3486_6[0], addr_3486_6, addr_positional[55779:55776], addr_13944_7);

wire[31:0] addr_13945_7;

Selector_2 s13945_7(wires_3486_6[1], addr_3486_6, addr_positional[55783:55780], addr_13945_7);

wire[31:0] addr_13946_7;

Selector_2 s13946_7(wires_3486_6[2], addr_3486_6, addr_positional[55787:55784], addr_13946_7);

wire[31:0] addr_13947_7;

Selector_2 s13947_7(wires_3486_6[3], addr_3486_6, addr_positional[55791:55788], addr_13947_7);

wire[31:0] addr_13948_7;

Selector_2 s13948_7(wires_3487_6[0], addr_3487_6, addr_positional[55795:55792], addr_13948_7);

wire[31:0] addr_13949_7;

Selector_2 s13949_7(wires_3487_6[1], addr_3487_6, addr_positional[55799:55796], addr_13949_7);

wire[31:0] addr_13950_7;

Selector_2 s13950_7(wires_3487_6[2], addr_3487_6, addr_positional[55803:55800], addr_13950_7);

wire[31:0] addr_13951_7;

Selector_2 s13951_7(wires_3487_6[3], addr_3487_6, addr_positional[55807:55804], addr_13951_7);

wire[31:0] addr_13952_7;

Selector_2 s13952_7(wires_3488_6[0], addr_3488_6, addr_positional[55811:55808], addr_13952_7);

wire[31:0] addr_13953_7;

Selector_2 s13953_7(wires_3488_6[1], addr_3488_6, addr_positional[55815:55812], addr_13953_7);

wire[31:0] addr_13954_7;

Selector_2 s13954_7(wires_3488_6[2], addr_3488_6, addr_positional[55819:55816], addr_13954_7);

wire[31:0] addr_13955_7;

Selector_2 s13955_7(wires_3488_6[3], addr_3488_6, addr_positional[55823:55820], addr_13955_7);

wire[31:0] addr_13956_7;

Selector_2 s13956_7(wires_3489_6[0], addr_3489_6, addr_positional[55827:55824], addr_13956_7);

wire[31:0] addr_13957_7;

Selector_2 s13957_7(wires_3489_6[1], addr_3489_6, addr_positional[55831:55828], addr_13957_7);

wire[31:0] addr_13958_7;

Selector_2 s13958_7(wires_3489_6[2], addr_3489_6, addr_positional[55835:55832], addr_13958_7);

wire[31:0] addr_13959_7;

Selector_2 s13959_7(wires_3489_6[3], addr_3489_6, addr_positional[55839:55836], addr_13959_7);

wire[31:0] addr_13960_7;

Selector_2 s13960_7(wires_3490_6[0], addr_3490_6, addr_positional[55843:55840], addr_13960_7);

wire[31:0] addr_13961_7;

Selector_2 s13961_7(wires_3490_6[1], addr_3490_6, addr_positional[55847:55844], addr_13961_7);

wire[31:0] addr_13962_7;

Selector_2 s13962_7(wires_3490_6[2], addr_3490_6, addr_positional[55851:55848], addr_13962_7);

wire[31:0] addr_13963_7;

Selector_2 s13963_7(wires_3490_6[3], addr_3490_6, addr_positional[55855:55852], addr_13963_7);

wire[31:0] addr_13964_7;

Selector_2 s13964_7(wires_3491_6[0], addr_3491_6, addr_positional[55859:55856], addr_13964_7);

wire[31:0] addr_13965_7;

Selector_2 s13965_7(wires_3491_6[1], addr_3491_6, addr_positional[55863:55860], addr_13965_7);

wire[31:0] addr_13966_7;

Selector_2 s13966_7(wires_3491_6[2], addr_3491_6, addr_positional[55867:55864], addr_13966_7);

wire[31:0] addr_13967_7;

Selector_2 s13967_7(wires_3491_6[3], addr_3491_6, addr_positional[55871:55868], addr_13967_7);

wire[31:0] addr_13968_7;

Selector_2 s13968_7(wires_3492_6[0], addr_3492_6, addr_positional[55875:55872], addr_13968_7);

wire[31:0] addr_13969_7;

Selector_2 s13969_7(wires_3492_6[1], addr_3492_6, addr_positional[55879:55876], addr_13969_7);

wire[31:0] addr_13970_7;

Selector_2 s13970_7(wires_3492_6[2], addr_3492_6, addr_positional[55883:55880], addr_13970_7);

wire[31:0] addr_13971_7;

Selector_2 s13971_7(wires_3492_6[3], addr_3492_6, addr_positional[55887:55884], addr_13971_7);

wire[31:0] addr_13972_7;

Selector_2 s13972_7(wires_3493_6[0], addr_3493_6, addr_positional[55891:55888], addr_13972_7);

wire[31:0] addr_13973_7;

Selector_2 s13973_7(wires_3493_6[1], addr_3493_6, addr_positional[55895:55892], addr_13973_7);

wire[31:0] addr_13974_7;

Selector_2 s13974_7(wires_3493_6[2], addr_3493_6, addr_positional[55899:55896], addr_13974_7);

wire[31:0] addr_13975_7;

Selector_2 s13975_7(wires_3493_6[3], addr_3493_6, addr_positional[55903:55900], addr_13975_7);

wire[31:0] addr_13976_7;

Selector_2 s13976_7(wires_3494_6[0], addr_3494_6, addr_positional[55907:55904], addr_13976_7);

wire[31:0] addr_13977_7;

Selector_2 s13977_7(wires_3494_6[1], addr_3494_6, addr_positional[55911:55908], addr_13977_7);

wire[31:0] addr_13978_7;

Selector_2 s13978_7(wires_3494_6[2], addr_3494_6, addr_positional[55915:55912], addr_13978_7);

wire[31:0] addr_13979_7;

Selector_2 s13979_7(wires_3494_6[3], addr_3494_6, addr_positional[55919:55916], addr_13979_7);

wire[31:0] addr_13980_7;

Selector_2 s13980_7(wires_3495_6[0], addr_3495_6, addr_positional[55923:55920], addr_13980_7);

wire[31:0] addr_13981_7;

Selector_2 s13981_7(wires_3495_6[1], addr_3495_6, addr_positional[55927:55924], addr_13981_7);

wire[31:0] addr_13982_7;

Selector_2 s13982_7(wires_3495_6[2], addr_3495_6, addr_positional[55931:55928], addr_13982_7);

wire[31:0] addr_13983_7;

Selector_2 s13983_7(wires_3495_6[3], addr_3495_6, addr_positional[55935:55932], addr_13983_7);

wire[31:0] addr_13984_7;

Selector_2 s13984_7(wires_3496_6[0], addr_3496_6, addr_positional[55939:55936], addr_13984_7);

wire[31:0] addr_13985_7;

Selector_2 s13985_7(wires_3496_6[1], addr_3496_6, addr_positional[55943:55940], addr_13985_7);

wire[31:0] addr_13986_7;

Selector_2 s13986_7(wires_3496_6[2], addr_3496_6, addr_positional[55947:55944], addr_13986_7);

wire[31:0] addr_13987_7;

Selector_2 s13987_7(wires_3496_6[3], addr_3496_6, addr_positional[55951:55948], addr_13987_7);

wire[31:0] addr_13988_7;

Selector_2 s13988_7(wires_3497_6[0], addr_3497_6, addr_positional[55955:55952], addr_13988_7);

wire[31:0] addr_13989_7;

Selector_2 s13989_7(wires_3497_6[1], addr_3497_6, addr_positional[55959:55956], addr_13989_7);

wire[31:0] addr_13990_7;

Selector_2 s13990_7(wires_3497_6[2], addr_3497_6, addr_positional[55963:55960], addr_13990_7);

wire[31:0] addr_13991_7;

Selector_2 s13991_7(wires_3497_6[3], addr_3497_6, addr_positional[55967:55964], addr_13991_7);

wire[31:0] addr_13992_7;

Selector_2 s13992_7(wires_3498_6[0], addr_3498_6, addr_positional[55971:55968], addr_13992_7);

wire[31:0] addr_13993_7;

Selector_2 s13993_7(wires_3498_6[1], addr_3498_6, addr_positional[55975:55972], addr_13993_7);

wire[31:0] addr_13994_7;

Selector_2 s13994_7(wires_3498_6[2], addr_3498_6, addr_positional[55979:55976], addr_13994_7);

wire[31:0] addr_13995_7;

Selector_2 s13995_7(wires_3498_6[3], addr_3498_6, addr_positional[55983:55980], addr_13995_7);

wire[31:0] addr_13996_7;

Selector_2 s13996_7(wires_3499_6[0], addr_3499_6, addr_positional[55987:55984], addr_13996_7);

wire[31:0] addr_13997_7;

Selector_2 s13997_7(wires_3499_6[1], addr_3499_6, addr_positional[55991:55988], addr_13997_7);

wire[31:0] addr_13998_7;

Selector_2 s13998_7(wires_3499_6[2], addr_3499_6, addr_positional[55995:55992], addr_13998_7);

wire[31:0] addr_13999_7;

Selector_2 s13999_7(wires_3499_6[3], addr_3499_6, addr_positional[55999:55996], addr_13999_7);

wire[31:0] addr_14000_7;

Selector_2 s14000_7(wires_3500_6[0], addr_3500_6, addr_positional[56003:56000], addr_14000_7);

wire[31:0] addr_14001_7;

Selector_2 s14001_7(wires_3500_6[1], addr_3500_6, addr_positional[56007:56004], addr_14001_7);

wire[31:0] addr_14002_7;

Selector_2 s14002_7(wires_3500_6[2], addr_3500_6, addr_positional[56011:56008], addr_14002_7);

wire[31:0] addr_14003_7;

Selector_2 s14003_7(wires_3500_6[3], addr_3500_6, addr_positional[56015:56012], addr_14003_7);

wire[31:0] addr_14004_7;

Selector_2 s14004_7(wires_3501_6[0], addr_3501_6, addr_positional[56019:56016], addr_14004_7);

wire[31:0] addr_14005_7;

Selector_2 s14005_7(wires_3501_6[1], addr_3501_6, addr_positional[56023:56020], addr_14005_7);

wire[31:0] addr_14006_7;

Selector_2 s14006_7(wires_3501_6[2], addr_3501_6, addr_positional[56027:56024], addr_14006_7);

wire[31:0] addr_14007_7;

Selector_2 s14007_7(wires_3501_6[3], addr_3501_6, addr_positional[56031:56028], addr_14007_7);

wire[31:0] addr_14008_7;

Selector_2 s14008_7(wires_3502_6[0], addr_3502_6, addr_positional[56035:56032], addr_14008_7);

wire[31:0] addr_14009_7;

Selector_2 s14009_7(wires_3502_6[1], addr_3502_6, addr_positional[56039:56036], addr_14009_7);

wire[31:0] addr_14010_7;

Selector_2 s14010_7(wires_3502_6[2], addr_3502_6, addr_positional[56043:56040], addr_14010_7);

wire[31:0] addr_14011_7;

Selector_2 s14011_7(wires_3502_6[3], addr_3502_6, addr_positional[56047:56044], addr_14011_7);

wire[31:0] addr_14012_7;

Selector_2 s14012_7(wires_3503_6[0], addr_3503_6, addr_positional[56051:56048], addr_14012_7);

wire[31:0] addr_14013_7;

Selector_2 s14013_7(wires_3503_6[1], addr_3503_6, addr_positional[56055:56052], addr_14013_7);

wire[31:0] addr_14014_7;

Selector_2 s14014_7(wires_3503_6[2], addr_3503_6, addr_positional[56059:56056], addr_14014_7);

wire[31:0] addr_14015_7;

Selector_2 s14015_7(wires_3503_6[3], addr_3503_6, addr_positional[56063:56060], addr_14015_7);

wire[31:0] addr_14016_7;

Selector_2 s14016_7(wires_3504_6[0], addr_3504_6, addr_positional[56067:56064], addr_14016_7);

wire[31:0] addr_14017_7;

Selector_2 s14017_7(wires_3504_6[1], addr_3504_6, addr_positional[56071:56068], addr_14017_7);

wire[31:0] addr_14018_7;

Selector_2 s14018_7(wires_3504_6[2], addr_3504_6, addr_positional[56075:56072], addr_14018_7);

wire[31:0] addr_14019_7;

Selector_2 s14019_7(wires_3504_6[3], addr_3504_6, addr_positional[56079:56076], addr_14019_7);

wire[31:0] addr_14020_7;

Selector_2 s14020_7(wires_3505_6[0], addr_3505_6, addr_positional[56083:56080], addr_14020_7);

wire[31:0] addr_14021_7;

Selector_2 s14021_7(wires_3505_6[1], addr_3505_6, addr_positional[56087:56084], addr_14021_7);

wire[31:0] addr_14022_7;

Selector_2 s14022_7(wires_3505_6[2], addr_3505_6, addr_positional[56091:56088], addr_14022_7);

wire[31:0] addr_14023_7;

Selector_2 s14023_7(wires_3505_6[3], addr_3505_6, addr_positional[56095:56092], addr_14023_7);

wire[31:0] addr_14024_7;

Selector_2 s14024_7(wires_3506_6[0], addr_3506_6, addr_positional[56099:56096], addr_14024_7);

wire[31:0] addr_14025_7;

Selector_2 s14025_7(wires_3506_6[1], addr_3506_6, addr_positional[56103:56100], addr_14025_7);

wire[31:0] addr_14026_7;

Selector_2 s14026_7(wires_3506_6[2], addr_3506_6, addr_positional[56107:56104], addr_14026_7);

wire[31:0] addr_14027_7;

Selector_2 s14027_7(wires_3506_6[3], addr_3506_6, addr_positional[56111:56108], addr_14027_7);

wire[31:0] addr_14028_7;

Selector_2 s14028_7(wires_3507_6[0], addr_3507_6, addr_positional[56115:56112], addr_14028_7);

wire[31:0] addr_14029_7;

Selector_2 s14029_7(wires_3507_6[1], addr_3507_6, addr_positional[56119:56116], addr_14029_7);

wire[31:0] addr_14030_7;

Selector_2 s14030_7(wires_3507_6[2], addr_3507_6, addr_positional[56123:56120], addr_14030_7);

wire[31:0] addr_14031_7;

Selector_2 s14031_7(wires_3507_6[3], addr_3507_6, addr_positional[56127:56124], addr_14031_7);

wire[31:0] addr_14032_7;

Selector_2 s14032_7(wires_3508_6[0], addr_3508_6, addr_positional[56131:56128], addr_14032_7);

wire[31:0] addr_14033_7;

Selector_2 s14033_7(wires_3508_6[1], addr_3508_6, addr_positional[56135:56132], addr_14033_7);

wire[31:0] addr_14034_7;

Selector_2 s14034_7(wires_3508_6[2], addr_3508_6, addr_positional[56139:56136], addr_14034_7);

wire[31:0] addr_14035_7;

Selector_2 s14035_7(wires_3508_6[3], addr_3508_6, addr_positional[56143:56140], addr_14035_7);

wire[31:0] addr_14036_7;

Selector_2 s14036_7(wires_3509_6[0], addr_3509_6, addr_positional[56147:56144], addr_14036_7);

wire[31:0] addr_14037_7;

Selector_2 s14037_7(wires_3509_6[1], addr_3509_6, addr_positional[56151:56148], addr_14037_7);

wire[31:0] addr_14038_7;

Selector_2 s14038_7(wires_3509_6[2], addr_3509_6, addr_positional[56155:56152], addr_14038_7);

wire[31:0] addr_14039_7;

Selector_2 s14039_7(wires_3509_6[3], addr_3509_6, addr_positional[56159:56156], addr_14039_7);

wire[31:0] addr_14040_7;

Selector_2 s14040_7(wires_3510_6[0], addr_3510_6, addr_positional[56163:56160], addr_14040_7);

wire[31:0] addr_14041_7;

Selector_2 s14041_7(wires_3510_6[1], addr_3510_6, addr_positional[56167:56164], addr_14041_7);

wire[31:0] addr_14042_7;

Selector_2 s14042_7(wires_3510_6[2], addr_3510_6, addr_positional[56171:56168], addr_14042_7);

wire[31:0] addr_14043_7;

Selector_2 s14043_7(wires_3510_6[3], addr_3510_6, addr_positional[56175:56172], addr_14043_7);

wire[31:0] addr_14044_7;

Selector_2 s14044_7(wires_3511_6[0], addr_3511_6, addr_positional[56179:56176], addr_14044_7);

wire[31:0] addr_14045_7;

Selector_2 s14045_7(wires_3511_6[1], addr_3511_6, addr_positional[56183:56180], addr_14045_7);

wire[31:0] addr_14046_7;

Selector_2 s14046_7(wires_3511_6[2], addr_3511_6, addr_positional[56187:56184], addr_14046_7);

wire[31:0] addr_14047_7;

Selector_2 s14047_7(wires_3511_6[3], addr_3511_6, addr_positional[56191:56188], addr_14047_7);

wire[31:0] addr_14048_7;

Selector_2 s14048_7(wires_3512_6[0], addr_3512_6, addr_positional[56195:56192], addr_14048_7);

wire[31:0] addr_14049_7;

Selector_2 s14049_7(wires_3512_6[1], addr_3512_6, addr_positional[56199:56196], addr_14049_7);

wire[31:0] addr_14050_7;

Selector_2 s14050_7(wires_3512_6[2], addr_3512_6, addr_positional[56203:56200], addr_14050_7);

wire[31:0] addr_14051_7;

Selector_2 s14051_7(wires_3512_6[3], addr_3512_6, addr_positional[56207:56204], addr_14051_7);

wire[31:0] addr_14052_7;

Selector_2 s14052_7(wires_3513_6[0], addr_3513_6, addr_positional[56211:56208], addr_14052_7);

wire[31:0] addr_14053_7;

Selector_2 s14053_7(wires_3513_6[1], addr_3513_6, addr_positional[56215:56212], addr_14053_7);

wire[31:0] addr_14054_7;

Selector_2 s14054_7(wires_3513_6[2], addr_3513_6, addr_positional[56219:56216], addr_14054_7);

wire[31:0] addr_14055_7;

Selector_2 s14055_7(wires_3513_6[3], addr_3513_6, addr_positional[56223:56220], addr_14055_7);

wire[31:0] addr_14056_7;

Selector_2 s14056_7(wires_3514_6[0], addr_3514_6, addr_positional[56227:56224], addr_14056_7);

wire[31:0] addr_14057_7;

Selector_2 s14057_7(wires_3514_6[1], addr_3514_6, addr_positional[56231:56228], addr_14057_7);

wire[31:0] addr_14058_7;

Selector_2 s14058_7(wires_3514_6[2], addr_3514_6, addr_positional[56235:56232], addr_14058_7);

wire[31:0] addr_14059_7;

Selector_2 s14059_7(wires_3514_6[3], addr_3514_6, addr_positional[56239:56236], addr_14059_7);

wire[31:0] addr_14060_7;

Selector_2 s14060_7(wires_3515_6[0], addr_3515_6, addr_positional[56243:56240], addr_14060_7);

wire[31:0] addr_14061_7;

Selector_2 s14061_7(wires_3515_6[1], addr_3515_6, addr_positional[56247:56244], addr_14061_7);

wire[31:0] addr_14062_7;

Selector_2 s14062_7(wires_3515_6[2], addr_3515_6, addr_positional[56251:56248], addr_14062_7);

wire[31:0] addr_14063_7;

Selector_2 s14063_7(wires_3515_6[3], addr_3515_6, addr_positional[56255:56252], addr_14063_7);

wire[31:0] addr_14064_7;

Selector_2 s14064_7(wires_3516_6[0], addr_3516_6, addr_positional[56259:56256], addr_14064_7);

wire[31:0] addr_14065_7;

Selector_2 s14065_7(wires_3516_6[1], addr_3516_6, addr_positional[56263:56260], addr_14065_7);

wire[31:0] addr_14066_7;

Selector_2 s14066_7(wires_3516_6[2], addr_3516_6, addr_positional[56267:56264], addr_14066_7);

wire[31:0] addr_14067_7;

Selector_2 s14067_7(wires_3516_6[3], addr_3516_6, addr_positional[56271:56268], addr_14067_7);

wire[31:0] addr_14068_7;

Selector_2 s14068_7(wires_3517_6[0], addr_3517_6, addr_positional[56275:56272], addr_14068_7);

wire[31:0] addr_14069_7;

Selector_2 s14069_7(wires_3517_6[1], addr_3517_6, addr_positional[56279:56276], addr_14069_7);

wire[31:0] addr_14070_7;

Selector_2 s14070_7(wires_3517_6[2], addr_3517_6, addr_positional[56283:56280], addr_14070_7);

wire[31:0] addr_14071_7;

Selector_2 s14071_7(wires_3517_6[3], addr_3517_6, addr_positional[56287:56284], addr_14071_7);

wire[31:0] addr_14072_7;

Selector_2 s14072_7(wires_3518_6[0], addr_3518_6, addr_positional[56291:56288], addr_14072_7);

wire[31:0] addr_14073_7;

Selector_2 s14073_7(wires_3518_6[1], addr_3518_6, addr_positional[56295:56292], addr_14073_7);

wire[31:0] addr_14074_7;

Selector_2 s14074_7(wires_3518_6[2], addr_3518_6, addr_positional[56299:56296], addr_14074_7);

wire[31:0] addr_14075_7;

Selector_2 s14075_7(wires_3518_6[3], addr_3518_6, addr_positional[56303:56300], addr_14075_7);

wire[31:0] addr_14076_7;

Selector_2 s14076_7(wires_3519_6[0], addr_3519_6, addr_positional[56307:56304], addr_14076_7);

wire[31:0] addr_14077_7;

Selector_2 s14077_7(wires_3519_6[1], addr_3519_6, addr_positional[56311:56308], addr_14077_7);

wire[31:0] addr_14078_7;

Selector_2 s14078_7(wires_3519_6[2], addr_3519_6, addr_positional[56315:56312], addr_14078_7);

wire[31:0] addr_14079_7;

Selector_2 s14079_7(wires_3519_6[3], addr_3519_6, addr_positional[56319:56316], addr_14079_7);

wire[31:0] addr_14080_7;

Selector_2 s14080_7(wires_3520_6[0], addr_3520_6, addr_positional[56323:56320], addr_14080_7);

wire[31:0] addr_14081_7;

Selector_2 s14081_7(wires_3520_6[1], addr_3520_6, addr_positional[56327:56324], addr_14081_7);

wire[31:0] addr_14082_7;

Selector_2 s14082_7(wires_3520_6[2], addr_3520_6, addr_positional[56331:56328], addr_14082_7);

wire[31:0] addr_14083_7;

Selector_2 s14083_7(wires_3520_6[3], addr_3520_6, addr_positional[56335:56332], addr_14083_7);

wire[31:0] addr_14084_7;

Selector_2 s14084_7(wires_3521_6[0], addr_3521_6, addr_positional[56339:56336], addr_14084_7);

wire[31:0] addr_14085_7;

Selector_2 s14085_7(wires_3521_6[1], addr_3521_6, addr_positional[56343:56340], addr_14085_7);

wire[31:0] addr_14086_7;

Selector_2 s14086_7(wires_3521_6[2], addr_3521_6, addr_positional[56347:56344], addr_14086_7);

wire[31:0] addr_14087_7;

Selector_2 s14087_7(wires_3521_6[3], addr_3521_6, addr_positional[56351:56348], addr_14087_7);

wire[31:0] addr_14088_7;

Selector_2 s14088_7(wires_3522_6[0], addr_3522_6, addr_positional[56355:56352], addr_14088_7);

wire[31:0] addr_14089_7;

Selector_2 s14089_7(wires_3522_6[1], addr_3522_6, addr_positional[56359:56356], addr_14089_7);

wire[31:0] addr_14090_7;

Selector_2 s14090_7(wires_3522_6[2], addr_3522_6, addr_positional[56363:56360], addr_14090_7);

wire[31:0] addr_14091_7;

Selector_2 s14091_7(wires_3522_6[3], addr_3522_6, addr_positional[56367:56364], addr_14091_7);

wire[31:0] addr_14092_7;

Selector_2 s14092_7(wires_3523_6[0], addr_3523_6, addr_positional[56371:56368], addr_14092_7);

wire[31:0] addr_14093_7;

Selector_2 s14093_7(wires_3523_6[1], addr_3523_6, addr_positional[56375:56372], addr_14093_7);

wire[31:0] addr_14094_7;

Selector_2 s14094_7(wires_3523_6[2], addr_3523_6, addr_positional[56379:56376], addr_14094_7);

wire[31:0] addr_14095_7;

Selector_2 s14095_7(wires_3523_6[3], addr_3523_6, addr_positional[56383:56380], addr_14095_7);

wire[31:0] addr_14096_7;

Selector_2 s14096_7(wires_3524_6[0], addr_3524_6, addr_positional[56387:56384], addr_14096_7);

wire[31:0] addr_14097_7;

Selector_2 s14097_7(wires_3524_6[1], addr_3524_6, addr_positional[56391:56388], addr_14097_7);

wire[31:0] addr_14098_7;

Selector_2 s14098_7(wires_3524_6[2], addr_3524_6, addr_positional[56395:56392], addr_14098_7);

wire[31:0] addr_14099_7;

Selector_2 s14099_7(wires_3524_6[3], addr_3524_6, addr_positional[56399:56396], addr_14099_7);

wire[31:0] addr_14100_7;

Selector_2 s14100_7(wires_3525_6[0], addr_3525_6, addr_positional[56403:56400], addr_14100_7);

wire[31:0] addr_14101_7;

Selector_2 s14101_7(wires_3525_6[1], addr_3525_6, addr_positional[56407:56404], addr_14101_7);

wire[31:0] addr_14102_7;

Selector_2 s14102_7(wires_3525_6[2], addr_3525_6, addr_positional[56411:56408], addr_14102_7);

wire[31:0] addr_14103_7;

Selector_2 s14103_7(wires_3525_6[3], addr_3525_6, addr_positional[56415:56412], addr_14103_7);

wire[31:0] addr_14104_7;

Selector_2 s14104_7(wires_3526_6[0], addr_3526_6, addr_positional[56419:56416], addr_14104_7);

wire[31:0] addr_14105_7;

Selector_2 s14105_7(wires_3526_6[1], addr_3526_6, addr_positional[56423:56420], addr_14105_7);

wire[31:0] addr_14106_7;

Selector_2 s14106_7(wires_3526_6[2], addr_3526_6, addr_positional[56427:56424], addr_14106_7);

wire[31:0] addr_14107_7;

Selector_2 s14107_7(wires_3526_6[3], addr_3526_6, addr_positional[56431:56428], addr_14107_7);

wire[31:0] addr_14108_7;

Selector_2 s14108_7(wires_3527_6[0], addr_3527_6, addr_positional[56435:56432], addr_14108_7);

wire[31:0] addr_14109_7;

Selector_2 s14109_7(wires_3527_6[1], addr_3527_6, addr_positional[56439:56436], addr_14109_7);

wire[31:0] addr_14110_7;

Selector_2 s14110_7(wires_3527_6[2], addr_3527_6, addr_positional[56443:56440], addr_14110_7);

wire[31:0] addr_14111_7;

Selector_2 s14111_7(wires_3527_6[3], addr_3527_6, addr_positional[56447:56444], addr_14111_7);

wire[31:0] addr_14112_7;

Selector_2 s14112_7(wires_3528_6[0], addr_3528_6, addr_positional[56451:56448], addr_14112_7);

wire[31:0] addr_14113_7;

Selector_2 s14113_7(wires_3528_6[1], addr_3528_6, addr_positional[56455:56452], addr_14113_7);

wire[31:0] addr_14114_7;

Selector_2 s14114_7(wires_3528_6[2], addr_3528_6, addr_positional[56459:56456], addr_14114_7);

wire[31:0] addr_14115_7;

Selector_2 s14115_7(wires_3528_6[3], addr_3528_6, addr_positional[56463:56460], addr_14115_7);

wire[31:0] addr_14116_7;

Selector_2 s14116_7(wires_3529_6[0], addr_3529_6, addr_positional[56467:56464], addr_14116_7);

wire[31:0] addr_14117_7;

Selector_2 s14117_7(wires_3529_6[1], addr_3529_6, addr_positional[56471:56468], addr_14117_7);

wire[31:0] addr_14118_7;

Selector_2 s14118_7(wires_3529_6[2], addr_3529_6, addr_positional[56475:56472], addr_14118_7);

wire[31:0] addr_14119_7;

Selector_2 s14119_7(wires_3529_6[3], addr_3529_6, addr_positional[56479:56476], addr_14119_7);

wire[31:0] addr_14120_7;

Selector_2 s14120_7(wires_3530_6[0], addr_3530_6, addr_positional[56483:56480], addr_14120_7);

wire[31:0] addr_14121_7;

Selector_2 s14121_7(wires_3530_6[1], addr_3530_6, addr_positional[56487:56484], addr_14121_7);

wire[31:0] addr_14122_7;

Selector_2 s14122_7(wires_3530_6[2], addr_3530_6, addr_positional[56491:56488], addr_14122_7);

wire[31:0] addr_14123_7;

Selector_2 s14123_7(wires_3530_6[3], addr_3530_6, addr_positional[56495:56492], addr_14123_7);

wire[31:0] addr_14124_7;

Selector_2 s14124_7(wires_3531_6[0], addr_3531_6, addr_positional[56499:56496], addr_14124_7);

wire[31:0] addr_14125_7;

Selector_2 s14125_7(wires_3531_6[1], addr_3531_6, addr_positional[56503:56500], addr_14125_7);

wire[31:0] addr_14126_7;

Selector_2 s14126_7(wires_3531_6[2], addr_3531_6, addr_positional[56507:56504], addr_14126_7);

wire[31:0] addr_14127_7;

Selector_2 s14127_7(wires_3531_6[3], addr_3531_6, addr_positional[56511:56508], addr_14127_7);

wire[31:0] addr_14128_7;

Selector_2 s14128_7(wires_3532_6[0], addr_3532_6, addr_positional[56515:56512], addr_14128_7);

wire[31:0] addr_14129_7;

Selector_2 s14129_7(wires_3532_6[1], addr_3532_6, addr_positional[56519:56516], addr_14129_7);

wire[31:0] addr_14130_7;

Selector_2 s14130_7(wires_3532_6[2], addr_3532_6, addr_positional[56523:56520], addr_14130_7);

wire[31:0] addr_14131_7;

Selector_2 s14131_7(wires_3532_6[3], addr_3532_6, addr_positional[56527:56524], addr_14131_7);

wire[31:0] addr_14132_7;

Selector_2 s14132_7(wires_3533_6[0], addr_3533_6, addr_positional[56531:56528], addr_14132_7);

wire[31:0] addr_14133_7;

Selector_2 s14133_7(wires_3533_6[1], addr_3533_6, addr_positional[56535:56532], addr_14133_7);

wire[31:0] addr_14134_7;

Selector_2 s14134_7(wires_3533_6[2], addr_3533_6, addr_positional[56539:56536], addr_14134_7);

wire[31:0] addr_14135_7;

Selector_2 s14135_7(wires_3533_6[3], addr_3533_6, addr_positional[56543:56540], addr_14135_7);

wire[31:0] addr_14136_7;

Selector_2 s14136_7(wires_3534_6[0], addr_3534_6, addr_positional[56547:56544], addr_14136_7);

wire[31:0] addr_14137_7;

Selector_2 s14137_7(wires_3534_6[1], addr_3534_6, addr_positional[56551:56548], addr_14137_7);

wire[31:0] addr_14138_7;

Selector_2 s14138_7(wires_3534_6[2], addr_3534_6, addr_positional[56555:56552], addr_14138_7);

wire[31:0] addr_14139_7;

Selector_2 s14139_7(wires_3534_6[3], addr_3534_6, addr_positional[56559:56556], addr_14139_7);

wire[31:0] addr_14140_7;

Selector_2 s14140_7(wires_3535_6[0], addr_3535_6, addr_positional[56563:56560], addr_14140_7);

wire[31:0] addr_14141_7;

Selector_2 s14141_7(wires_3535_6[1], addr_3535_6, addr_positional[56567:56564], addr_14141_7);

wire[31:0] addr_14142_7;

Selector_2 s14142_7(wires_3535_6[2], addr_3535_6, addr_positional[56571:56568], addr_14142_7);

wire[31:0] addr_14143_7;

Selector_2 s14143_7(wires_3535_6[3], addr_3535_6, addr_positional[56575:56572], addr_14143_7);

wire[31:0] addr_14144_7;

Selector_2 s14144_7(wires_3536_6[0], addr_3536_6, addr_positional[56579:56576], addr_14144_7);

wire[31:0] addr_14145_7;

Selector_2 s14145_7(wires_3536_6[1], addr_3536_6, addr_positional[56583:56580], addr_14145_7);

wire[31:0] addr_14146_7;

Selector_2 s14146_7(wires_3536_6[2], addr_3536_6, addr_positional[56587:56584], addr_14146_7);

wire[31:0] addr_14147_7;

Selector_2 s14147_7(wires_3536_6[3], addr_3536_6, addr_positional[56591:56588], addr_14147_7);

wire[31:0] addr_14148_7;

Selector_2 s14148_7(wires_3537_6[0], addr_3537_6, addr_positional[56595:56592], addr_14148_7);

wire[31:0] addr_14149_7;

Selector_2 s14149_7(wires_3537_6[1], addr_3537_6, addr_positional[56599:56596], addr_14149_7);

wire[31:0] addr_14150_7;

Selector_2 s14150_7(wires_3537_6[2], addr_3537_6, addr_positional[56603:56600], addr_14150_7);

wire[31:0] addr_14151_7;

Selector_2 s14151_7(wires_3537_6[3], addr_3537_6, addr_positional[56607:56604], addr_14151_7);

wire[31:0] addr_14152_7;

Selector_2 s14152_7(wires_3538_6[0], addr_3538_6, addr_positional[56611:56608], addr_14152_7);

wire[31:0] addr_14153_7;

Selector_2 s14153_7(wires_3538_6[1], addr_3538_6, addr_positional[56615:56612], addr_14153_7);

wire[31:0] addr_14154_7;

Selector_2 s14154_7(wires_3538_6[2], addr_3538_6, addr_positional[56619:56616], addr_14154_7);

wire[31:0] addr_14155_7;

Selector_2 s14155_7(wires_3538_6[3], addr_3538_6, addr_positional[56623:56620], addr_14155_7);

wire[31:0] addr_14156_7;

Selector_2 s14156_7(wires_3539_6[0], addr_3539_6, addr_positional[56627:56624], addr_14156_7);

wire[31:0] addr_14157_7;

Selector_2 s14157_7(wires_3539_6[1], addr_3539_6, addr_positional[56631:56628], addr_14157_7);

wire[31:0] addr_14158_7;

Selector_2 s14158_7(wires_3539_6[2], addr_3539_6, addr_positional[56635:56632], addr_14158_7);

wire[31:0] addr_14159_7;

Selector_2 s14159_7(wires_3539_6[3], addr_3539_6, addr_positional[56639:56636], addr_14159_7);

wire[31:0] addr_14160_7;

Selector_2 s14160_7(wires_3540_6[0], addr_3540_6, addr_positional[56643:56640], addr_14160_7);

wire[31:0] addr_14161_7;

Selector_2 s14161_7(wires_3540_6[1], addr_3540_6, addr_positional[56647:56644], addr_14161_7);

wire[31:0] addr_14162_7;

Selector_2 s14162_7(wires_3540_6[2], addr_3540_6, addr_positional[56651:56648], addr_14162_7);

wire[31:0] addr_14163_7;

Selector_2 s14163_7(wires_3540_6[3], addr_3540_6, addr_positional[56655:56652], addr_14163_7);

wire[31:0] addr_14164_7;

Selector_2 s14164_7(wires_3541_6[0], addr_3541_6, addr_positional[56659:56656], addr_14164_7);

wire[31:0] addr_14165_7;

Selector_2 s14165_7(wires_3541_6[1], addr_3541_6, addr_positional[56663:56660], addr_14165_7);

wire[31:0] addr_14166_7;

Selector_2 s14166_7(wires_3541_6[2], addr_3541_6, addr_positional[56667:56664], addr_14166_7);

wire[31:0] addr_14167_7;

Selector_2 s14167_7(wires_3541_6[3], addr_3541_6, addr_positional[56671:56668], addr_14167_7);

wire[31:0] addr_14168_7;

Selector_2 s14168_7(wires_3542_6[0], addr_3542_6, addr_positional[56675:56672], addr_14168_7);

wire[31:0] addr_14169_7;

Selector_2 s14169_7(wires_3542_6[1], addr_3542_6, addr_positional[56679:56676], addr_14169_7);

wire[31:0] addr_14170_7;

Selector_2 s14170_7(wires_3542_6[2], addr_3542_6, addr_positional[56683:56680], addr_14170_7);

wire[31:0] addr_14171_7;

Selector_2 s14171_7(wires_3542_6[3], addr_3542_6, addr_positional[56687:56684], addr_14171_7);

wire[31:0] addr_14172_7;

Selector_2 s14172_7(wires_3543_6[0], addr_3543_6, addr_positional[56691:56688], addr_14172_7);

wire[31:0] addr_14173_7;

Selector_2 s14173_7(wires_3543_6[1], addr_3543_6, addr_positional[56695:56692], addr_14173_7);

wire[31:0] addr_14174_7;

Selector_2 s14174_7(wires_3543_6[2], addr_3543_6, addr_positional[56699:56696], addr_14174_7);

wire[31:0] addr_14175_7;

Selector_2 s14175_7(wires_3543_6[3], addr_3543_6, addr_positional[56703:56700], addr_14175_7);

wire[31:0] addr_14176_7;

Selector_2 s14176_7(wires_3544_6[0], addr_3544_6, addr_positional[56707:56704], addr_14176_7);

wire[31:0] addr_14177_7;

Selector_2 s14177_7(wires_3544_6[1], addr_3544_6, addr_positional[56711:56708], addr_14177_7);

wire[31:0] addr_14178_7;

Selector_2 s14178_7(wires_3544_6[2], addr_3544_6, addr_positional[56715:56712], addr_14178_7);

wire[31:0] addr_14179_7;

Selector_2 s14179_7(wires_3544_6[3], addr_3544_6, addr_positional[56719:56716], addr_14179_7);

wire[31:0] addr_14180_7;

Selector_2 s14180_7(wires_3545_6[0], addr_3545_6, addr_positional[56723:56720], addr_14180_7);

wire[31:0] addr_14181_7;

Selector_2 s14181_7(wires_3545_6[1], addr_3545_6, addr_positional[56727:56724], addr_14181_7);

wire[31:0] addr_14182_7;

Selector_2 s14182_7(wires_3545_6[2], addr_3545_6, addr_positional[56731:56728], addr_14182_7);

wire[31:0] addr_14183_7;

Selector_2 s14183_7(wires_3545_6[3], addr_3545_6, addr_positional[56735:56732], addr_14183_7);

wire[31:0] addr_14184_7;

Selector_2 s14184_7(wires_3546_6[0], addr_3546_6, addr_positional[56739:56736], addr_14184_7);

wire[31:0] addr_14185_7;

Selector_2 s14185_7(wires_3546_6[1], addr_3546_6, addr_positional[56743:56740], addr_14185_7);

wire[31:0] addr_14186_7;

Selector_2 s14186_7(wires_3546_6[2], addr_3546_6, addr_positional[56747:56744], addr_14186_7);

wire[31:0] addr_14187_7;

Selector_2 s14187_7(wires_3546_6[3], addr_3546_6, addr_positional[56751:56748], addr_14187_7);

wire[31:0] addr_14188_7;

Selector_2 s14188_7(wires_3547_6[0], addr_3547_6, addr_positional[56755:56752], addr_14188_7);

wire[31:0] addr_14189_7;

Selector_2 s14189_7(wires_3547_6[1], addr_3547_6, addr_positional[56759:56756], addr_14189_7);

wire[31:0] addr_14190_7;

Selector_2 s14190_7(wires_3547_6[2], addr_3547_6, addr_positional[56763:56760], addr_14190_7);

wire[31:0] addr_14191_7;

Selector_2 s14191_7(wires_3547_6[3], addr_3547_6, addr_positional[56767:56764], addr_14191_7);

wire[31:0] addr_14192_7;

Selector_2 s14192_7(wires_3548_6[0], addr_3548_6, addr_positional[56771:56768], addr_14192_7);

wire[31:0] addr_14193_7;

Selector_2 s14193_7(wires_3548_6[1], addr_3548_6, addr_positional[56775:56772], addr_14193_7);

wire[31:0] addr_14194_7;

Selector_2 s14194_7(wires_3548_6[2], addr_3548_6, addr_positional[56779:56776], addr_14194_7);

wire[31:0] addr_14195_7;

Selector_2 s14195_7(wires_3548_6[3], addr_3548_6, addr_positional[56783:56780], addr_14195_7);

wire[31:0] addr_14196_7;

Selector_2 s14196_7(wires_3549_6[0], addr_3549_6, addr_positional[56787:56784], addr_14196_7);

wire[31:0] addr_14197_7;

Selector_2 s14197_7(wires_3549_6[1], addr_3549_6, addr_positional[56791:56788], addr_14197_7);

wire[31:0] addr_14198_7;

Selector_2 s14198_7(wires_3549_6[2], addr_3549_6, addr_positional[56795:56792], addr_14198_7);

wire[31:0] addr_14199_7;

Selector_2 s14199_7(wires_3549_6[3], addr_3549_6, addr_positional[56799:56796], addr_14199_7);

wire[31:0] addr_14200_7;

Selector_2 s14200_7(wires_3550_6[0], addr_3550_6, addr_positional[56803:56800], addr_14200_7);

wire[31:0] addr_14201_7;

Selector_2 s14201_7(wires_3550_6[1], addr_3550_6, addr_positional[56807:56804], addr_14201_7);

wire[31:0] addr_14202_7;

Selector_2 s14202_7(wires_3550_6[2], addr_3550_6, addr_positional[56811:56808], addr_14202_7);

wire[31:0] addr_14203_7;

Selector_2 s14203_7(wires_3550_6[3], addr_3550_6, addr_positional[56815:56812], addr_14203_7);

wire[31:0] addr_14204_7;

Selector_2 s14204_7(wires_3551_6[0], addr_3551_6, addr_positional[56819:56816], addr_14204_7);

wire[31:0] addr_14205_7;

Selector_2 s14205_7(wires_3551_6[1], addr_3551_6, addr_positional[56823:56820], addr_14205_7);

wire[31:0] addr_14206_7;

Selector_2 s14206_7(wires_3551_6[2], addr_3551_6, addr_positional[56827:56824], addr_14206_7);

wire[31:0] addr_14207_7;

Selector_2 s14207_7(wires_3551_6[3], addr_3551_6, addr_positional[56831:56828], addr_14207_7);

wire[31:0] addr_14208_7;

Selector_2 s14208_7(wires_3552_6[0], addr_3552_6, addr_positional[56835:56832], addr_14208_7);

wire[31:0] addr_14209_7;

Selector_2 s14209_7(wires_3552_6[1], addr_3552_6, addr_positional[56839:56836], addr_14209_7);

wire[31:0] addr_14210_7;

Selector_2 s14210_7(wires_3552_6[2], addr_3552_6, addr_positional[56843:56840], addr_14210_7);

wire[31:0] addr_14211_7;

Selector_2 s14211_7(wires_3552_6[3], addr_3552_6, addr_positional[56847:56844], addr_14211_7);

wire[31:0] addr_14212_7;

Selector_2 s14212_7(wires_3553_6[0], addr_3553_6, addr_positional[56851:56848], addr_14212_7);

wire[31:0] addr_14213_7;

Selector_2 s14213_7(wires_3553_6[1], addr_3553_6, addr_positional[56855:56852], addr_14213_7);

wire[31:0] addr_14214_7;

Selector_2 s14214_7(wires_3553_6[2], addr_3553_6, addr_positional[56859:56856], addr_14214_7);

wire[31:0] addr_14215_7;

Selector_2 s14215_7(wires_3553_6[3], addr_3553_6, addr_positional[56863:56860], addr_14215_7);

wire[31:0] addr_14216_7;

Selector_2 s14216_7(wires_3554_6[0], addr_3554_6, addr_positional[56867:56864], addr_14216_7);

wire[31:0] addr_14217_7;

Selector_2 s14217_7(wires_3554_6[1], addr_3554_6, addr_positional[56871:56868], addr_14217_7);

wire[31:0] addr_14218_7;

Selector_2 s14218_7(wires_3554_6[2], addr_3554_6, addr_positional[56875:56872], addr_14218_7);

wire[31:0] addr_14219_7;

Selector_2 s14219_7(wires_3554_6[3], addr_3554_6, addr_positional[56879:56876], addr_14219_7);

wire[31:0] addr_14220_7;

Selector_2 s14220_7(wires_3555_6[0], addr_3555_6, addr_positional[56883:56880], addr_14220_7);

wire[31:0] addr_14221_7;

Selector_2 s14221_7(wires_3555_6[1], addr_3555_6, addr_positional[56887:56884], addr_14221_7);

wire[31:0] addr_14222_7;

Selector_2 s14222_7(wires_3555_6[2], addr_3555_6, addr_positional[56891:56888], addr_14222_7);

wire[31:0] addr_14223_7;

Selector_2 s14223_7(wires_3555_6[3], addr_3555_6, addr_positional[56895:56892], addr_14223_7);

wire[31:0] addr_14224_7;

Selector_2 s14224_7(wires_3556_6[0], addr_3556_6, addr_positional[56899:56896], addr_14224_7);

wire[31:0] addr_14225_7;

Selector_2 s14225_7(wires_3556_6[1], addr_3556_6, addr_positional[56903:56900], addr_14225_7);

wire[31:0] addr_14226_7;

Selector_2 s14226_7(wires_3556_6[2], addr_3556_6, addr_positional[56907:56904], addr_14226_7);

wire[31:0] addr_14227_7;

Selector_2 s14227_7(wires_3556_6[3], addr_3556_6, addr_positional[56911:56908], addr_14227_7);

wire[31:0] addr_14228_7;

Selector_2 s14228_7(wires_3557_6[0], addr_3557_6, addr_positional[56915:56912], addr_14228_7);

wire[31:0] addr_14229_7;

Selector_2 s14229_7(wires_3557_6[1], addr_3557_6, addr_positional[56919:56916], addr_14229_7);

wire[31:0] addr_14230_7;

Selector_2 s14230_7(wires_3557_6[2], addr_3557_6, addr_positional[56923:56920], addr_14230_7);

wire[31:0] addr_14231_7;

Selector_2 s14231_7(wires_3557_6[3], addr_3557_6, addr_positional[56927:56924], addr_14231_7);

wire[31:0] addr_14232_7;

Selector_2 s14232_7(wires_3558_6[0], addr_3558_6, addr_positional[56931:56928], addr_14232_7);

wire[31:0] addr_14233_7;

Selector_2 s14233_7(wires_3558_6[1], addr_3558_6, addr_positional[56935:56932], addr_14233_7);

wire[31:0] addr_14234_7;

Selector_2 s14234_7(wires_3558_6[2], addr_3558_6, addr_positional[56939:56936], addr_14234_7);

wire[31:0] addr_14235_7;

Selector_2 s14235_7(wires_3558_6[3], addr_3558_6, addr_positional[56943:56940], addr_14235_7);

wire[31:0] addr_14236_7;

Selector_2 s14236_7(wires_3559_6[0], addr_3559_6, addr_positional[56947:56944], addr_14236_7);

wire[31:0] addr_14237_7;

Selector_2 s14237_7(wires_3559_6[1], addr_3559_6, addr_positional[56951:56948], addr_14237_7);

wire[31:0] addr_14238_7;

Selector_2 s14238_7(wires_3559_6[2], addr_3559_6, addr_positional[56955:56952], addr_14238_7);

wire[31:0] addr_14239_7;

Selector_2 s14239_7(wires_3559_6[3], addr_3559_6, addr_positional[56959:56956], addr_14239_7);

wire[31:0] addr_14240_7;

Selector_2 s14240_7(wires_3560_6[0], addr_3560_6, addr_positional[56963:56960], addr_14240_7);

wire[31:0] addr_14241_7;

Selector_2 s14241_7(wires_3560_6[1], addr_3560_6, addr_positional[56967:56964], addr_14241_7);

wire[31:0] addr_14242_7;

Selector_2 s14242_7(wires_3560_6[2], addr_3560_6, addr_positional[56971:56968], addr_14242_7);

wire[31:0] addr_14243_7;

Selector_2 s14243_7(wires_3560_6[3], addr_3560_6, addr_positional[56975:56972], addr_14243_7);

wire[31:0] addr_14244_7;

Selector_2 s14244_7(wires_3561_6[0], addr_3561_6, addr_positional[56979:56976], addr_14244_7);

wire[31:0] addr_14245_7;

Selector_2 s14245_7(wires_3561_6[1], addr_3561_6, addr_positional[56983:56980], addr_14245_7);

wire[31:0] addr_14246_7;

Selector_2 s14246_7(wires_3561_6[2], addr_3561_6, addr_positional[56987:56984], addr_14246_7);

wire[31:0] addr_14247_7;

Selector_2 s14247_7(wires_3561_6[3], addr_3561_6, addr_positional[56991:56988], addr_14247_7);

wire[31:0] addr_14248_7;

Selector_2 s14248_7(wires_3562_6[0], addr_3562_6, addr_positional[56995:56992], addr_14248_7);

wire[31:0] addr_14249_7;

Selector_2 s14249_7(wires_3562_6[1], addr_3562_6, addr_positional[56999:56996], addr_14249_7);

wire[31:0] addr_14250_7;

Selector_2 s14250_7(wires_3562_6[2], addr_3562_6, addr_positional[57003:57000], addr_14250_7);

wire[31:0] addr_14251_7;

Selector_2 s14251_7(wires_3562_6[3], addr_3562_6, addr_positional[57007:57004], addr_14251_7);

wire[31:0] addr_14252_7;

Selector_2 s14252_7(wires_3563_6[0], addr_3563_6, addr_positional[57011:57008], addr_14252_7);

wire[31:0] addr_14253_7;

Selector_2 s14253_7(wires_3563_6[1], addr_3563_6, addr_positional[57015:57012], addr_14253_7);

wire[31:0] addr_14254_7;

Selector_2 s14254_7(wires_3563_6[2], addr_3563_6, addr_positional[57019:57016], addr_14254_7);

wire[31:0] addr_14255_7;

Selector_2 s14255_7(wires_3563_6[3], addr_3563_6, addr_positional[57023:57020], addr_14255_7);

wire[31:0] addr_14256_7;

Selector_2 s14256_7(wires_3564_6[0], addr_3564_6, addr_positional[57027:57024], addr_14256_7);

wire[31:0] addr_14257_7;

Selector_2 s14257_7(wires_3564_6[1], addr_3564_6, addr_positional[57031:57028], addr_14257_7);

wire[31:0] addr_14258_7;

Selector_2 s14258_7(wires_3564_6[2], addr_3564_6, addr_positional[57035:57032], addr_14258_7);

wire[31:0] addr_14259_7;

Selector_2 s14259_7(wires_3564_6[3], addr_3564_6, addr_positional[57039:57036], addr_14259_7);

wire[31:0] addr_14260_7;

Selector_2 s14260_7(wires_3565_6[0], addr_3565_6, addr_positional[57043:57040], addr_14260_7);

wire[31:0] addr_14261_7;

Selector_2 s14261_7(wires_3565_6[1], addr_3565_6, addr_positional[57047:57044], addr_14261_7);

wire[31:0] addr_14262_7;

Selector_2 s14262_7(wires_3565_6[2], addr_3565_6, addr_positional[57051:57048], addr_14262_7);

wire[31:0] addr_14263_7;

Selector_2 s14263_7(wires_3565_6[3], addr_3565_6, addr_positional[57055:57052], addr_14263_7);

wire[31:0] addr_14264_7;

Selector_2 s14264_7(wires_3566_6[0], addr_3566_6, addr_positional[57059:57056], addr_14264_7);

wire[31:0] addr_14265_7;

Selector_2 s14265_7(wires_3566_6[1], addr_3566_6, addr_positional[57063:57060], addr_14265_7);

wire[31:0] addr_14266_7;

Selector_2 s14266_7(wires_3566_6[2], addr_3566_6, addr_positional[57067:57064], addr_14266_7);

wire[31:0] addr_14267_7;

Selector_2 s14267_7(wires_3566_6[3], addr_3566_6, addr_positional[57071:57068], addr_14267_7);

wire[31:0] addr_14268_7;

Selector_2 s14268_7(wires_3567_6[0], addr_3567_6, addr_positional[57075:57072], addr_14268_7);

wire[31:0] addr_14269_7;

Selector_2 s14269_7(wires_3567_6[1], addr_3567_6, addr_positional[57079:57076], addr_14269_7);

wire[31:0] addr_14270_7;

Selector_2 s14270_7(wires_3567_6[2], addr_3567_6, addr_positional[57083:57080], addr_14270_7);

wire[31:0] addr_14271_7;

Selector_2 s14271_7(wires_3567_6[3], addr_3567_6, addr_positional[57087:57084], addr_14271_7);

wire[31:0] addr_14272_7;

Selector_2 s14272_7(wires_3568_6[0], addr_3568_6, addr_positional[57091:57088], addr_14272_7);

wire[31:0] addr_14273_7;

Selector_2 s14273_7(wires_3568_6[1], addr_3568_6, addr_positional[57095:57092], addr_14273_7);

wire[31:0] addr_14274_7;

Selector_2 s14274_7(wires_3568_6[2], addr_3568_6, addr_positional[57099:57096], addr_14274_7);

wire[31:0] addr_14275_7;

Selector_2 s14275_7(wires_3568_6[3], addr_3568_6, addr_positional[57103:57100], addr_14275_7);

wire[31:0] addr_14276_7;

Selector_2 s14276_7(wires_3569_6[0], addr_3569_6, addr_positional[57107:57104], addr_14276_7);

wire[31:0] addr_14277_7;

Selector_2 s14277_7(wires_3569_6[1], addr_3569_6, addr_positional[57111:57108], addr_14277_7);

wire[31:0] addr_14278_7;

Selector_2 s14278_7(wires_3569_6[2], addr_3569_6, addr_positional[57115:57112], addr_14278_7);

wire[31:0] addr_14279_7;

Selector_2 s14279_7(wires_3569_6[3], addr_3569_6, addr_positional[57119:57116], addr_14279_7);

wire[31:0] addr_14280_7;

Selector_2 s14280_7(wires_3570_6[0], addr_3570_6, addr_positional[57123:57120], addr_14280_7);

wire[31:0] addr_14281_7;

Selector_2 s14281_7(wires_3570_6[1], addr_3570_6, addr_positional[57127:57124], addr_14281_7);

wire[31:0] addr_14282_7;

Selector_2 s14282_7(wires_3570_6[2], addr_3570_6, addr_positional[57131:57128], addr_14282_7);

wire[31:0] addr_14283_7;

Selector_2 s14283_7(wires_3570_6[3], addr_3570_6, addr_positional[57135:57132], addr_14283_7);

wire[31:0] addr_14284_7;

Selector_2 s14284_7(wires_3571_6[0], addr_3571_6, addr_positional[57139:57136], addr_14284_7);

wire[31:0] addr_14285_7;

Selector_2 s14285_7(wires_3571_6[1], addr_3571_6, addr_positional[57143:57140], addr_14285_7);

wire[31:0] addr_14286_7;

Selector_2 s14286_7(wires_3571_6[2], addr_3571_6, addr_positional[57147:57144], addr_14286_7);

wire[31:0] addr_14287_7;

Selector_2 s14287_7(wires_3571_6[3], addr_3571_6, addr_positional[57151:57148], addr_14287_7);

wire[31:0] addr_14288_7;

Selector_2 s14288_7(wires_3572_6[0], addr_3572_6, addr_positional[57155:57152], addr_14288_7);

wire[31:0] addr_14289_7;

Selector_2 s14289_7(wires_3572_6[1], addr_3572_6, addr_positional[57159:57156], addr_14289_7);

wire[31:0] addr_14290_7;

Selector_2 s14290_7(wires_3572_6[2], addr_3572_6, addr_positional[57163:57160], addr_14290_7);

wire[31:0] addr_14291_7;

Selector_2 s14291_7(wires_3572_6[3], addr_3572_6, addr_positional[57167:57164], addr_14291_7);

wire[31:0] addr_14292_7;

Selector_2 s14292_7(wires_3573_6[0], addr_3573_6, addr_positional[57171:57168], addr_14292_7);

wire[31:0] addr_14293_7;

Selector_2 s14293_7(wires_3573_6[1], addr_3573_6, addr_positional[57175:57172], addr_14293_7);

wire[31:0] addr_14294_7;

Selector_2 s14294_7(wires_3573_6[2], addr_3573_6, addr_positional[57179:57176], addr_14294_7);

wire[31:0] addr_14295_7;

Selector_2 s14295_7(wires_3573_6[3], addr_3573_6, addr_positional[57183:57180], addr_14295_7);

wire[31:0] addr_14296_7;

Selector_2 s14296_7(wires_3574_6[0], addr_3574_6, addr_positional[57187:57184], addr_14296_7);

wire[31:0] addr_14297_7;

Selector_2 s14297_7(wires_3574_6[1], addr_3574_6, addr_positional[57191:57188], addr_14297_7);

wire[31:0] addr_14298_7;

Selector_2 s14298_7(wires_3574_6[2], addr_3574_6, addr_positional[57195:57192], addr_14298_7);

wire[31:0] addr_14299_7;

Selector_2 s14299_7(wires_3574_6[3], addr_3574_6, addr_positional[57199:57196], addr_14299_7);

wire[31:0] addr_14300_7;

Selector_2 s14300_7(wires_3575_6[0], addr_3575_6, addr_positional[57203:57200], addr_14300_7);

wire[31:0] addr_14301_7;

Selector_2 s14301_7(wires_3575_6[1], addr_3575_6, addr_positional[57207:57204], addr_14301_7);

wire[31:0] addr_14302_7;

Selector_2 s14302_7(wires_3575_6[2], addr_3575_6, addr_positional[57211:57208], addr_14302_7);

wire[31:0] addr_14303_7;

Selector_2 s14303_7(wires_3575_6[3], addr_3575_6, addr_positional[57215:57212], addr_14303_7);

wire[31:0] addr_14304_7;

Selector_2 s14304_7(wires_3576_6[0], addr_3576_6, addr_positional[57219:57216], addr_14304_7);

wire[31:0] addr_14305_7;

Selector_2 s14305_7(wires_3576_6[1], addr_3576_6, addr_positional[57223:57220], addr_14305_7);

wire[31:0] addr_14306_7;

Selector_2 s14306_7(wires_3576_6[2], addr_3576_6, addr_positional[57227:57224], addr_14306_7);

wire[31:0] addr_14307_7;

Selector_2 s14307_7(wires_3576_6[3], addr_3576_6, addr_positional[57231:57228], addr_14307_7);

wire[31:0] addr_14308_7;

Selector_2 s14308_7(wires_3577_6[0], addr_3577_6, addr_positional[57235:57232], addr_14308_7);

wire[31:0] addr_14309_7;

Selector_2 s14309_7(wires_3577_6[1], addr_3577_6, addr_positional[57239:57236], addr_14309_7);

wire[31:0] addr_14310_7;

Selector_2 s14310_7(wires_3577_6[2], addr_3577_6, addr_positional[57243:57240], addr_14310_7);

wire[31:0] addr_14311_7;

Selector_2 s14311_7(wires_3577_6[3], addr_3577_6, addr_positional[57247:57244], addr_14311_7);

wire[31:0] addr_14312_7;

Selector_2 s14312_7(wires_3578_6[0], addr_3578_6, addr_positional[57251:57248], addr_14312_7);

wire[31:0] addr_14313_7;

Selector_2 s14313_7(wires_3578_6[1], addr_3578_6, addr_positional[57255:57252], addr_14313_7);

wire[31:0] addr_14314_7;

Selector_2 s14314_7(wires_3578_6[2], addr_3578_6, addr_positional[57259:57256], addr_14314_7);

wire[31:0] addr_14315_7;

Selector_2 s14315_7(wires_3578_6[3], addr_3578_6, addr_positional[57263:57260], addr_14315_7);

wire[31:0] addr_14316_7;

Selector_2 s14316_7(wires_3579_6[0], addr_3579_6, addr_positional[57267:57264], addr_14316_7);

wire[31:0] addr_14317_7;

Selector_2 s14317_7(wires_3579_6[1], addr_3579_6, addr_positional[57271:57268], addr_14317_7);

wire[31:0] addr_14318_7;

Selector_2 s14318_7(wires_3579_6[2], addr_3579_6, addr_positional[57275:57272], addr_14318_7);

wire[31:0] addr_14319_7;

Selector_2 s14319_7(wires_3579_6[3], addr_3579_6, addr_positional[57279:57276], addr_14319_7);

wire[31:0] addr_14320_7;

Selector_2 s14320_7(wires_3580_6[0], addr_3580_6, addr_positional[57283:57280], addr_14320_7);

wire[31:0] addr_14321_7;

Selector_2 s14321_7(wires_3580_6[1], addr_3580_6, addr_positional[57287:57284], addr_14321_7);

wire[31:0] addr_14322_7;

Selector_2 s14322_7(wires_3580_6[2], addr_3580_6, addr_positional[57291:57288], addr_14322_7);

wire[31:0] addr_14323_7;

Selector_2 s14323_7(wires_3580_6[3], addr_3580_6, addr_positional[57295:57292], addr_14323_7);

wire[31:0] addr_14324_7;

Selector_2 s14324_7(wires_3581_6[0], addr_3581_6, addr_positional[57299:57296], addr_14324_7);

wire[31:0] addr_14325_7;

Selector_2 s14325_7(wires_3581_6[1], addr_3581_6, addr_positional[57303:57300], addr_14325_7);

wire[31:0] addr_14326_7;

Selector_2 s14326_7(wires_3581_6[2], addr_3581_6, addr_positional[57307:57304], addr_14326_7);

wire[31:0] addr_14327_7;

Selector_2 s14327_7(wires_3581_6[3], addr_3581_6, addr_positional[57311:57308], addr_14327_7);

wire[31:0] addr_14328_7;

Selector_2 s14328_7(wires_3582_6[0], addr_3582_6, addr_positional[57315:57312], addr_14328_7);

wire[31:0] addr_14329_7;

Selector_2 s14329_7(wires_3582_6[1], addr_3582_6, addr_positional[57319:57316], addr_14329_7);

wire[31:0] addr_14330_7;

Selector_2 s14330_7(wires_3582_6[2], addr_3582_6, addr_positional[57323:57320], addr_14330_7);

wire[31:0] addr_14331_7;

Selector_2 s14331_7(wires_3582_6[3], addr_3582_6, addr_positional[57327:57324], addr_14331_7);

wire[31:0] addr_14332_7;

Selector_2 s14332_7(wires_3583_6[0], addr_3583_6, addr_positional[57331:57328], addr_14332_7);

wire[31:0] addr_14333_7;

Selector_2 s14333_7(wires_3583_6[1], addr_3583_6, addr_positional[57335:57332], addr_14333_7);

wire[31:0] addr_14334_7;

Selector_2 s14334_7(wires_3583_6[2], addr_3583_6, addr_positional[57339:57336], addr_14334_7);

wire[31:0] addr_14335_7;

Selector_2 s14335_7(wires_3583_6[3], addr_3583_6, addr_positional[57343:57340], addr_14335_7);

wire[31:0] addr_14336_7;

Selector_2 s14336_7(wires_3584_6[0], addr_3584_6, addr_positional[57347:57344], addr_14336_7);

wire[31:0] addr_14337_7;

Selector_2 s14337_7(wires_3584_6[1], addr_3584_6, addr_positional[57351:57348], addr_14337_7);

wire[31:0] addr_14338_7;

Selector_2 s14338_7(wires_3584_6[2], addr_3584_6, addr_positional[57355:57352], addr_14338_7);

wire[31:0] addr_14339_7;

Selector_2 s14339_7(wires_3584_6[3], addr_3584_6, addr_positional[57359:57356], addr_14339_7);

wire[31:0] addr_14340_7;

Selector_2 s14340_7(wires_3585_6[0], addr_3585_6, addr_positional[57363:57360], addr_14340_7);

wire[31:0] addr_14341_7;

Selector_2 s14341_7(wires_3585_6[1], addr_3585_6, addr_positional[57367:57364], addr_14341_7);

wire[31:0] addr_14342_7;

Selector_2 s14342_7(wires_3585_6[2], addr_3585_6, addr_positional[57371:57368], addr_14342_7);

wire[31:0] addr_14343_7;

Selector_2 s14343_7(wires_3585_6[3], addr_3585_6, addr_positional[57375:57372], addr_14343_7);

wire[31:0] addr_14344_7;

Selector_2 s14344_7(wires_3586_6[0], addr_3586_6, addr_positional[57379:57376], addr_14344_7);

wire[31:0] addr_14345_7;

Selector_2 s14345_7(wires_3586_6[1], addr_3586_6, addr_positional[57383:57380], addr_14345_7);

wire[31:0] addr_14346_7;

Selector_2 s14346_7(wires_3586_6[2], addr_3586_6, addr_positional[57387:57384], addr_14346_7);

wire[31:0] addr_14347_7;

Selector_2 s14347_7(wires_3586_6[3], addr_3586_6, addr_positional[57391:57388], addr_14347_7);

wire[31:0] addr_14348_7;

Selector_2 s14348_7(wires_3587_6[0], addr_3587_6, addr_positional[57395:57392], addr_14348_7);

wire[31:0] addr_14349_7;

Selector_2 s14349_7(wires_3587_6[1], addr_3587_6, addr_positional[57399:57396], addr_14349_7);

wire[31:0] addr_14350_7;

Selector_2 s14350_7(wires_3587_6[2], addr_3587_6, addr_positional[57403:57400], addr_14350_7);

wire[31:0] addr_14351_7;

Selector_2 s14351_7(wires_3587_6[3], addr_3587_6, addr_positional[57407:57404], addr_14351_7);

wire[31:0] addr_14352_7;

Selector_2 s14352_7(wires_3588_6[0], addr_3588_6, addr_positional[57411:57408], addr_14352_7);

wire[31:0] addr_14353_7;

Selector_2 s14353_7(wires_3588_6[1], addr_3588_6, addr_positional[57415:57412], addr_14353_7);

wire[31:0] addr_14354_7;

Selector_2 s14354_7(wires_3588_6[2], addr_3588_6, addr_positional[57419:57416], addr_14354_7);

wire[31:0] addr_14355_7;

Selector_2 s14355_7(wires_3588_6[3], addr_3588_6, addr_positional[57423:57420], addr_14355_7);

wire[31:0] addr_14356_7;

Selector_2 s14356_7(wires_3589_6[0], addr_3589_6, addr_positional[57427:57424], addr_14356_7);

wire[31:0] addr_14357_7;

Selector_2 s14357_7(wires_3589_6[1], addr_3589_6, addr_positional[57431:57428], addr_14357_7);

wire[31:0] addr_14358_7;

Selector_2 s14358_7(wires_3589_6[2], addr_3589_6, addr_positional[57435:57432], addr_14358_7);

wire[31:0] addr_14359_7;

Selector_2 s14359_7(wires_3589_6[3], addr_3589_6, addr_positional[57439:57436], addr_14359_7);

wire[31:0] addr_14360_7;

Selector_2 s14360_7(wires_3590_6[0], addr_3590_6, addr_positional[57443:57440], addr_14360_7);

wire[31:0] addr_14361_7;

Selector_2 s14361_7(wires_3590_6[1], addr_3590_6, addr_positional[57447:57444], addr_14361_7);

wire[31:0] addr_14362_7;

Selector_2 s14362_7(wires_3590_6[2], addr_3590_6, addr_positional[57451:57448], addr_14362_7);

wire[31:0] addr_14363_7;

Selector_2 s14363_7(wires_3590_6[3], addr_3590_6, addr_positional[57455:57452], addr_14363_7);

wire[31:0] addr_14364_7;

Selector_2 s14364_7(wires_3591_6[0], addr_3591_6, addr_positional[57459:57456], addr_14364_7);

wire[31:0] addr_14365_7;

Selector_2 s14365_7(wires_3591_6[1], addr_3591_6, addr_positional[57463:57460], addr_14365_7);

wire[31:0] addr_14366_7;

Selector_2 s14366_7(wires_3591_6[2], addr_3591_6, addr_positional[57467:57464], addr_14366_7);

wire[31:0] addr_14367_7;

Selector_2 s14367_7(wires_3591_6[3], addr_3591_6, addr_positional[57471:57468], addr_14367_7);

wire[31:0] addr_14368_7;

Selector_2 s14368_7(wires_3592_6[0], addr_3592_6, addr_positional[57475:57472], addr_14368_7);

wire[31:0] addr_14369_7;

Selector_2 s14369_7(wires_3592_6[1], addr_3592_6, addr_positional[57479:57476], addr_14369_7);

wire[31:0] addr_14370_7;

Selector_2 s14370_7(wires_3592_6[2], addr_3592_6, addr_positional[57483:57480], addr_14370_7);

wire[31:0] addr_14371_7;

Selector_2 s14371_7(wires_3592_6[3], addr_3592_6, addr_positional[57487:57484], addr_14371_7);

wire[31:0] addr_14372_7;

Selector_2 s14372_7(wires_3593_6[0], addr_3593_6, addr_positional[57491:57488], addr_14372_7);

wire[31:0] addr_14373_7;

Selector_2 s14373_7(wires_3593_6[1], addr_3593_6, addr_positional[57495:57492], addr_14373_7);

wire[31:0] addr_14374_7;

Selector_2 s14374_7(wires_3593_6[2], addr_3593_6, addr_positional[57499:57496], addr_14374_7);

wire[31:0] addr_14375_7;

Selector_2 s14375_7(wires_3593_6[3], addr_3593_6, addr_positional[57503:57500], addr_14375_7);

wire[31:0] addr_14376_7;

Selector_2 s14376_7(wires_3594_6[0], addr_3594_6, addr_positional[57507:57504], addr_14376_7);

wire[31:0] addr_14377_7;

Selector_2 s14377_7(wires_3594_6[1], addr_3594_6, addr_positional[57511:57508], addr_14377_7);

wire[31:0] addr_14378_7;

Selector_2 s14378_7(wires_3594_6[2], addr_3594_6, addr_positional[57515:57512], addr_14378_7);

wire[31:0] addr_14379_7;

Selector_2 s14379_7(wires_3594_6[3], addr_3594_6, addr_positional[57519:57516], addr_14379_7);

wire[31:0] addr_14380_7;

Selector_2 s14380_7(wires_3595_6[0], addr_3595_6, addr_positional[57523:57520], addr_14380_7);

wire[31:0] addr_14381_7;

Selector_2 s14381_7(wires_3595_6[1], addr_3595_6, addr_positional[57527:57524], addr_14381_7);

wire[31:0] addr_14382_7;

Selector_2 s14382_7(wires_3595_6[2], addr_3595_6, addr_positional[57531:57528], addr_14382_7);

wire[31:0] addr_14383_7;

Selector_2 s14383_7(wires_3595_6[3], addr_3595_6, addr_positional[57535:57532], addr_14383_7);

wire[31:0] addr_14384_7;

Selector_2 s14384_7(wires_3596_6[0], addr_3596_6, addr_positional[57539:57536], addr_14384_7);

wire[31:0] addr_14385_7;

Selector_2 s14385_7(wires_3596_6[1], addr_3596_6, addr_positional[57543:57540], addr_14385_7);

wire[31:0] addr_14386_7;

Selector_2 s14386_7(wires_3596_6[2], addr_3596_6, addr_positional[57547:57544], addr_14386_7);

wire[31:0] addr_14387_7;

Selector_2 s14387_7(wires_3596_6[3], addr_3596_6, addr_positional[57551:57548], addr_14387_7);

wire[31:0] addr_14388_7;

Selector_2 s14388_7(wires_3597_6[0], addr_3597_6, addr_positional[57555:57552], addr_14388_7);

wire[31:0] addr_14389_7;

Selector_2 s14389_7(wires_3597_6[1], addr_3597_6, addr_positional[57559:57556], addr_14389_7);

wire[31:0] addr_14390_7;

Selector_2 s14390_7(wires_3597_6[2], addr_3597_6, addr_positional[57563:57560], addr_14390_7);

wire[31:0] addr_14391_7;

Selector_2 s14391_7(wires_3597_6[3], addr_3597_6, addr_positional[57567:57564], addr_14391_7);

wire[31:0] addr_14392_7;

Selector_2 s14392_7(wires_3598_6[0], addr_3598_6, addr_positional[57571:57568], addr_14392_7);

wire[31:0] addr_14393_7;

Selector_2 s14393_7(wires_3598_6[1], addr_3598_6, addr_positional[57575:57572], addr_14393_7);

wire[31:0] addr_14394_7;

Selector_2 s14394_7(wires_3598_6[2], addr_3598_6, addr_positional[57579:57576], addr_14394_7);

wire[31:0] addr_14395_7;

Selector_2 s14395_7(wires_3598_6[3], addr_3598_6, addr_positional[57583:57580], addr_14395_7);

wire[31:0] addr_14396_7;

Selector_2 s14396_7(wires_3599_6[0], addr_3599_6, addr_positional[57587:57584], addr_14396_7);

wire[31:0] addr_14397_7;

Selector_2 s14397_7(wires_3599_6[1], addr_3599_6, addr_positional[57591:57588], addr_14397_7);

wire[31:0] addr_14398_7;

Selector_2 s14398_7(wires_3599_6[2], addr_3599_6, addr_positional[57595:57592], addr_14398_7);

wire[31:0] addr_14399_7;

Selector_2 s14399_7(wires_3599_6[3], addr_3599_6, addr_positional[57599:57596], addr_14399_7);

wire[31:0] addr_14400_7;

Selector_2 s14400_7(wires_3600_6[0], addr_3600_6, addr_positional[57603:57600], addr_14400_7);

wire[31:0] addr_14401_7;

Selector_2 s14401_7(wires_3600_6[1], addr_3600_6, addr_positional[57607:57604], addr_14401_7);

wire[31:0] addr_14402_7;

Selector_2 s14402_7(wires_3600_6[2], addr_3600_6, addr_positional[57611:57608], addr_14402_7);

wire[31:0] addr_14403_7;

Selector_2 s14403_7(wires_3600_6[3], addr_3600_6, addr_positional[57615:57612], addr_14403_7);

wire[31:0] addr_14404_7;

Selector_2 s14404_7(wires_3601_6[0], addr_3601_6, addr_positional[57619:57616], addr_14404_7);

wire[31:0] addr_14405_7;

Selector_2 s14405_7(wires_3601_6[1], addr_3601_6, addr_positional[57623:57620], addr_14405_7);

wire[31:0] addr_14406_7;

Selector_2 s14406_7(wires_3601_6[2], addr_3601_6, addr_positional[57627:57624], addr_14406_7);

wire[31:0] addr_14407_7;

Selector_2 s14407_7(wires_3601_6[3], addr_3601_6, addr_positional[57631:57628], addr_14407_7);

wire[31:0] addr_14408_7;

Selector_2 s14408_7(wires_3602_6[0], addr_3602_6, addr_positional[57635:57632], addr_14408_7);

wire[31:0] addr_14409_7;

Selector_2 s14409_7(wires_3602_6[1], addr_3602_6, addr_positional[57639:57636], addr_14409_7);

wire[31:0] addr_14410_7;

Selector_2 s14410_7(wires_3602_6[2], addr_3602_6, addr_positional[57643:57640], addr_14410_7);

wire[31:0] addr_14411_7;

Selector_2 s14411_7(wires_3602_6[3], addr_3602_6, addr_positional[57647:57644], addr_14411_7);

wire[31:0] addr_14412_7;

Selector_2 s14412_7(wires_3603_6[0], addr_3603_6, addr_positional[57651:57648], addr_14412_7);

wire[31:0] addr_14413_7;

Selector_2 s14413_7(wires_3603_6[1], addr_3603_6, addr_positional[57655:57652], addr_14413_7);

wire[31:0] addr_14414_7;

Selector_2 s14414_7(wires_3603_6[2], addr_3603_6, addr_positional[57659:57656], addr_14414_7);

wire[31:0] addr_14415_7;

Selector_2 s14415_7(wires_3603_6[3], addr_3603_6, addr_positional[57663:57660], addr_14415_7);

wire[31:0] addr_14416_7;

Selector_2 s14416_7(wires_3604_6[0], addr_3604_6, addr_positional[57667:57664], addr_14416_7);

wire[31:0] addr_14417_7;

Selector_2 s14417_7(wires_3604_6[1], addr_3604_6, addr_positional[57671:57668], addr_14417_7);

wire[31:0] addr_14418_7;

Selector_2 s14418_7(wires_3604_6[2], addr_3604_6, addr_positional[57675:57672], addr_14418_7);

wire[31:0] addr_14419_7;

Selector_2 s14419_7(wires_3604_6[3], addr_3604_6, addr_positional[57679:57676], addr_14419_7);

wire[31:0] addr_14420_7;

Selector_2 s14420_7(wires_3605_6[0], addr_3605_6, addr_positional[57683:57680], addr_14420_7);

wire[31:0] addr_14421_7;

Selector_2 s14421_7(wires_3605_6[1], addr_3605_6, addr_positional[57687:57684], addr_14421_7);

wire[31:0] addr_14422_7;

Selector_2 s14422_7(wires_3605_6[2], addr_3605_6, addr_positional[57691:57688], addr_14422_7);

wire[31:0] addr_14423_7;

Selector_2 s14423_7(wires_3605_6[3], addr_3605_6, addr_positional[57695:57692], addr_14423_7);

wire[31:0] addr_14424_7;

Selector_2 s14424_7(wires_3606_6[0], addr_3606_6, addr_positional[57699:57696], addr_14424_7);

wire[31:0] addr_14425_7;

Selector_2 s14425_7(wires_3606_6[1], addr_3606_6, addr_positional[57703:57700], addr_14425_7);

wire[31:0] addr_14426_7;

Selector_2 s14426_7(wires_3606_6[2], addr_3606_6, addr_positional[57707:57704], addr_14426_7);

wire[31:0] addr_14427_7;

Selector_2 s14427_7(wires_3606_6[3], addr_3606_6, addr_positional[57711:57708], addr_14427_7);

wire[31:0] addr_14428_7;

Selector_2 s14428_7(wires_3607_6[0], addr_3607_6, addr_positional[57715:57712], addr_14428_7);

wire[31:0] addr_14429_7;

Selector_2 s14429_7(wires_3607_6[1], addr_3607_6, addr_positional[57719:57716], addr_14429_7);

wire[31:0] addr_14430_7;

Selector_2 s14430_7(wires_3607_6[2], addr_3607_6, addr_positional[57723:57720], addr_14430_7);

wire[31:0] addr_14431_7;

Selector_2 s14431_7(wires_3607_6[3], addr_3607_6, addr_positional[57727:57724], addr_14431_7);

wire[31:0] addr_14432_7;

Selector_2 s14432_7(wires_3608_6[0], addr_3608_6, addr_positional[57731:57728], addr_14432_7);

wire[31:0] addr_14433_7;

Selector_2 s14433_7(wires_3608_6[1], addr_3608_6, addr_positional[57735:57732], addr_14433_7);

wire[31:0] addr_14434_7;

Selector_2 s14434_7(wires_3608_6[2], addr_3608_6, addr_positional[57739:57736], addr_14434_7);

wire[31:0] addr_14435_7;

Selector_2 s14435_7(wires_3608_6[3], addr_3608_6, addr_positional[57743:57740], addr_14435_7);

wire[31:0] addr_14436_7;

Selector_2 s14436_7(wires_3609_6[0], addr_3609_6, addr_positional[57747:57744], addr_14436_7);

wire[31:0] addr_14437_7;

Selector_2 s14437_7(wires_3609_6[1], addr_3609_6, addr_positional[57751:57748], addr_14437_7);

wire[31:0] addr_14438_7;

Selector_2 s14438_7(wires_3609_6[2], addr_3609_6, addr_positional[57755:57752], addr_14438_7);

wire[31:0] addr_14439_7;

Selector_2 s14439_7(wires_3609_6[3], addr_3609_6, addr_positional[57759:57756], addr_14439_7);

wire[31:0] addr_14440_7;

Selector_2 s14440_7(wires_3610_6[0], addr_3610_6, addr_positional[57763:57760], addr_14440_7);

wire[31:0] addr_14441_7;

Selector_2 s14441_7(wires_3610_6[1], addr_3610_6, addr_positional[57767:57764], addr_14441_7);

wire[31:0] addr_14442_7;

Selector_2 s14442_7(wires_3610_6[2], addr_3610_6, addr_positional[57771:57768], addr_14442_7);

wire[31:0] addr_14443_7;

Selector_2 s14443_7(wires_3610_6[3], addr_3610_6, addr_positional[57775:57772], addr_14443_7);

wire[31:0] addr_14444_7;

Selector_2 s14444_7(wires_3611_6[0], addr_3611_6, addr_positional[57779:57776], addr_14444_7);

wire[31:0] addr_14445_7;

Selector_2 s14445_7(wires_3611_6[1], addr_3611_6, addr_positional[57783:57780], addr_14445_7);

wire[31:0] addr_14446_7;

Selector_2 s14446_7(wires_3611_6[2], addr_3611_6, addr_positional[57787:57784], addr_14446_7);

wire[31:0] addr_14447_7;

Selector_2 s14447_7(wires_3611_6[3], addr_3611_6, addr_positional[57791:57788], addr_14447_7);

wire[31:0] addr_14448_7;

Selector_2 s14448_7(wires_3612_6[0], addr_3612_6, addr_positional[57795:57792], addr_14448_7);

wire[31:0] addr_14449_7;

Selector_2 s14449_7(wires_3612_6[1], addr_3612_6, addr_positional[57799:57796], addr_14449_7);

wire[31:0] addr_14450_7;

Selector_2 s14450_7(wires_3612_6[2], addr_3612_6, addr_positional[57803:57800], addr_14450_7);

wire[31:0] addr_14451_7;

Selector_2 s14451_7(wires_3612_6[3], addr_3612_6, addr_positional[57807:57804], addr_14451_7);

wire[31:0] addr_14452_7;

Selector_2 s14452_7(wires_3613_6[0], addr_3613_6, addr_positional[57811:57808], addr_14452_7);

wire[31:0] addr_14453_7;

Selector_2 s14453_7(wires_3613_6[1], addr_3613_6, addr_positional[57815:57812], addr_14453_7);

wire[31:0] addr_14454_7;

Selector_2 s14454_7(wires_3613_6[2], addr_3613_6, addr_positional[57819:57816], addr_14454_7);

wire[31:0] addr_14455_7;

Selector_2 s14455_7(wires_3613_6[3], addr_3613_6, addr_positional[57823:57820], addr_14455_7);

wire[31:0] addr_14456_7;

Selector_2 s14456_7(wires_3614_6[0], addr_3614_6, addr_positional[57827:57824], addr_14456_7);

wire[31:0] addr_14457_7;

Selector_2 s14457_7(wires_3614_6[1], addr_3614_6, addr_positional[57831:57828], addr_14457_7);

wire[31:0] addr_14458_7;

Selector_2 s14458_7(wires_3614_6[2], addr_3614_6, addr_positional[57835:57832], addr_14458_7);

wire[31:0] addr_14459_7;

Selector_2 s14459_7(wires_3614_6[3], addr_3614_6, addr_positional[57839:57836], addr_14459_7);

wire[31:0] addr_14460_7;

Selector_2 s14460_7(wires_3615_6[0], addr_3615_6, addr_positional[57843:57840], addr_14460_7);

wire[31:0] addr_14461_7;

Selector_2 s14461_7(wires_3615_6[1], addr_3615_6, addr_positional[57847:57844], addr_14461_7);

wire[31:0] addr_14462_7;

Selector_2 s14462_7(wires_3615_6[2], addr_3615_6, addr_positional[57851:57848], addr_14462_7);

wire[31:0] addr_14463_7;

Selector_2 s14463_7(wires_3615_6[3], addr_3615_6, addr_positional[57855:57852], addr_14463_7);

wire[31:0] addr_14464_7;

Selector_2 s14464_7(wires_3616_6[0], addr_3616_6, addr_positional[57859:57856], addr_14464_7);

wire[31:0] addr_14465_7;

Selector_2 s14465_7(wires_3616_6[1], addr_3616_6, addr_positional[57863:57860], addr_14465_7);

wire[31:0] addr_14466_7;

Selector_2 s14466_7(wires_3616_6[2], addr_3616_6, addr_positional[57867:57864], addr_14466_7);

wire[31:0] addr_14467_7;

Selector_2 s14467_7(wires_3616_6[3], addr_3616_6, addr_positional[57871:57868], addr_14467_7);

wire[31:0] addr_14468_7;

Selector_2 s14468_7(wires_3617_6[0], addr_3617_6, addr_positional[57875:57872], addr_14468_7);

wire[31:0] addr_14469_7;

Selector_2 s14469_7(wires_3617_6[1], addr_3617_6, addr_positional[57879:57876], addr_14469_7);

wire[31:0] addr_14470_7;

Selector_2 s14470_7(wires_3617_6[2], addr_3617_6, addr_positional[57883:57880], addr_14470_7);

wire[31:0] addr_14471_7;

Selector_2 s14471_7(wires_3617_6[3], addr_3617_6, addr_positional[57887:57884], addr_14471_7);

wire[31:0] addr_14472_7;

Selector_2 s14472_7(wires_3618_6[0], addr_3618_6, addr_positional[57891:57888], addr_14472_7);

wire[31:0] addr_14473_7;

Selector_2 s14473_7(wires_3618_6[1], addr_3618_6, addr_positional[57895:57892], addr_14473_7);

wire[31:0] addr_14474_7;

Selector_2 s14474_7(wires_3618_6[2], addr_3618_6, addr_positional[57899:57896], addr_14474_7);

wire[31:0] addr_14475_7;

Selector_2 s14475_7(wires_3618_6[3], addr_3618_6, addr_positional[57903:57900], addr_14475_7);

wire[31:0] addr_14476_7;

Selector_2 s14476_7(wires_3619_6[0], addr_3619_6, addr_positional[57907:57904], addr_14476_7);

wire[31:0] addr_14477_7;

Selector_2 s14477_7(wires_3619_6[1], addr_3619_6, addr_positional[57911:57908], addr_14477_7);

wire[31:0] addr_14478_7;

Selector_2 s14478_7(wires_3619_6[2], addr_3619_6, addr_positional[57915:57912], addr_14478_7);

wire[31:0] addr_14479_7;

Selector_2 s14479_7(wires_3619_6[3], addr_3619_6, addr_positional[57919:57916], addr_14479_7);

wire[31:0] addr_14480_7;

Selector_2 s14480_7(wires_3620_6[0], addr_3620_6, addr_positional[57923:57920], addr_14480_7);

wire[31:0] addr_14481_7;

Selector_2 s14481_7(wires_3620_6[1], addr_3620_6, addr_positional[57927:57924], addr_14481_7);

wire[31:0] addr_14482_7;

Selector_2 s14482_7(wires_3620_6[2], addr_3620_6, addr_positional[57931:57928], addr_14482_7);

wire[31:0] addr_14483_7;

Selector_2 s14483_7(wires_3620_6[3], addr_3620_6, addr_positional[57935:57932], addr_14483_7);

wire[31:0] addr_14484_7;

Selector_2 s14484_7(wires_3621_6[0], addr_3621_6, addr_positional[57939:57936], addr_14484_7);

wire[31:0] addr_14485_7;

Selector_2 s14485_7(wires_3621_6[1], addr_3621_6, addr_positional[57943:57940], addr_14485_7);

wire[31:0] addr_14486_7;

Selector_2 s14486_7(wires_3621_6[2], addr_3621_6, addr_positional[57947:57944], addr_14486_7);

wire[31:0] addr_14487_7;

Selector_2 s14487_7(wires_3621_6[3], addr_3621_6, addr_positional[57951:57948], addr_14487_7);

wire[31:0] addr_14488_7;

Selector_2 s14488_7(wires_3622_6[0], addr_3622_6, addr_positional[57955:57952], addr_14488_7);

wire[31:0] addr_14489_7;

Selector_2 s14489_7(wires_3622_6[1], addr_3622_6, addr_positional[57959:57956], addr_14489_7);

wire[31:0] addr_14490_7;

Selector_2 s14490_7(wires_3622_6[2], addr_3622_6, addr_positional[57963:57960], addr_14490_7);

wire[31:0] addr_14491_7;

Selector_2 s14491_7(wires_3622_6[3], addr_3622_6, addr_positional[57967:57964], addr_14491_7);

wire[31:0] addr_14492_7;

Selector_2 s14492_7(wires_3623_6[0], addr_3623_6, addr_positional[57971:57968], addr_14492_7);

wire[31:0] addr_14493_7;

Selector_2 s14493_7(wires_3623_6[1], addr_3623_6, addr_positional[57975:57972], addr_14493_7);

wire[31:0] addr_14494_7;

Selector_2 s14494_7(wires_3623_6[2], addr_3623_6, addr_positional[57979:57976], addr_14494_7);

wire[31:0] addr_14495_7;

Selector_2 s14495_7(wires_3623_6[3], addr_3623_6, addr_positional[57983:57980], addr_14495_7);

wire[31:0] addr_14496_7;

Selector_2 s14496_7(wires_3624_6[0], addr_3624_6, addr_positional[57987:57984], addr_14496_7);

wire[31:0] addr_14497_7;

Selector_2 s14497_7(wires_3624_6[1], addr_3624_6, addr_positional[57991:57988], addr_14497_7);

wire[31:0] addr_14498_7;

Selector_2 s14498_7(wires_3624_6[2], addr_3624_6, addr_positional[57995:57992], addr_14498_7);

wire[31:0] addr_14499_7;

Selector_2 s14499_7(wires_3624_6[3], addr_3624_6, addr_positional[57999:57996], addr_14499_7);

wire[31:0] addr_14500_7;

Selector_2 s14500_7(wires_3625_6[0], addr_3625_6, addr_positional[58003:58000], addr_14500_7);

wire[31:0] addr_14501_7;

Selector_2 s14501_7(wires_3625_6[1], addr_3625_6, addr_positional[58007:58004], addr_14501_7);

wire[31:0] addr_14502_7;

Selector_2 s14502_7(wires_3625_6[2], addr_3625_6, addr_positional[58011:58008], addr_14502_7);

wire[31:0] addr_14503_7;

Selector_2 s14503_7(wires_3625_6[3], addr_3625_6, addr_positional[58015:58012], addr_14503_7);

wire[31:0] addr_14504_7;

Selector_2 s14504_7(wires_3626_6[0], addr_3626_6, addr_positional[58019:58016], addr_14504_7);

wire[31:0] addr_14505_7;

Selector_2 s14505_7(wires_3626_6[1], addr_3626_6, addr_positional[58023:58020], addr_14505_7);

wire[31:0] addr_14506_7;

Selector_2 s14506_7(wires_3626_6[2], addr_3626_6, addr_positional[58027:58024], addr_14506_7);

wire[31:0] addr_14507_7;

Selector_2 s14507_7(wires_3626_6[3], addr_3626_6, addr_positional[58031:58028], addr_14507_7);

wire[31:0] addr_14508_7;

Selector_2 s14508_7(wires_3627_6[0], addr_3627_6, addr_positional[58035:58032], addr_14508_7);

wire[31:0] addr_14509_7;

Selector_2 s14509_7(wires_3627_6[1], addr_3627_6, addr_positional[58039:58036], addr_14509_7);

wire[31:0] addr_14510_7;

Selector_2 s14510_7(wires_3627_6[2], addr_3627_6, addr_positional[58043:58040], addr_14510_7);

wire[31:0] addr_14511_7;

Selector_2 s14511_7(wires_3627_6[3], addr_3627_6, addr_positional[58047:58044], addr_14511_7);

wire[31:0] addr_14512_7;

Selector_2 s14512_7(wires_3628_6[0], addr_3628_6, addr_positional[58051:58048], addr_14512_7);

wire[31:0] addr_14513_7;

Selector_2 s14513_7(wires_3628_6[1], addr_3628_6, addr_positional[58055:58052], addr_14513_7);

wire[31:0] addr_14514_7;

Selector_2 s14514_7(wires_3628_6[2], addr_3628_6, addr_positional[58059:58056], addr_14514_7);

wire[31:0] addr_14515_7;

Selector_2 s14515_7(wires_3628_6[3], addr_3628_6, addr_positional[58063:58060], addr_14515_7);

wire[31:0] addr_14516_7;

Selector_2 s14516_7(wires_3629_6[0], addr_3629_6, addr_positional[58067:58064], addr_14516_7);

wire[31:0] addr_14517_7;

Selector_2 s14517_7(wires_3629_6[1], addr_3629_6, addr_positional[58071:58068], addr_14517_7);

wire[31:0] addr_14518_7;

Selector_2 s14518_7(wires_3629_6[2], addr_3629_6, addr_positional[58075:58072], addr_14518_7);

wire[31:0] addr_14519_7;

Selector_2 s14519_7(wires_3629_6[3], addr_3629_6, addr_positional[58079:58076], addr_14519_7);

wire[31:0] addr_14520_7;

Selector_2 s14520_7(wires_3630_6[0], addr_3630_6, addr_positional[58083:58080], addr_14520_7);

wire[31:0] addr_14521_7;

Selector_2 s14521_7(wires_3630_6[1], addr_3630_6, addr_positional[58087:58084], addr_14521_7);

wire[31:0] addr_14522_7;

Selector_2 s14522_7(wires_3630_6[2], addr_3630_6, addr_positional[58091:58088], addr_14522_7);

wire[31:0] addr_14523_7;

Selector_2 s14523_7(wires_3630_6[3], addr_3630_6, addr_positional[58095:58092], addr_14523_7);

wire[31:0] addr_14524_7;

Selector_2 s14524_7(wires_3631_6[0], addr_3631_6, addr_positional[58099:58096], addr_14524_7);

wire[31:0] addr_14525_7;

Selector_2 s14525_7(wires_3631_6[1], addr_3631_6, addr_positional[58103:58100], addr_14525_7);

wire[31:0] addr_14526_7;

Selector_2 s14526_7(wires_3631_6[2], addr_3631_6, addr_positional[58107:58104], addr_14526_7);

wire[31:0] addr_14527_7;

Selector_2 s14527_7(wires_3631_6[3], addr_3631_6, addr_positional[58111:58108], addr_14527_7);

wire[31:0] addr_14528_7;

Selector_2 s14528_7(wires_3632_6[0], addr_3632_6, addr_positional[58115:58112], addr_14528_7);

wire[31:0] addr_14529_7;

Selector_2 s14529_7(wires_3632_6[1], addr_3632_6, addr_positional[58119:58116], addr_14529_7);

wire[31:0] addr_14530_7;

Selector_2 s14530_7(wires_3632_6[2], addr_3632_6, addr_positional[58123:58120], addr_14530_7);

wire[31:0] addr_14531_7;

Selector_2 s14531_7(wires_3632_6[3], addr_3632_6, addr_positional[58127:58124], addr_14531_7);

wire[31:0] addr_14532_7;

Selector_2 s14532_7(wires_3633_6[0], addr_3633_6, addr_positional[58131:58128], addr_14532_7);

wire[31:0] addr_14533_7;

Selector_2 s14533_7(wires_3633_6[1], addr_3633_6, addr_positional[58135:58132], addr_14533_7);

wire[31:0] addr_14534_7;

Selector_2 s14534_7(wires_3633_6[2], addr_3633_6, addr_positional[58139:58136], addr_14534_7);

wire[31:0] addr_14535_7;

Selector_2 s14535_7(wires_3633_6[3], addr_3633_6, addr_positional[58143:58140], addr_14535_7);

wire[31:0] addr_14536_7;

Selector_2 s14536_7(wires_3634_6[0], addr_3634_6, addr_positional[58147:58144], addr_14536_7);

wire[31:0] addr_14537_7;

Selector_2 s14537_7(wires_3634_6[1], addr_3634_6, addr_positional[58151:58148], addr_14537_7);

wire[31:0] addr_14538_7;

Selector_2 s14538_7(wires_3634_6[2], addr_3634_6, addr_positional[58155:58152], addr_14538_7);

wire[31:0] addr_14539_7;

Selector_2 s14539_7(wires_3634_6[3], addr_3634_6, addr_positional[58159:58156], addr_14539_7);

wire[31:0] addr_14540_7;

Selector_2 s14540_7(wires_3635_6[0], addr_3635_6, addr_positional[58163:58160], addr_14540_7);

wire[31:0] addr_14541_7;

Selector_2 s14541_7(wires_3635_6[1], addr_3635_6, addr_positional[58167:58164], addr_14541_7);

wire[31:0] addr_14542_7;

Selector_2 s14542_7(wires_3635_6[2], addr_3635_6, addr_positional[58171:58168], addr_14542_7);

wire[31:0] addr_14543_7;

Selector_2 s14543_7(wires_3635_6[3], addr_3635_6, addr_positional[58175:58172], addr_14543_7);

wire[31:0] addr_14544_7;

Selector_2 s14544_7(wires_3636_6[0], addr_3636_6, addr_positional[58179:58176], addr_14544_7);

wire[31:0] addr_14545_7;

Selector_2 s14545_7(wires_3636_6[1], addr_3636_6, addr_positional[58183:58180], addr_14545_7);

wire[31:0] addr_14546_7;

Selector_2 s14546_7(wires_3636_6[2], addr_3636_6, addr_positional[58187:58184], addr_14546_7);

wire[31:0] addr_14547_7;

Selector_2 s14547_7(wires_3636_6[3], addr_3636_6, addr_positional[58191:58188], addr_14547_7);

wire[31:0] addr_14548_7;

Selector_2 s14548_7(wires_3637_6[0], addr_3637_6, addr_positional[58195:58192], addr_14548_7);

wire[31:0] addr_14549_7;

Selector_2 s14549_7(wires_3637_6[1], addr_3637_6, addr_positional[58199:58196], addr_14549_7);

wire[31:0] addr_14550_7;

Selector_2 s14550_7(wires_3637_6[2], addr_3637_6, addr_positional[58203:58200], addr_14550_7);

wire[31:0] addr_14551_7;

Selector_2 s14551_7(wires_3637_6[3], addr_3637_6, addr_positional[58207:58204], addr_14551_7);

wire[31:0] addr_14552_7;

Selector_2 s14552_7(wires_3638_6[0], addr_3638_6, addr_positional[58211:58208], addr_14552_7);

wire[31:0] addr_14553_7;

Selector_2 s14553_7(wires_3638_6[1], addr_3638_6, addr_positional[58215:58212], addr_14553_7);

wire[31:0] addr_14554_7;

Selector_2 s14554_7(wires_3638_6[2], addr_3638_6, addr_positional[58219:58216], addr_14554_7);

wire[31:0] addr_14555_7;

Selector_2 s14555_7(wires_3638_6[3], addr_3638_6, addr_positional[58223:58220], addr_14555_7);

wire[31:0] addr_14556_7;

Selector_2 s14556_7(wires_3639_6[0], addr_3639_6, addr_positional[58227:58224], addr_14556_7);

wire[31:0] addr_14557_7;

Selector_2 s14557_7(wires_3639_6[1], addr_3639_6, addr_positional[58231:58228], addr_14557_7);

wire[31:0] addr_14558_7;

Selector_2 s14558_7(wires_3639_6[2], addr_3639_6, addr_positional[58235:58232], addr_14558_7);

wire[31:0] addr_14559_7;

Selector_2 s14559_7(wires_3639_6[3], addr_3639_6, addr_positional[58239:58236], addr_14559_7);

wire[31:0] addr_14560_7;

Selector_2 s14560_7(wires_3640_6[0], addr_3640_6, addr_positional[58243:58240], addr_14560_7);

wire[31:0] addr_14561_7;

Selector_2 s14561_7(wires_3640_6[1], addr_3640_6, addr_positional[58247:58244], addr_14561_7);

wire[31:0] addr_14562_7;

Selector_2 s14562_7(wires_3640_6[2], addr_3640_6, addr_positional[58251:58248], addr_14562_7);

wire[31:0] addr_14563_7;

Selector_2 s14563_7(wires_3640_6[3], addr_3640_6, addr_positional[58255:58252], addr_14563_7);

wire[31:0] addr_14564_7;

Selector_2 s14564_7(wires_3641_6[0], addr_3641_6, addr_positional[58259:58256], addr_14564_7);

wire[31:0] addr_14565_7;

Selector_2 s14565_7(wires_3641_6[1], addr_3641_6, addr_positional[58263:58260], addr_14565_7);

wire[31:0] addr_14566_7;

Selector_2 s14566_7(wires_3641_6[2], addr_3641_6, addr_positional[58267:58264], addr_14566_7);

wire[31:0] addr_14567_7;

Selector_2 s14567_7(wires_3641_6[3], addr_3641_6, addr_positional[58271:58268], addr_14567_7);

wire[31:0] addr_14568_7;

Selector_2 s14568_7(wires_3642_6[0], addr_3642_6, addr_positional[58275:58272], addr_14568_7);

wire[31:0] addr_14569_7;

Selector_2 s14569_7(wires_3642_6[1], addr_3642_6, addr_positional[58279:58276], addr_14569_7);

wire[31:0] addr_14570_7;

Selector_2 s14570_7(wires_3642_6[2], addr_3642_6, addr_positional[58283:58280], addr_14570_7);

wire[31:0] addr_14571_7;

Selector_2 s14571_7(wires_3642_6[3], addr_3642_6, addr_positional[58287:58284], addr_14571_7);

wire[31:0] addr_14572_7;

Selector_2 s14572_7(wires_3643_6[0], addr_3643_6, addr_positional[58291:58288], addr_14572_7);

wire[31:0] addr_14573_7;

Selector_2 s14573_7(wires_3643_6[1], addr_3643_6, addr_positional[58295:58292], addr_14573_7);

wire[31:0] addr_14574_7;

Selector_2 s14574_7(wires_3643_6[2], addr_3643_6, addr_positional[58299:58296], addr_14574_7);

wire[31:0] addr_14575_7;

Selector_2 s14575_7(wires_3643_6[3], addr_3643_6, addr_positional[58303:58300], addr_14575_7);

wire[31:0] addr_14576_7;

Selector_2 s14576_7(wires_3644_6[0], addr_3644_6, addr_positional[58307:58304], addr_14576_7);

wire[31:0] addr_14577_7;

Selector_2 s14577_7(wires_3644_6[1], addr_3644_6, addr_positional[58311:58308], addr_14577_7);

wire[31:0] addr_14578_7;

Selector_2 s14578_7(wires_3644_6[2], addr_3644_6, addr_positional[58315:58312], addr_14578_7);

wire[31:0] addr_14579_7;

Selector_2 s14579_7(wires_3644_6[3], addr_3644_6, addr_positional[58319:58316], addr_14579_7);

wire[31:0] addr_14580_7;

Selector_2 s14580_7(wires_3645_6[0], addr_3645_6, addr_positional[58323:58320], addr_14580_7);

wire[31:0] addr_14581_7;

Selector_2 s14581_7(wires_3645_6[1], addr_3645_6, addr_positional[58327:58324], addr_14581_7);

wire[31:0] addr_14582_7;

Selector_2 s14582_7(wires_3645_6[2], addr_3645_6, addr_positional[58331:58328], addr_14582_7);

wire[31:0] addr_14583_7;

Selector_2 s14583_7(wires_3645_6[3], addr_3645_6, addr_positional[58335:58332], addr_14583_7);

wire[31:0] addr_14584_7;

Selector_2 s14584_7(wires_3646_6[0], addr_3646_6, addr_positional[58339:58336], addr_14584_7);

wire[31:0] addr_14585_7;

Selector_2 s14585_7(wires_3646_6[1], addr_3646_6, addr_positional[58343:58340], addr_14585_7);

wire[31:0] addr_14586_7;

Selector_2 s14586_7(wires_3646_6[2], addr_3646_6, addr_positional[58347:58344], addr_14586_7);

wire[31:0] addr_14587_7;

Selector_2 s14587_7(wires_3646_6[3], addr_3646_6, addr_positional[58351:58348], addr_14587_7);

wire[31:0] addr_14588_7;

Selector_2 s14588_7(wires_3647_6[0], addr_3647_6, addr_positional[58355:58352], addr_14588_7);

wire[31:0] addr_14589_7;

Selector_2 s14589_7(wires_3647_6[1], addr_3647_6, addr_positional[58359:58356], addr_14589_7);

wire[31:0] addr_14590_7;

Selector_2 s14590_7(wires_3647_6[2], addr_3647_6, addr_positional[58363:58360], addr_14590_7);

wire[31:0] addr_14591_7;

Selector_2 s14591_7(wires_3647_6[3], addr_3647_6, addr_positional[58367:58364], addr_14591_7);

wire[31:0] addr_14592_7;

Selector_2 s14592_7(wires_3648_6[0], addr_3648_6, addr_positional[58371:58368], addr_14592_7);

wire[31:0] addr_14593_7;

Selector_2 s14593_7(wires_3648_6[1], addr_3648_6, addr_positional[58375:58372], addr_14593_7);

wire[31:0] addr_14594_7;

Selector_2 s14594_7(wires_3648_6[2], addr_3648_6, addr_positional[58379:58376], addr_14594_7);

wire[31:0] addr_14595_7;

Selector_2 s14595_7(wires_3648_6[3], addr_3648_6, addr_positional[58383:58380], addr_14595_7);

wire[31:0] addr_14596_7;

Selector_2 s14596_7(wires_3649_6[0], addr_3649_6, addr_positional[58387:58384], addr_14596_7);

wire[31:0] addr_14597_7;

Selector_2 s14597_7(wires_3649_6[1], addr_3649_6, addr_positional[58391:58388], addr_14597_7);

wire[31:0] addr_14598_7;

Selector_2 s14598_7(wires_3649_6[2], addr_3649_6, addr_positional[58395:58392], addr_14598_7);

wire[31:0] addr_14599_7;

Selector_2 s14599_7(wires_3649_6[3], addr_3649_6, addr_positional[58399:58396], addr_14599_7);

wire[31:0] addr_14600_7;

Selector_2 s14600_7(wires_3650_6[0], addr_3650_6, addr_positional[58403:58400], addr_14600_7);

wire[31:0] addr_14601_7;

Selector_2 s14601_7(wires_3650_6[1], addr_3650_6, addr_positional[58407:58404], addr_14601_7);

wire[31:0] addr_14602_7;

Selector_2 s14602_7(wires_3650_6[2], addr_3650_6, addr_positional[58411:58408], addr_14602_7);

wire[31:0] addr_14603_7;

Selector_2 s14603_7(wires_3650_6[3], addr_3650_6, addr_positional[58415:58412], addr_14603_7);

wire[31:0] addr_14604_7;

Selector_2 s14604_7(wires_3651_6[0], addr_3651_6, addr_positional[58419:58416], addr_14604_7);

wire[31:0] addr_14605_7;

Selector_2 s14605_7(wires_3651_6[1], addr_3651_6, addr_positional[58423:58420], addr_14605_7);

wire[31:0] addr_14606_7;

Selector_2 s14606_7(wires_3651_6[2], addr_3651_6, addr_positional[58427:58424], addr_14606_7);

wire[31:0] addr_14607_7;

Selector_2 s14607_7(wires_3651_6[3], addr_3651_6, addr_positional[58431:58428], addr_14607_7);

wire[31:0] addr_14608_7;

Selector_2 s14608_7(wires_3652_6[0], addr_3652_6, addr_positional[58435:58432], addr_14608_7);

wire[31:0] addr_14609_7;

Selector_2 s14609_7(wires_3652_6[1], addr_3652_6, addr_positional[58439:58436], addr_14609_7);

wire[31:0] addr_14610_7;

Selector_2 s14610_7(wires_3652_6[2], addr_3652_6, addr_positional[58443:58440], addr_14610_7);

wire[31:0] addr_14611_7;

Selector_2 s14611_7(wires_3652_6[3], addr_3652_6, addr_positional[58447:58444], addr_14611_7);

wire[31:0] addr_14612_7;

Selector_2 s14612_7(wires_3653_6[0], addr_3653_6, addr_positional[58451:58448], addr_14612_7);

wire[31:0] addr_14613_7;

Selector_2 s14613_7(wires_3653_6[1], addr_3653_6, addr_positional[58455:58452], addr_14613_7);

wire[31:0] addr_14614_7;

Selector_2 s14614_7(wires_3653_6[2], addr_3653_6, addr_positional[58459:58456], addr_14614_7);

wire[31:0] addr_14615_7;

Selector_2 s14615_7(wires_3653_6[3], addr_3653_6, addr_positional[58463:58460], addr_14615_7);

wire[31:0] addr_14616_7;

Selector_2 s14616_7(wires_3654_6[0], addr_3654_6, addr_positional[58467:58464], addr_14616_7);

wire[31:0] addr_14617_7;

Selector_2 s14617_7(wires_3654_6[1], addr_3654_6, addr_positional[58471:58468], addr_14617_7);

wire[31:0] addr_14618_7;

Selector_2 s14618_7(wires_3654_6[2], addr_3654_6, addr_positional[58475:58472], addr_14618_7);

wire[31:0] addr_14619_7;

Selector_2 s14619_7(wires_3654_6[3], addr_3654_6, addr_positional[58479:58476], addr_14619_7);

wire[31:0] addr_14620_7;

Selector_2 s14620_7(wires_3655_6[0], addr_3655_6, addr_positional[58483:58480], addr_14620_7);

wire[31:0] addr_14621_7;

Selector_2 s14621_7(wires_3655_6[1], addr_3655_6, addr_positional[58487:58484], addr_14621_7);

wire[31:0] addr_14622_7;

Selector_2 s14622_7(wires_3655_6[2], addr_3655_6, addr_positional[58491:58488], addr_14622_7);

wire[31:0] addr_14623_7;

Selector_2 s14623_7(wires_3655_6[3], addr_3655_6, addr_positional[58495:58492], addr_14623_7);

wire[31:0] addr_14624_7;

Selector_2 s14624_7(wires_3656_6[0], addr_3656_6, addr_positional[58499:58496], addr_14624_7);

wire[31:0] addr_14625_7;

Selector_2 s14625_7(wires_3656_6[1], addr_3656_6, addr_positional[58503:58500], addr_14625_7);

wire[31:0] addr_14626_7;

Selector_2 s14626_7(wires_3656_6[2], addr_3656_6, addr_positional[58507:58504], addr_14626_7);

wire[31:0] addr_14627_7;

Selector_2 s14627_7(wires_3656_6[3], addr_3656_6, addr_positional[58511:58508], addr_14627_7);

wire[31:0] addr_14628_7;

Selector_2 s14628_7(wires_3657_6[0], addr_3657_6, addr_positional[58515:58512], addr_14628_7);

wire[31:0] addr_14629_7;

Selector_2 s14629_7(wires_3657_6[1], addr_3657_6, addr_positional[58519:58516], addr_14629_7);

wire[31:0] addr_14630_7;

Selector_2 s14630_7(wires_3657_6[2], addr_3657_6, addr_positional[58523:58520], addr_14630_7);

wire[31:0] addr_14631_7;

Selector_2 s14631_7(wires_3657_6[3], addr_3657_6, addr_positional[58527:58524], addr_14631_7);

wire[31:0] addr_14632_7;

Selector_2 s14632_7(wires_3658_6[0], addr_3658_6, addr_positional[58531:58528], addr_14632_7);

wire[31:0] addr_14633_7;

Selector_2 s14633_7(wires_3658_6[1], addr_3658_6, addr_positional[58535:58532], addr_14633_7);

wire[31:0] addr_14634_7;

Selector_2 s14634_7(wires_3658_6[2], addr_3658_6, addr_positional[58539:58536], addr_14634_7);

wire[31:0] addr_14635_7;

Selector_2 s14635_7(wires_3658_6[3], addr_3658_6, addr_positional[58543:58540], addr_14635_7);

wire[31:0] addr_14636_7;

Selector_2 s14636_7(wires_3659_6[0], addr_3659_6, addr_positional[58547:58544], addr_14636_7);

wire[31:0] addr_14637_7;

Selector_2 s14637_7(wires_3659_6[1], addr_3659_6, addr_positional[58551:58548], addr_14637_7);

wire[31:0] addr_14638_7;

Selector_2 s14638_7(wires_3659_6[2], addr_3659_6, addr_positional[58555:58552], addr_14638_7);

wire[31:0] addr_14639_7;

Selector_2 s14639_7(wires_3659_6[3], addr_3659_6, addr_positional[58559:58556], addr_14639_7);

wire[31:0] addr_14640_7;

Selector_2 s14640_7(wires_3660_6[0], addr_3660_6, addr_positional[58563:58560], addr_14640_7);

wire[31:0] addr_14641_7;

Selector_2 s14641_7(wires_3660_6[1], addr_3660_6, addr_positional[58567:58564], addr_14641_7);

wire[31:0] addr_14642_7;

Selector_2 s14642_7(wires_3660_6[2], addr_3660_6, addr_positional[58571:58568], addr_14642_7);

wire[31:0] addr_14643_7;

Selector_2 s14643_7(wires_3660_6[3], addr_3660_6, addr_positional[58575:58572], addr_14643_7);

wire[31:0] addr_14644_7;

Selector_2 s14644_7(wires_3661_6[0], addr_3661_6, addr_positional[58579:58576], addr_14644_7);

wire[31:0] addr_14645_7;

Selector_2 s14645_7(wires_3661_6[1], addr_3661_6, addr_positional[58583:58580], addr_14645_7);

wire[31:0] addr_14646_7;

Selector_2 s14646_7(wires_3661_6[2], addr_3661_6, addr_positional[58587:58584], addr_14646_7);

wire[31:0] addr_14647_7;

Selector_2 s14647_7(wires_3661_6[3], addr_3661_6, addr_positional[58591:58588], addr_14647_7);

wire[31:0] addr_14648_7;

Selector_2 s14648_7(wires_3662_6[0], addr_3662_6, addr_positional[58595:58592], addr_14648_7);

wire[31:0] addr_14649_7;

Selector_2 s14649_7(wires_3662_6[1], addr_3662_6, addr_positional[58599:58596], addr_14649_7);

wire[31:0] addr_14650_7;

Selector_2 s14650_7(wires_3662_6[2], addr_3662_6, addr_positional[58603:58600], addr_14650_7);

wire[31:0] addr_14651_7;

Selector_2 s14651_7(wires_3662_6[3], addr_3662_6, addr_positional[58607:58604], addr_14651_7);

wire[31:0] addr_14652_7;

Selector_2 s14652_7(wires_3663_6[0], addr_3663_6, addr_positional[58611:58608], addr_14652_7);

wire[31:0] addr_14653_7;

Selector_2 s14653_7(wires_3663_6[1], addr_3663_6, addr_positional[58615:58612], addr_14653_7);

wire[31:0] addr_14654_7;

Selector_2 s14654_7(wires_3663_6[2], addr_3663_6, addr_positional[58619:58616], addr_14654_7);

wire[31:0] addr_14655_7;

Selector_2 s14655_7(wires_3663_6[3], addr_3663_6, addr_positional[58623:58620], addr_14655_7);

wire[31:0] addr_14656_7;

Selector_2 s14656_7(wires_3664_6[0], addr_3664_6, addr_positional[58627:58624], addr_14656_7);

wire[31:0] addr_14657_7;

Selector_2 s14657_7(wires_3664_6[1], addr_3664_6, addr_positional[58631:58628], addr_14657_7);

wire[31:0] addr_14658_7;

Selector_2 s14658_7(wires_3664_6[2], addr_3664_6, addr_positional[58635:58632], addr_14658_7);

wire[31:0] addr_14659_7;

Selector_2 s14659_7(wires_3664_6[3], addr_3664_6, addr_positional[58639:58636], addr_14659_7);

wire[31:0] addr_14660_7;

Selector_2 s14660_7(wires_3665_6[0], addr_3665_6, addr_positional[58643:58640], addr_14660_7);

wire[31:0] addr_14661_7;

Selector_2 s14661_7(wires_3665_6[1], addr_3665_6, addr_positional[58647:58644], addr_14661_7);

wire[31:0] addr_14662_7;

Selector_2 s14662_7(wires_3665_6[2], addr_3665_6, addr_positional[58651:58648], addr_14662_7);

wire[31:0] addr_14663_7;

Selector_2 s14663_7(wires_3665_6[3], addr_3665_6, addr_positional[58655:58652], addr_14663_7);

wire[31:0] addr_14664_7;

Selector_2 s14664_7(wires_3666_6[0], addr_3666_6, addr_positional[58659:58656], addr_14664_7);

wire[31:0] addr_14665_7;

Selector_2 s14665_7(wires_3666_6[1], addr_3666_6, addr_positional[58663:58660], addr_14665_7);

wire[31:0] addr_14666_7;

Selector_2 s14666_7(wires_3666_6[2], addr_3666_6, addr_positional[58667:58664], addr_14666_7);

wire[31:0] addr_14667_7;

Selector_2 s14667_7(wires_3666_6[3], addr_3666_6, addr_positional[58671:58668], addr_14667_7);

wire[31:0] addr_14668_7;

Selector_2 s14668_7(wires_3667_6[0], addr_3667_6, addr_positional[58675:58672], addr_14668_7);

wire[31:0] addr_14669_7;

Selector_2 s14669_7(wires_3667_6[1], addr_3667_6, addr_positional[58679:58676], addr_14669_7);

wire[31:0] addr_14670_7;

Selector_2 s14670_7(wires_3667_6[2], addr_3667_6, addr_positional[58683:58680], addr_14670_7);

wire[31:0] addr_14671_7;

Selector_2 s14671_7(wires_3667_6[3], addr_3667_6, addr_positional[58687:58684], addr_14671_7);

wire[31:0] addr_14672_7;

Selector_2 s14672_7(wires_3668_6[0], addr_3668_6, addr_positional[58691:58688], addr_14672_7);

wire[31:0] addr_14673_7;

Selector_2 s14673_7(wires_3668_6[1], addr_3668_6, addr_positional[58695:58692], addr_14673_7);

wire[31:0] addr_14674_7;

Selector_2 s14674_7(wires_3668_6[2], addr_3668_6, addr_positional[58699:58696], addr_14674_7);

wire[31:0] addr_14675_7;

Selector_2 s14675_7(wires_3668_6[3], addr_3668_6, addr_positional[58703:58700], addr_14675_7);

wire[31:0] addr_14676_7;

Selector_2 s14676_7(wires_3669_6[0], addr_3669_6, addr_positional[58707:58704], addr_14676_7);

wire[31:0] addr_14677_7;

Selector_2 s14677_7(wires_3669_6[1], addr_3669_6, addr_positional[58711:58708], addr_14677_7);

wire[31:0] addr_14678_7;

Selector_2 s14678_7(wires_3669_6[2], addr_3669_6, addr_positional[58715:58712], addr_14678_7);

wire[31:0] addr_14679_7;

Selector_2 s14679_7(wires_3669_6[3], addr_3669_6, addr_positional[58719:58716], addr_14679_7);

wire[31:0] addr_14680_7;

Selector_2 s14680_7(wires_3670_6[0], addr_3670_6, addr_positional[58723:58720], addr_14680_7);

wire[31:0] addr_14681_7;

Selector_2 s14681_7(wires_3670_6[1], addr_3670_6, addr_positional[58727:58724], addr_14681_7);

wire[31:0] addr_14682_7;

Selector_2 s14682_7(wires_3670_6[2], addr_3670_6, addr_positional[58731:58728], addr_14682_7);

wire[31:0] addr_14683_7;

Selector_2 s14683_7(wires_3670_6[3], addr_3670_6, addr_positional[58735:58732], addr_14683_7);

wire[31:0] addr_14684_7;

Selector_2 s14684_7(wires_3671_6[0], addr_3671_6, addr_positional[58739:58736], addr_14684_7);

wire[31:0] addr_14685_7;

Selector_2 s14685_7(wires_3671_6[1], addr_3671_6, addr_positional[58743:58740], addr_14685_7);

wire[31:0] addr_14686_7;

Selector_2 s14686_7(wires_3671_6[2], addr_3671_6, addr_positional[58747:58744], addr_14686_7);

wire[31:0] addr_14687_7;

Selector_2 s14687_7(wires_3671_6[3], addr_3671_6, addr_positional[58751:58748], addr_14687_7);

wire[31:0] addr_14688_7;

Selector_2 s14688_7(wires_3672_6[0], addr_3672_6, addr_positional[58755:58752], addr_14688_7);

wire[31:0] addr_14689_7;

Selector_2 s14689_7(wires_3672_6[1], addr_3672_6, addr_positional[58759:58756], addr_14689_7);

wire[31:0] addr_14690_7;

Selector_2 s14690_7(wires_3672_6[2], addr_3672_6, addr_positional[58763:58760], addr_14690_7);

wire[31:0] addr_14691_7;

Selector_2 s14691_7(wires_3672_6[3], addr_3672_6, addr_positional[58767:58764], addr_14691_7);

wire[31:0] addr_14692_7;

Selector_2 s14692_7(wires_3673_6[0], addr_3673_6, addr_positional[58771:58768], addr_14692_7);

wire[31:0] addr_14693_7;

Selector_2 s14693_7(wires_3673_6[1], addr_3673_6, addr_positional[58775:58772], addr_14693_7);

wire[31:0] addr_14694_7;

Selector_2 s14694_7(wires_3673_6[2], addr_3673_6, addr_positional[58779:58776], addr_14694_7);

wire[31:0] addr_14695_7;

Selector_2 s14695_7(wires_3673_6[3], addr_3673_6, addr_positional[58783:58780], addr_14695_7);

wire[31:0] addr_14696_7;

Selector_2 s14696_7(wires_3674_6[0], addr_3674_6, addr_positional[58787:58784], addr_14696_7);

wire[31:0] addr_14697_7;

Selector_2 s14697_7(wires_3674_6[1], addr_3674_6, addr_positional[58791:58788], addr_14697_7);

wire[31:0] addr_14698_7;

Selector_2 s14698_7(wires_3674_6[2], addr_3674_6, addr_positional[58795:58792], addr_14698_7);

wire[31:0] addr_14699_7;

Selector_2 s14699_7(wires_3674_6[3], addr_3674_6, addr_positional[58799:58796], addr_14699_7);

wire[31:0] addr_14700_7;

Selector_2 s14700_7(wires_3675_6[0], addr_3675_6, addr_positional[58803:58800], addr_14700_7);

wire[31:0] addr_14701_7;

Selector_2 s14701_7(wires_3675_6[1], addr_3675_6, addr_positional[58807:58804], addr_14701_7);

wire[31:0] addr_14702_7;

Selector_2 s14702_7(wires_3675_6[2], addr_3675_6, addr_positional[58811:58808], addr_14702_7);

wire[31:0] addr_14703_7;

Selector_2 s14703_7(wires_3675_6[3], addr_3675_6, addr_positional[58815:58812], addr_14703_7);

wire[31:0] addr_14704_7;

Selector_2 s14704_7(wires_3676_6[0], addr_3676_6, addr_positional[58819:58816], addr_14704_7);

wire[31:0] addr_14705_7;

Selector_2 s14705_7(wires_3676_6[1], addr_3676_6, addr_positional[58823:58820], addr_14705_7);

wire[31:0] addr_14706_7;

Selector_2 s14706_7(wires_3676_6[2], addr_3676_6, addr_positional[58827:58824], addr_14706_7);

wire[31:0] addr_14707_7;

Selector_2 s14707_7(wires_3676_6[3], addr_3676_6, addr_positional[58831:58828], addr_14707_7);

wire[31:0] addr_14708_7;

Selector_2 s14708_7(wires_3677_6[0], addr_3677_6, addr_positional[58835:58832], addr_14708_7);

wire[31:0] addr_14709_7;

Selector_2 s14709_7(wires_3677_6[1], addr_3677_6, addr_positional[58839:58836], addr_14709_7);

wire[31:0] addr_14710_7;

Selector_2 s14710_7(wires_3677_6[2], addr_3677_6, addr_positional[58843:58840], addr_14710_7);

wire[31:0] addr_14711_7;

Selector_2 s14711_7(wires_3677_6[3], addr_3677_6, addr_positional[58847:58844], addr_14711_7);

wire[31:0] addr_14712_7;

Selector_2 s14712_7(wires_3678_6[0], addr_3678_6, addr_positional[58851:58848], addr_14712_7);

wire[31:0] addr_14713_7;

Selector_2 s14713_7(wires_3678_6[1], addr_3678_6, addr_positional[58855:58852], addr_14713_7);

wire[31:0] addr_14714_7;

Selector_2 s14714_7(wires_3678_6[2], addr_3678_6, addr_positional[58859:58856], addr_14714_7);

wire[31:0] addr_14715_7;

Selector_2 s14715_7(wires_3678_6[3], addr_3678_6, addr_positional[58863:58860], addr_14715_7);

wire[31:0] addr_14716_7;

Selector_2 s14716_7(wires_3679_6[0], addr_3679_6, addr_positional[58867:58864], addr_14716_7);

wire[31:0] addr_14717_7;

Selector_2 s14717_7(wires_3679_6[1], addr_3679_6, addr_positional[58871:58868], addr_14717_7);

wire[31:0] addr_14718_7;

Selector_2 s14718_7(wires_3679_6[2], addr_3679_6, addr_positional[58875:58872], addr_14718_7);

wire[31:0] addr_14719_7;

Selector_2 s14719_7(wires_3679_6[3], addr_3679_6, addr_positional[58879:58876], addr_14719_7);

wire[31:0] addr_14720_7;

Selector_2 s14720_7(wires_3680_6[0], addr_3680_6, addr_positional[58883:58880], addr_14720_7);

wire[31:0] addr_14721_7;

Selector_2 s14721_7(wires_3680_6[1], addr_3680_6, addr_positional[58887:58884], addr_14721_7);

wire[31:0] addr_14722_7;

Selector_2 s14722_7(wires_3680_6[2], addr_3680_6, addr_positional[58891:58888], addr_14722_7);

wire[31:0] addr_14723_7;

Selector_2 s14723_7(wires_3680_6[3], addr_3680_6, addr_positional[58895:58892], addr_14723_7);

wire[31:0] addr_14724_7;

Selector_2 s14724_7(wires_3681_6[0], addr_3681_6, addr_positional[58899:58896], addr_14724_7);

wire[31:0] addr_14725_7;

Selector_2 s14725_7(wires_3681_6[1], addr_3681_6, addr_positional[58903:58900], addr_14725_7);

wire[31:0] addr_14726_7;

Selector_2 s14726_7(wires_3681_6[2], addr_3681_6, addr_positional[58907:58904], addr_14726_7);

wire[31:0] addr_14727_7;

Selector_2 s14727_7(wires_3681_6[3], addr_3681_6, addr_positional[58911:58908], addr_14727_7);

wire[31:0] addr_14728_7;

Selector_2 s14728_7(wires_3682_6[0], addr_3682_6, addr_positional[58915:58912], addr_14728_7);

wire[31:0] addr_14729_7;

Selector_2 s14729_7(wires_3682_6[1], addr_3682_6, addr_positional[58919:58916], addr_14729_7);

wire[31:0] addr_14730_7;

Selector_2 s14730_7(wires_3682_6[2], addr_3682_6, addr_positional[58923:58920], addr_14730_7);

wire[31:0] addr_14731_7;

Selector_2 s14731_7(wires_3682_6[3], addr_3682_6, addr_positional[58927:58924], addr_14731_7);

wire[31:0] addr_14732_7;

Selector_2 s14732_7(wires_3683_6[0], addr_3683_6, addr_positional[58931:58928], addr_14732_7);

wire[31:0] addr_14733_7;

Selector_2 s14733_7(wires_3683_6[1], addr_3683_6, addr_positional[58935:58932], addr_14733_7);

wire[31:0] addr_14734_7;

Selector_2 s14734_7(wires_3683_6[2], addr_3683_6, addr_positional[58939:58936], addr_14734_7);

wire[31:0] addr_14735_7;

Selector_2 s14735_7(wires_3683_6[3], addr_3683_6, addr_positional[58943:58940], addr_14735_7);

wire[31:0] addr_14736_7;

Selector_2 s14736_7(wires_3684_6[0], addr_3684_6, addr_positional[58947:58944], addr_14736_7);

wire[31:0] addr_14737_7;

Selector_2 s14737_7(wires_3684_6[1], addr_3684_6, addr_positional[58951:58948], addr_14737_7);

wire[31:0] addr_14738_7;

Selector_2 s14738_7(wires_3684_6[2], addr_3684_6, addr_positional[58955:58952], addr_14738_7);

wire[31:0] addr_14739_7;

Selector_2 s14739_7(wires_3684_6[3], addr_3684_6, addr_positional[58959:58956], addr_14739_7);

wire[31:0] addr_14740_7;

Selector_2 s14740_7(wires_3685_6[0], addr_3685_6, addr_positional[58963:58960], addr_14740_7);

wire[31:0] addr_14741_7;

Selector_2 s14741_7(wires_3685_6[1], addr_3685_6, addr_positional[58967:58964], addr_14741_7);

wire[31:0] addr_14742_7;

Selector_2 s14742_7(wires_3685_6[2], addr_3685_6, addr_positional[58971:58968], addr_14742_7);

wire[31:0] addr_14743_7;

Selector_2 s14743_7(wires_3685_6[3], addr_3685_6, addr_positional[58975:58972], addr_14743_7);

wire[31:0] addr_14744_7;

Selector_2 s14744_7(wires_3686_6[0], addr_3686_6, addr_positional[58979:58976], addr_14744_7);

wire[31:0] addr_14745_7;

Selector_2 s14745_7(wires_3686_6[1], addr_3686_6, addr_positional[58983:58980], addr_14745_7);

wire[31:0] addr_14746_7;

Selector_2 s14746_7(wires_3686_6[2], addr_3686_6, addr_positional[58987:58984], addr_14746_7);

wire[31:0] addr_14747_7;

Selector_2 s14747_7(wires_3686_6[3], addr_3686_6, addr_positional[58991:58988], addr_14747_7);

wire[31:0] addr_14748_7;

Selector_2 s14748_7(wires_3687_6[0], addr_3687_6, addr_positional[58995:58992], addr_14748_7);

wire[31:0] addr_14749_7;

Selector_2 s14749_7(wires_3687_6[1], addr_3687_6, addr_positional[58999:58996], addr_14749_7);

wire[31:0] addr_14750_7;

Selector_2 s14750_7(wires_3687_6[2], addr_3687_6, addr_positional[59003:59000], addr_14750_7);

wire[31:0] addr_14751_7;

Selector_2 s14751_7(wires_3687_6[3], addr_3687_6, addr_positional[59007:59004], addr_14751_7);

wire[31:0] addr_14752_7;

Selector_2 s14752_7(wires_3688_6[0], addr_3688_6, addr_positional[59011:59008], addr_14752_7);

wire[31:0] addr_14753_7;

Selector_2 s14753_7(wires_3688_6[1], addr_3688_6, addr_positional[59015:59012], addr_14753_7);

wire[31:0] addr_14754_7;

Selector_2 s14754_7(wires_3688_6[2], addr_3688_6, addr_positional[59019:59016], addr_14754_7);

wire[31:0] addr_14755_7;

Selector_2 s14755_7(wires_3688_6[3], addr_3688_6, addr_positional[59023:59020], addr_14755_7);

wire[31:0] addr_14756_7;

Selector_2 s14756_7(wires_3689_6[0], addr_3689_6, addr_positional[59027:59024], addr_14756_7);

wire[31:0] addr_14757_7;

Selector_2 s14757_7(wires_3689_6[1], addr_3689_6, addr_positional[59031:59028], addr_14757_7);

wire[31:0] addr_14758_7;

Selector_2 s14758_7(wires_3689_6[2], addr_3689_6, addr_positional[59035:59032], addr_14758_7);

wire[31:0] addr_14759_7;

Selector_2 s14759_7(wires_3689_6[3], addr_3689_6, addr_positional[59039:59036], addr_14759_7);

wire[31:0] addr_14760_7;

Selector_2 s14760_7(wires_3690_6[0], addr_3690_6, addr_positional[59043:59040], addr_14760_7);

wire[31:0] addr_14761_7;

Selector_2 s14761_7(wires_3690_6[1], addr_3690_6, addr_positional[59047:59044], addr_14761_7);

wire[31:0] addr_14762_7;

Selector_2 s14762_7(wires_3690_6[2], addr_3690_6, addr_positional[59051:59048], addr_14762_7);

wire[31:0] addr_14763_7;

Selector_2 s14763_7(wires_3690_6[3], addr_3690_6, addr_positional[59055:59052], addr_14763_7);

wire[31:0] addr_14764_7;

Selector_2 s14764_7(wires_3691_6[0], addr_3691_6, addr_positional[59059:59056], addr_14764_7);

wire[31:0] addr_14765_7;

Selector_2 s14765_7(wires_3691_6[1], addr_3691_6, addr_positional[59063:59060], addr_14765_7);

wire[31:0] addr_14766_7;

Selector_2 s14766_7(wires_3691_6[2], addr_3691_6, addr_positional[59067:59064], addr_14766_7);

wire[31:0] addr_14767_7;

Selector_2 s14767_7(wires_3691_6[3], addr_3691_6, addr_positional[59071:59068], addr_14767_7);

wire[31:0] addr_14768_7;

Selector_2 s14768_7(wires_3692_6[0], addr_3692_6, addr_positional[59075:59072], addr_14768_7);

wire[31:0] addr_14769_7;

Selector_2 s14769_7(wires_3692_6[1], addr_3692_6, addr_positional[59079:59076], addr_14769_7);

wire[31:0] addr_14770_7;

Selector_2 s14770_7(wires_3692_6[2], addr_3692_6, addr_positional[59083:59080], addr_14770_7);

wire[31:0] addr_14771_7;

Selector_2 s14771_7(wires_3692_6[3], addr_3692_6, addr_positional[59087:59084], addr_14771_7);

wire[31:0] addr_14772_7;

Selector_2 s14772_7(wires_3693_6[0], addr_3693_6, addr_positional[59091:59088], addr_14772_7);

wire[31:0] addr_14773_7;

Selector_2 s14773_7(wires_3693_6[1], addr_3693_6, addr_positional[59095:59092], addr_14773_7);

wire[31:0] addr_14774_7;

Selector_2 s14774_7(wires_3693_6[2], addr_3693_6, addr_positional[59099:59096], addr_14774_7);

wire[31:0] addr_14775_7;

Selector_2 s14775_7(wires_3693_6[3], addr_3693_6, addr_positional[59103:59100], addr_14775_7);

wire[31:0] addr_14776_7;

Selector_2 s14776_7(wires_3694_6[0], addr_3694_6, addr_positional[59107:59104], addr_14776_7);

wire[31:0] addr_14777_7;

Selector_2 s14777_7(wires_3694_6[1], addr_3694_6, addr_positional[59111:59108], addr_14777_7);

wire[31:0] addr_14778_7;

Selector_2 s14778_7(wires_3694_6[2], addr_3694_6, addr_positional[59115:59112], addr_14778_7);

wire[31:0] addr_14779_7;

Selector_2 s14779_7(wires_3694_6[3], addr_3694_6, addr_positional[59119:59116], addr_14779_7);

wire[31:0] addr_14780_7;

Selector_2 s14780_7(wires_3695_6[0], addr_3695_6, addr_positional[59123:59120], addr_14780_7);

wire[31:0] addr_14781_7;

Selector_2 s14781_7(wires_3695_6[1], addr_3695_6, addr_positional[59127:59124], addr_14781_7);

wire[31:0] addr_14782_7;

Selector_2 s14782_7(wires_3695_6[2], addr_3695_6, addr_positional[59131:59128], addr_14782_7);

wire[31:0] addr_14783_7;

Selector_2 s14783_7(wires_3695_6[3], addr_3695_6, addr_positional[59135:59132], addr_14783_7);

wire[31:0] addr_14784_7;

Selector_2 s14784_7(wires_3696_6[0], addr_3696_6, addr_positional[59139:59136], addr_14784_7);

wire[31:0] addr_14785_7;

Selector_2 s14785_7(wires_3696_6[1], addr_3696_6, addr_positional[59143:59140], addr_14785_7);

wire[31:0] addr_14786_7;

Selector_2 s14786_7(wires_3696_6[2], addr_3696_6, addr_positional[59147:59144], addr_14786_7);

wire[31:0] addr_14787_7;

Selector_2 s14787_7(wires_3696_6[3], addr_3696_6, addr_positional[59151:59148], addr_14787_7);

wire[31:0] addr_14788_7;

Selector_2 s14788_7(wires_3697_6[0], addr_3697_6, addr_positional[59155:59152], addr_14788_7);

wire[31:0] addr_14789_7;

Selector_2 s14789_7(wires_3697_6[1], addr_3697_6, addr_positional[59159:59156], addr_14789_7);

wire[31:0] addr_14790_7;

Selector_2 s14790_7(wires_3697_6[2], addr_3697_6, addr_positional[59163:59160], addr_14790_7);

wire[31:0] addr_14791_7;

Selector_2 s14791_7(wires_3697_6[3], addr_3697_6, addr_positional[59167:59164], addr_14791_7);

wire[31:0] addr_14792_7;

Selector_2 s14792_7(wires_3698_6[0], addr_3698_6, addr_positional[59171:59168], addr_14792_7);

wire[31:0] addr_14793_7;

Selector_2 s14793_7(wires_3698_6[1], addr_3698_6, addr_positional[59175:59172], addr_14793_7);

wire[31:0] addr_14794_7;

Selector_2 s14794_7(wires_3698_6[2], addr_3698_6, addr_positional[59179:59176], addr_14794_7);

wire[31:0] addr_14795_7;

Selector_2 s14795_7(wires_3698_6[3], addr_3698_6, addr_positional[59183:59180], addr_14795_7);

wire[31:0] addr_14796_7;

Selector_2 s14796_7(wires_3699_6[0], addr_3699_6, addr_positional[59187:59184], addr_14796_7);

wire[31:0] addr_14797_7;

Selector_2 s14797_7(wires_3699_6[1], addr_3699_6, addr_positional[59191:59188], addr_14797_7);

wire[31:0] addr_14798_7;

Selector_2 s14798_7(wires_3699_6[2], addr_3699_6, addr_positional[59195:59192], addr_14798_7);

wire[31:0] addr_14799_7;

Selector_2 s14799_7(wires_3699_6[3], addr_3699_6, addr_positional[59199:59196], addr_14799_7);

wire[31:0] addr_14800_7;

Selector_2 s14800_7(wires_3700_6[0], addr_3700_6, addr_positional[59203:59200], addr_14800_7);

wire[31:0] addr_14801_7;

Selector_2 s14801_7(wires_3700_6[1], addr_3700_6, addr_positional[59207:59204], addr_14801_7);

wire[31:0] addr_14802_7;

Selector_2 s14802_7(wires_3700_6[2], addr_3700_6, addr_positional[59211:59208], addr_14802_7);

wire[31:0] addr_14803_7;

Selector_2 s14803_7(wires_3700_6[3], addr_3700_6, addr_positional[59215:59212], addr_14803_7);

wire[31:0] addr_14804_7;

Selector_2 s14804_7(wires_3701_6[0], addr_3701_6, addr_positional[59219:59216], addr_14804_7);

wire[31:0] addr_14805_7;

Selector_2 s14805_7(wires_3701_6[1], addr_3701_6, addr_positional[59223:59220], addr_14805_7);

wire[31:0] addr_14806_7;

Selector_2 s14806_7(wires_3701_6[2], addr_3701_6, addr_positional[59227:59224], addr_14806_7);

wire[31:0] addr_14807_7;

Selector_2 s14807_7(wires_3701_6[3], addr_3701_6, addr_positional[59231:59228], addr_14807_7);

wire[31:0] addr_14808_7;

Selector_2 s14808_7(wires_3702_6[0], addr_3702_6, addr_positional[59235:59232], addr_14808_7);

wire[31:0] addr_14809_7;

Selector_2 s14809_7(wires_3702_6[1], addr_3702_6, addr_positional[59239:59236], addr_14809_7);

wire[31:0] addr_14810_7;

Selector_2 s14810_7(wires_3702_6[2], addr_3702_6, addr_positional[59243:59240], addr_14810_7);

wire[31:0] addr_14811_7;

Selector_2 s14811_7(wires_3702_6[3], addr_3702_6, addr_positional[59247:59244], addr_14811_7);

wire[31:0] addr_14812_7;

Selector_2 s14812_7(wires_3703_6[0], addr_3703_6, addr_positional[59251:59248], addr_14812_7);

wire[31:0] addr_14813_7;

Selector_2 s14813_7(wires_3703_6[1], addr_3703_6, addr_positional[59255:59252], addr_14813_7);

wire[31:0] addr_14814_7;

Selector_2 s14814_7(wires_3703_6[2], addr_3703_6, addr_positional[59259:59256], addr_14814_7);

wire[31:0] addr_14815_7;

Selector_2 s14815_7(wires_3703_6[3], addr_3703_6, addr_positional[59263:59260], addr_14815_7);

wire[31:0] addr_14816_7;

Selector_2 s14816_7(wires_3704_6[0], addr_3704_6, addr_positional[59267:59264], addr_14816_7);

wire[31:0] addr_14817_7;

Selector_2 s14817_7(wires_3704_6[1], addr_3704_6, addr_positional[59271:59268], addr_14817_7);

wire[31:0] addr_14818_7;

Selector_2 s14818_7(wires_3704_6[2], addr_3704_6, addr_positional[59275:59272], addr_14818_7);

wire[31:0] addr_14819_7;

Selector_2 s14819_7(wires_3704_6[3], addr_3704_6, addr_positional[59279:59276], addr_14819_7);

wire[31:0] addr_14820_7;

Selector_2 s14820_7(wires_3705_6[0], addr_3705_6, addr_positional[59283:59280], addr_14820_7);

wire[31:0] addr_14821_7;

Selector_2 s14821_7(wires_3705_6[1], addr_3705_6, addr_positional[59287:59284], addr_14821_7);

wire[31:0] addr_14822_7;

Selector_2 s14822_7(wires_3705_6[2], addr_3705_6, addr_positional[59291:59288], addr_14822_7);

wire[31:0] addr_14823_7;

Selector_2 s14823_7(wires_3705_6[3], addr_3705_6, addr_positional[59295:59292], addr_14823_7);

wire[31:0] addr_14824_7;

Selector_2 s14824_7(wires_3706_6[0], addr_3706_6, addr_positional[59299:59296], addr_14824_7);

wire[31:0] addr_14825_7;

Selector_2 s14825_7(wires_3706_6[1], addr_3706_6, addr_positional[59303:59300], addr_14825_7);

wire[31:0] addr_14826_7;

Selector_2 s14826_7(wires_3706_6[2], addr_3706_6, addr_positional[59307:59304], addr_14826_7);

wire[31:0] addr_14827_7;

Selector_2 s14827_7(wires_3706_6[3], addr_3706_6, addr_positional[59311:59308], addr_14827_7);

wire[31:0] addr_14828_7;

Selector_2 s14828_7(wires_3707_6[0], addr_3707_6, addr_positional[59315:59312], addr_14828_7);

wire[31:0] addr_14829_7;

Selector_2 s14829_7(wires_3707_6[1], addr_3707_6, addr_positional[59319:59316], addr_14829_7);

wire[31:0] addr_14830_7;

Selector_2 s14830_7(wires_3707_6[2], addr_3707_6, addr_positional[59323:59320], addr_14830_7);

wire[31:0] addr_14831_7;

Selector_2 s14831_7(wires_3707_6[3], addr_3707_6, addr_positional[59327:59324], addr_14831_7);

wire[31:0] addr_14832_7;

Selector_2 s14832_7(wires_3708_6[0], addr_3708_6, addr_positional[59331:59328], addr_14832_7);

wire[31:0] addr_14833_7;

Selector_2 s14833_7(wires_3708_6[1], addr_3708_6, addr_positional[59335:59332], addr_14833_7);

wire[31:0] addr_14834_7;

Selector_2 s14834_7(wires_3708_6[2], addr_3708_6, addr_positional[59339:59336], addr_14834_7);

wire[31:0] addr_14835_7;

Selector_2 s14835_7(wires_3708_6[3], addr_3708_6, addr_positional[59343:59340], addr_14835_7);

wire[31:0] addr_14836_7;

Selector_2 s14836_7(wires_3709_6[0], addr_3709_6, addr_positional[59347:59344], addr_14836_7);

wire[31:0] addr_14837_7;

Selector_2 s14837_7(wires_3709_6[1], addr_3709_6, addr_positional[59351:59348], addr_14837_7);

wire[31:0] addr_14838_7;

Selector_2 s14838_7(wires_3709_6[2], addr_3709_6, addr_positional[59355:59352], addr_14838_7);

wire[31:0] addr_14839_7;

Selector_2 s14839_7(wires_3709_6[3], addr_3709_6, addr_positional[59359:59356], addr_14839_7);

wire[31:0] addr_14840_7;

Selector_2 s14840_7(wires_3710_6[0], addr_3710_6, addr_positional[59363:59360], addr_14840_7);

wire[31:0] addr_14841_7;

Selector_2 s14841_7(wires_3710_6[1], addr_3710_6, addr_positional[59367:59364], addr_14841_7);

wire[31:0] addr_14842_7;

Selector_2 s14842_7(wires_3710_6[2], addr_3710_6, addr_positional[59371:59368], addr_14842_7);

wire[31:0] addr_14843_7;

Selector_2 s14843_7(wires_3710_6[3], addr_3710_6, addr_positional[59375:59372], addr_14843_7);

wire[31:0] addr_14844_7;

Selector_2 s14844_7(wires_3711_6[0], addr_3711_6, addr_positional[59379:59376], addr_14844_7);

wire[31:0] addr_14845_7;

Selector_2 s14845_7(wires_3711_6[1], addr_3711_6, addr_positional[59383:59380], addr_14845_7);

wire[31:0] addr_14846_7;

Selector_2 s14846_7(wires_3711_6[2], addr_3711_6, addr_positional[59387:59384], addr_14846_7);

wire[31:0] addr_14847_7;

Selector_2 s14847_7(wires_3711_6[3], addr_3711_6, addr_positional[59391:59388], addr_14847_7);

wire[31:0] addr_14848_7;

Selector_2 s14848_7(wires_3712_6[0], addr_3712_6, addr_positional[59395:59392], addr_14848_7);

wire[31:0] addr_14849_7;

Selector_2 s14849_7(wires_3712_6[1], addr_3712_6, addr_positional[59399:59396], addr_14849_7);

wire[31:0] addr_14850_7;

Selector_2 s14850_7(wires_3712_6[2], addr_3712_6, addr_positional[59403:59400], addr_14850_7);

wire[31:0] addr_14851_7;

Selector_2 s14851_7(wires_3712_6[3], addr_3712_6, addr_positional[59407:59404], addr_14851_7);

wire[31:0] addr_14852_7;

Selector_2 s14852_7(wires_3713_6[0], addr_3713_6, addr_positional[59411:59408], addr_14852_7);

wire[31:0] addr_14853_7;

Selector_2 s14853_7(wires_3713_6[1], addr_3713_6, addr_positional[59415:59412], addr_14853_7);

wire[31:0] addr_14854_7;

Selector_2 s14854_7(wires_3713_6[2], addr_3713_6, addr_positional[59419:59416], addr_14854_7);

wire[31:0] addr_14855_7;

Selector_2 s14855_7(wires_3713_6[3], addr_3713_6, addr_positional[59423:59420], addr_14855_7);

wire[31:0] addr_14856_7;

Selector_2 s14856_7(wires_3714_6[0], addr_3714_6, addr_positional[59427:59424], addr_14856_7);

wire[31:0] addr_14857_7;

Selector_2 s14857_7(wires_3714_6[1], addr_3714_6, addr_positional[59431:59428], addr_14857_7);

wire[31:0] addr_14858_7;

Selector_2 s14858_7(wires_3714_6[2], addr_3714_6, addr_positional[59435:59432], addr_14858_7);

wire[31:0] addr_14859_7;

Selector_2 s14859_7(wires_3714_6[3], addr_3714_6, addr_positional[59439:59436], addr_14859_7);

wire[31:0] addr_14860_7;

Selector_2 s14860_7(wires_3715_6[0], addr_3715_6, addr_positional[59443:59440], addr_14860_7);

wire[31:0] addr_14861_7;

Selector_2 s14861_7(wires_3715_6[1], addr_3715_6, addr_positional[59447:59444], addr_14861_7);

wire[31:0] addr_14862_7;

Selector_2 s14862_7(wires_3715_6[2], addr_3715_6, addr_positional[59451:59448], addr_14862_7);

wire[31:0] addr_14863_7;

Selector_2 s14863_7(wires_3715_6[3], addr_3715_6, addr_positional[59455:59452], addr_14863_7);

wire[31:0] addr_14864_7;

Selector_2 s14864_7(wires_3716_6[0], addr_3716_6, addr_positional[59459:59456], addr_14864_7);

wire[31:0] addr_14865_7;

Selector_2 s14865_7(wires_3716_6[1], addr_3716_6, addr_positional[59463:59460], addr_14865_7);

wire[31:0] addr_14866_7;

Selector_2 s14866_7(wires_3716_6[2], addr_3716_6, addr_positional[59467:59464], addr_14866_7);

wire[31:0] addr_14867_7;

Selector_2 s14867_7(wires_3716_6[3], addr_3716_6, addr_positional[59471:59468], addr_14867_7);

wire[31:0] addr_14868_7;

Selector_2 s14868_7(wires_3717_6[0], addr_3717_6, addr_positional[59475:59472], addr_14868_7);

wire[31:0] addr_14869_7;

Selector_2 s14869_7(wires_3717_6[1], addr_3717_6, addr_positional[59479:59476], addr_14869_7);

wire[31:0] addr_14870_7;

Selector_2 s14870_7(wires_3717_6[2], addr_3717_6, addr_positional[59483:59480], addr_14870_7);

wire[31:0] addr_14871_7;

Selector_2 s14871_7(wires_3717_6[3], addr_3717_6, addr_positional[59487:59484], addr_14871_7);

wire[31:0] addr_14872_7;

Selector_2 s14872_7(wires_3718_6[0], addr_3718_6, addr_positional[59491:59488], addr_14872_7);

wire[31:0] addr_14873_7;

Selector_2 s14873_7(wires_3718_6[1], addr_3718_6, addr_positional[59495:59492], addr_14873_7);

wire[31:0] addr_14874_7;

Selector_2 s14874_7(wires_3718_6[2], addr_3718_6, addr_positional[59499:59496], addr_14874_7);

wire[31:0] addr_14875_7;

Selector_2 s14875_7(wires_3718_6[3], addr_3718_6, addr_positional[59503:59500], addr_14875_7);

wire[31:0] addr_14876_7;

Selector_2 s14876_7(wires_3719_6[0], addr_3719_6, addr_positional[59507:59504], addr_14876_7);

wire[31:0] addr_14877_7;

Selector_2 s14877_7(wires_3719_6[1], addr_3719_6, addr_positional[59511:59508], addr_14877_7);

wire[31:0] addr_14878_7;

Selector_2 s14878_7(wires_3719_6[2], addr_3719_6, addr_positional[59515:59512], addr_14878_7);

wire[31:0] addr_14879_7;

Selector_2 s14879_7(wires_3719_6[3], addr_3719_6, addr_positional[59519:59516], addr_14879_7);

wire[31:0] addr_14880_7;

Selector_2 s14880_7(wires_3720_6[0], addr_3720_6, addr_positional[59523:59520], addr_14880_7);

wire[31:0] addr_14881_7;

Selector_2 s14881_7(wires_3720_6[1], addr_3720_6, addr_positional[59527:59524], addr_14881_7);

wire[31:0] addr_14882_7;

Selector_2 s14882_7(wires_3720_6[2], addr_3720_6, addr_positional[59531:59528], addr_14882_7);

wire[31:0] addr_14883_7;

Selector_2 s14883_7(wires_3720_6[3], addr_3720_6, addr_positional[59535:59532], addr_14883_7);

wire[31:0] addr_14884_7;

Selector_2 s14884_7(wires_3721_6[0], addr_3721_6, addr_positional[59539:59536], addr_14884_7);

wire[31:0] addr_14885_7;

Selector_2 s14885_7(wires_3721_6[1], addr_3721_6, addr_positional[59543:59540], addr_14885_7);

wire[31:0] addr_14886_7;

Selector_2 s14886_7(wires_3721_6[2], addr_3721_6, addr_positional[59547:59544], addr_14886_7);

wire[31:0] addr_14887_7;

Selector_2 s14887_7(wires_3721_6[3], addr_3721_6, addr_positional[59551:59548], addr_14887_7);

wire[31:0] addr_14888_7;

Selector_2 s14888_7(wires_3722_6[0], addr_3722_6, addr_positional[59555:59552], addr_14888_7);

wire[31:0] addr_14889_7;

Selector_2 s14889_7(wires_3722_6[1], addr_3722_6, addr_positional[59559:59556], addr_14889_7);

wire[31:0] addr_14890_7;

Selector_2 s14890_7(wires_3722_6[2], addr_3722_6, addr_positional[59563:59560], addr_14890_7);

wire[31:0] addr_14891_7;

Selector_2 s14891_7(wires_3722_6[3], addr_3722_6, addr_positional[59567:59564], addr_14891_7);

wire[31:0] addr_14892_7;

Selector_2 s14892_7(wires_3723_6[0], addr_3723_6, addr_positional[59571:59568], addr_14892_7);

wire[31:0] addr_14893_7;

Selector_2 s14893_7(wires_3723_6[1], addr_3723_6, addr_positional[59575:59572], addr_14893_7);

wire[31:0] addr_14894_7;

Selector_2 s14894_7(wires_3723_6[2], addr_3723_6, addr_positional[59579:59576], addr_14894_7);

wire[31:0] addr_14895_7;

Selector_2 s14895_7(wires_3723_6[3], addr_3723_6, addr_positional[59583:59580], addr_14895_7);

wire[31:0] addr_14896_7;

Selector_2 s14896_7(wires_3724_6[0], addr_3724_6, addr_positional[59587:59584], addr_14896_7);

wire[31:0] addr_14897_7;

Selector_2 s14897_7(wires_3724_6[1], addr_3724_6, addr_positional[59591:59588], addr_14897_7);

wire[31:0] addr_14898_7;

Selector_2 s14898_7(wires_3724_6[2], addr_3724_6, addr_positional[59595:59592], addr_14898_7);

wire[31:0] addr_14899_7;

Selector_2 s14899_7(wires_3724_6[3], addr_3724_6, addr_positional[59599:59596], addr_14899_7);

wire[31:0] addr_14900_7;

Selector_2 s14900_7(wires_3725_6[0], addr_3725_6, addr_positional[59603:59600], addr_14900_7);

wire[31:0] addr_14901_7;

Selector_2 s14901_7(wires_3725_6[1], addr_3725_6, addr_positional[59607:59604], addr_14901_7);

wire[31:0] addr_14902_7;

Selector_2 s14902_7(wires_3725_6[2], addr_3725_6, addr_positional[59611:59608], addr_14902_7);

wire[31:0] addr_14903_7;

Selector_2 s14903_7(wires_3725_6[3], addr_3725_6, addr_positional[59615:59612], addr_14903_7);

wire[31:0] addr_14904_7;

Selector_2 s14904_7(wires_3726_6[0], addr_3726_6, addr_positional[59619:59616], addr_14904_7);

wire[31:0] addr_14905_7;

Selector_2 s14905_7(wires_3726_6[1], addr_3726_6, addr_positional[59623:59620], addr_14905_7);

wire[31:0] addr_14906_7;

Selector_2 s14906_7(wires_3726_6[2], addr_3726_6, addr_positional[59627:59624], addr_14906_7);

wire[31:0] addr_14907_7;

Selector_2 s14907_7(wires_3726_6[3], addr_3726_6, addr_positional[59631:59628], addr_14907_7);

wire[31:0] addr_14908_7;

Selector_2 s14908_7(wires_3727_6[0], addr_3727_6, addr_positional[59635:59632], addr_14908_7);

wire[31:0] addr_14909_7;

Selector_2 s14909_7(wires_3727_6[1], addr_3727_6, addr_positional[59639:59636], addr_14909_7);

wire[31:0] addr_14910_7;

Selector_2 s14910_7(wires_3727_6[2], addr_3727_6, addr_positional[59643:59640], addr_14910_7);

wire[31:0] addr_14911_7;

Selector_2 s14911_7(wires_3727_6[3], addr_3727_6, addr_positional[59647:59644], addr_14911_7);

wire[31:0] addr_14912_7;

Selector_2 s14912_7(wires_3728_6[0], addr_3728_6, addr_positional[59651:59648], addr_14912_7);

wire[31:0] addr_14913_7;

Selector_2 s14913_7(wires_3728_6[1], addr_3728_6, addr_positional[59655:59652], addr_14913_7);

wire[31:0] addr_14914_7;

Selector_2 s14914_7(wires_3728_6[2], addr_3728_6, addr_positional[59659:59656], addr_14914_7);

wire[31:0] addr_14915_7;

Selector_2 s14915_7(wires_3728_6[3], addr_3728_6, addr_positional[59663:59660], addr_14915_7);

wire[31:0] addr_14916_7;

Selector_2 s14916_7(wires_3729_6[0], addr_3729_6, addr_positional[59667:59664], addr_14916_7);

wire[31:0] addr_14917_7;

Selector_2 s14917_7(wires_3729_6[1], addr_3729_6, addr_positional[59671:59668], addr_14917_7);

wire[31:0] addr_14918_7;

Selector_2 s14918_7(wires_3729_6[2], addr_3729_6, addr_positional[59675:59672], addr_14918_7);

wire[31:0] addr_14919_7;

Selector_2 s14919_7(wires_3729_6[3], addr_3729_6, addr_positional[59679:59676], addr_14919_7);

wire[31:0] addr_14920_7;

Selector_2 s14920_7(wires_3730_6[0], addr_3730_6, addr_positional[59683:59680], addr_14920_7);

wire[31:0] addr_14921_7;

Selector_2 s14921_7(wires_3730_6[1], addr_3730_6, addr_positional[59687:59684], addr_14921_7);

wire[31:0] addr_14922_7;

Selector_2 s14922_7(wires_3730_6[2], addr_3730_6, addr_positional[59691:59688], addr_14922_7);

wire[31:0] addr_14923_7;

Selector_2 s14923_7(wires_3730_6[3], addr_3730_6, addr_positional[59695:59692], addr_14923_7);

wire[31:0] addr_14924_7;

Selector_2 s14924_7(wires_3731_6[0], addr_3731_6, addr_positional[59699:59696], addr_14924_7);

wire[31:0] addr_14925_7;

Selector_2 s14925_7(wires_3731_6[1], addr_3731_6, addr_positional[59703:59700], addr_14925_7);

wire[31:0] addr_14926_7;

Selector_2 s14926_7(wires_3731_6[2], addr_3731_6, addr_positional[59707:59704], addr_14926_7);

wire[31:0] addr_14927_7;

Selector_2 s14927_7(wires_3731_6[3], addr_3731_6, addr_positional[59711:59708], addr_14927_7);

wire[31:0] addr_14928_7;

Selector_2 s14928_7(wires_3732_6[0], addr_3732_6, addr_positional[59715:59712], addr_14928_7);

wire[31:0] addr_14929_7;

Selector_2 s14929_7(wires_3732_6[1], addr_3732_6, addr_positional[59719:59716], addr_14929_7);

wire[31:0] addr_14930_7;

Selector_2 s14930_7(wires_3732_6[2], addr_3732_6, addr_positional[59723:59720], addr_14930_7);

wire[31:0] addr_14931_7;

Selector_2 s14931_7(wires_3732_6[3], addr_3732_6, addr_positional[59727:59724], addr_14931_7);

wire[31:0] addr_14932_7;

Selector_2 s14932_7(wires_3733_6[0], addr_3733_6, addr_positional[59731:59728], addr_14932_7);

wire[31:0] addr_14933_7;

Selector_2 s14933_7(wires_3733_6[1], addr_3733_6, addr_positional[59735:59732], addr_14933_7);

wire[31:0] addr_14934_7;

Selector_2 s14934_7(wires_3733_6[2], addr_3733_6, addr_positional[59739:59736], addr_14934_7);

wire[31:0] addr_14935_7;

Selector_2 s14935_7(wires_3733_6[3], addr_3733_6, addr_positional[59743:59740], addr_14935_7);

wire[31:0] addr_14936_7;

Selector_2 s14936_7(wires_3734_6[0], addr_3734_6, addr_positional[59747:59744], addr_14936_7);

wire[31:0] addr_14937_7;

Selector_2 s14937_7(wires_3734_6[1], addr_3734_6, addr_positional[59751:59748], addr_14937_7);

wire[31:0] addr_14938_7;

Selector_2 s14938_7(wires_3734_6[2], addr_3734_6, addr_positional[59755:59752], addr_14938_7);

wire[31:0] addr_14939_7;

Selector_2 s14939_7(wires_3734_6[3], addr_3734_6, addr_positional[59759:59756], addr_14939_7);

wire[31:0] addr_14940_7;

Selector_2 s14940_7(wires_3735_6[0], addr_3735_6, addr_positional[59763:59760], addr_14940_7);

wire[31:0] addr_14941_7;

Selector_2 s14941_7(wires_3735_6[1], addr_3735_6, addr_positional[59767:59764], addr_14941_7);

wire[31:0] addr_14942_7;

Selector_2 s14942_7(wires_3735_6[2], addr_3735_6, addr_positional[59771:59768], addr_14942_7);

wire[31:0] addr_14943_7;

Selector_2 s14943_7(wires_3735_6[3], addr_3735_6, addr_positional[59775:59772], addr_14943_7);

wire[31:0] addr_14944_7;

Selector_2 s14944_7(wires_3736_6[0], addr_3736_6, addr_positional[59779:59776], addr_14944_7);

wire[31:0] addr_14945_7;

Selector_2 s14945_7(wires_3736_6[1], addr_3736_6, addr_positional[59783:59780], addr_14945_7);

wire[31:0] addr_14946_7;

Selector_2 s14946_7(wires_3736_6[2], addr_3736_6, addr_positional[59787:59784], addr_14946_7);

wire[31:0] addr_14947_7;

Selector_2 s14947_7(wires_3736_6[3], addr_3736_6, addr_positional[59791:59788], addr_14947_7);

wire[31:0] addr_14948_7;

Selector_2 s14948_7(wires_3737_6[0], addr_3737_6, addr_positional[59795:59792], addr_14948_7);

wire[31:0] addr_14949_7;

Selector_2 s14949_7(wires_3737_6[1], addr_3737_6, addr_positional[59799:59796], addr_14949_7);

wire[31:0] addr_14950_7;

Selector_2 s14950_7(wires_3737_6[2], addr_3737_6, addr_positional[59803:59800], addr_14950_7);

wire[31:0] addr_14951_7;

Selector_2 s14951_7(wires_3737_6[3], addr_3737_6, addr_positional[59807:59804], addr_14951_7);

wire[31:0] addr_14952_7;

Selector_2 s14952_7(wires_3738_6[0], addr_3738_6, addr_positional[59811:59808], addr_14952_7);

wire[31:0] addr_14953_7;

Selector_2 s14953_7(wires_3738_6[1], addr_3738_6, addr_positional[59815:59812], addr_14953_7);

wire[31:0] addr_14954_7;

Selector_2 s14954_7(wires_3738_6[2], addr_3738_6, addr_positional[59819:59816], addr_14954_7);

wire[31:0] addr_14955_7;

Selector_2 s14955_7(wires_3738_6[3], addr_3738_6, addr_positional[59823:59820], addr_14955_7);

wire[31:0] addr_14956_7;

Selector_2 s14956_7(wires_3739_6[0], addr_3739_6, addr_positional[59827:59824], addr_14956_7);

wire[31:0] addr_14957_7;

Selector_2 s14957_7(wires_3739_6[1], addr_3739_6, addr_positional[59831:59828], addr_14957_7);

wire[31:0] addr_14958_7;

Selector_2 s14958_7(wires_3739_6[2], addr_3739_6, addr_positional[59835:59832], addr_14958_7);

wire[31:0] addr_14959_7;

Selector_2 s14959_7(wires_3739_6[3], addr_3739_6, addr_positional[59839:59836], addr_14959_7);

wire[31:0] addr_14960_7;

Selector_2 s14960_7(wires_3740_6[0], addr_3740_6, addr_positional[59843:59840], addr_14960_7);

wire[31:0] addr_14961_7;

Selector_2 s14961_7(wires_3740_6[1], addr_3740_6, addr_positional[59847:59844], addr_14961_7);

wire[31:0] addr_14962_7;

Selector_2 s14962_7(wires_3740_6[2], addr_3740_6, addr_positional[59851:59848], addr_14962_7);

wire[31:0] addr_14963_7;

Selector_2 s14963_7(wires_3740_6[3], addr_3740_6, addr_positional[59855:59852], addr_14963_7);

wire[31:0] addr_14964_7;

Selector_2 s14964_7(wires_3741_6[0], addr_3741_6, addr_positional[59859:59856], addr_14964_7);

wire[31:0] addr_14965_7;

Selector_2 s14965_7(wires_3741_6[1], addr_3741_6, addr_positional[59863:59860], addr_14965_7);

wire[31:0] addr_14966_7;

Selector_2 s14966_7(wires_3741_6[2], addr_3741_6, addr_positional[59867:59864], addr_14966_7);

wire[31:0] addr_14967_7;

Selector_2 s14967_7(wires_3741_6[3], addr_3741_6, addr_positional[59871:59868], addr_14967_7);

wire[31:0] addr_14968_7;

Selector_2 s14968_7(wires_3742_6[0], addr_3742_6, addr_positional[59875:59872], addr_14968_7);

wire[31:0] addr_14969_7;

Selector_2 s14969_7(wires_3742_6[1], addr_3742_6, addr_positional[59879:59876], addr_14969_7);

wire[31:0] addr_14970_7;

Selector_2 s14970_7(wires_3742_6[2], addr_3742_6, addr_positional[59883:59880], addr_14970_7);

wire[31:0] addr_14971_7;

Selector_2 s14971_7(wires_3742_6[3], addr_3742_6, addr_positional[59887:59884], addr_14971_7);

wire[31:0] addr_14972_7;

Selector_2 s14972_7(wires_3743_6[0], addr_3743_6, addr_positional[59891:59888], addr_14972_7);

wire[31:0] addr_14973_7;

Selector_2 s14973_7(wires_3743_6[1], addr_3743_6, addr_positional[59895:59892], addr_14973_7);

wire[31:0] addr_14974_7;

Selector_2 s14974_7(wires_3743_6[2], addr_3743_6, addr_positional[59899:59896], addr_14974_7);

wire[31:0] addr_14975_7;

Selector_2 s14975_7(wires_3743_6[3], addr_3743_6, addr_positional[59903:59900], addr_14975_7);

wire[31:0] addr_14976_7;

Selector_2 s14976_7(wires_3744_6[0], addr_3744_6, addr_positional[59907:59904], addr_14976_7);

wire[31:0] addr_14977_7;

Selector_2 s14977_7(wires_3744_6[1], addr_3744_6, addr_positional[59911:59908], addr_14977_7);

wire[31:0] addr_14978_7;

Selector_2 s14978_7(wires_3744_6[2], addr_3744_6, addr_positional[59915:59912], addr_14978_7);

wire[31:0] addr_14979_7;

Selector_2 s14979_7(wires_3744_6[3], addr_3744_6, addr_positional[59919:59916], addr_14979_7);

wire[31:0] addr_14980_7;

Selector_2 s14980_7(wires_3745_6[0], addr_3745_6, addr_positional[59923:59920], addr_14980_7);

wire[31:0] addr_14981_7;

Selector_2 s14981_7(wires_3745_6[1], addr_3745_6, addr_positional[59927:59924], addr_14981_7);

wire[31:0] addr_14982_7;

Selector_2 s14982_7(wires_3745_6[2], addr_3745_6, addr_positional[59931:59928], addr_14982_7);

wire[31:0] addr_14983_7;

Selector_2 s14983_7(wires_3745_6[3], addr_3745_6, addr_positional[59935:59932], addr_14983_7);

wire[31:0] addr_14984_7;

Selector_2 s14984_7(wires_3746_6[0], addr_3746_6, addr_positional[59939:59936], addr_14984_7);

wire[31:0] addr_14985_7;

Selector_2 s14985_7(wires_3746_6[1], addr_3746_6, addr_positional[59943:59940], addr_14985_7);

wire[31:0] addr_14986_7;

Selector_2 s14986_7(wires_3746_6[2], addr_3746_6, addr_positional[59947:59944], addr_14986_7);

wire[31:0] addr_14987_7;

Selector_2 s14987_7(wires_3746_6[3], addr_3746_6, addr_positional[59951:59948], addr_14987_7);

wire[31:0] addr_14988_7;

Selector_2 s14988_7(wires_3747_6[0], addr_3747_6, addr_positional[59955:59952], addr_14988_7);

wire[31:0] addr_14989_7;

Selector_2 s14989_7(wires_3747_6[1], addr_3747_6, addr_positional[59959:59956], addr_14989_7);

wire[31:0] addr_14990_7;

Selector_2 s14990_7(wires_3747_6[2], addr_3747_6, addr_positional[59963:59960], addr_14990_7);

wire[31:0] addr_14991_7;

Selector_2 s14991_7(wires_3747_6[3], addr_3747_6, addr_positional[59967:59964], addr_14991_7);

wire[31:0] addr_14992_7;

Selector_2 s14992_7(wires_3748_6[0], addr_3748_6, addr_positional[59971:59968], addr_14992_7);

wire[31:0] addr_14993_7;

Selector_2 s14993_7(wires_3748_6[1], addr_3748_6, addr_positional[59975:59972], addr_14993_7);

wire[31:0] addr_14994_7;

Selector_2 s14994_7(wires_3748_6[2], addr_3748_6, addr_positional[59979:59976], addr_14994_7);

wire[31:0] addr_14995_7;

Selector_2 s14995_7(wires_3748_6[3], addr_3748_6, addr_positional[59983:59980], addr_14995_7);

wire[31:0] addr_14996_7;

Selector_2 s14996_7(wires_3749_6[0], addr_3749_6, addr_positional[59987:59984], addr_14996_7);

wire[31:0] addr_14997_7;

Selector_2 s14997_7(wires_3749_6[1], addr_3749_6, addr_positional[59991:59988], addr_14997_7);

wire[31:0] addr_14998_7;

Selector_2 s14998_7(wires_3749_6[2], addr_3749_6, addr_positional[59995:59992], addr_14998_7);

wire[31:0] addr_14999_7;

Selector_2 s14999_7(wires_3749_6[3], addr_3749_6, addr_positional[59999:59996], addr_14999_7);

wire[31:0] addr_15000_7;

Selector_2 s15000_7(wires_3750_6[0], addr_3750_6, addr_positional[60003:60000], addr_15000_7);

wire[31:0] addr_15001_7;

Selector_2 s15001_7(wires_3750_6[1], addr_3750_6, addr_positional[60007:60004], addr_15001_7);

wire[31:0] addr_15002_7;

Selector_2 s15002_7(wires_3750_6[2], addr_3750_6, addr_positional[60011:60008], addr_15002_7);

wire[31:0] addr_15003_7;

Selector_2 s15003_7(wires_3750_6[3], addr_3750_6, addr_positional[60015:60012], addr_15003_7);

wire[31:0] addr_15004_7;

Selector_2 s15004_7(wires_3751_6[0], addr_3751_6, addr_positional[60019:60016], addr_15004_7);

wire[31:0] addr_15005_7;

Selector_2 s15005_7(wires_3751_6[1], addr_3751_6, addr_positional[60023:60020], addr_15005_7);

wire[31:0] addr_15006_7;

Selector_2 s15006_7(wires_3751_6[2], addr_3751_6, addr_positional[60027:60024], addr_15006_7);

wire[31:0] addr_15007_7;

Selector_2 s15007_7(wires_3751_6[3], addr_3751_6, addr_positional[60031:60028], addr_15007_7);

wire[31:0] addr_15008_7;

Selector_2 s15008_7(wires_3752_6[0], addr_3752_6, addr_positional[60035:60032], addr_15008_7);

wire[31:0] addr_15009_7;

Selector_2 s15009_7(wires_3752_6[1], addr_3752_6, addr_positional[60039:60036], addr_15009_7);

wire[31:0] addr_15010_7;

Selector_2 s15010_7(wires_3752_6[2], addr_3752_6, addr_positional[60043:60040], addr_15010_7);

wire[31:0] addr_15011_7;

Selector_2 s15011_7(wires_3752_6[3], addr_3752_6, addr_positional[60047:60044], addr_15011_7);

wire[31:0] addr_15012_7;

Selector_2 s15012_7(wires_3753_6[0], addr_3753_6, addr_positional[60051:60048], addr_15012_7);

wire[31:0] addr_15013_7;

Selector_2 s15013_7(wires_3753_6[1], addr_3753_6, addr_positional[60055:60052], addr_15013_7);

wire[31:0] addr_15014_7;

Selector_2 s15014_7(wires_3753_6[2], addr_3753_6, addr_positional[60059:60056], addr_15014_7);

wire[31:0] addr_15015_7;

Selector_2 s15015_7(wires_3753_6[3], addr_3753_6, addr_positional[60063:60060], addr_15015_7);

wire[31:0] addr_15016_7;

Selector_2 s15016_7(wires_3754_6[0], addr_3754_6, addr_positional[60067:60064], addr_15016_7);

wire[31:0] addr_15017_7;

Selector_2 s15017_7(wires_3754_6[1], addr_3754_6, addr_positional[60071:60068], addr_15017_7);

wire[31:0] addr_15018_7;

Selector_2 s15018_7(wires_3754_6[2], addr_3754_6, addr_positional[60075:60072], addr_15018_7);

wire[31:0] addr_15019_7;

Selector_2 s15019_7(wires_3754_6[3], addr_3754_6, addr_positional[60079:60076], addr_15019_7);

wire[31:0] addr_15020_7;

Selector_2 s15020_7(wires_3755_6[0], addr_3755_6, addr_positional[60083:60080], addr_15020_7);

wire[31:0] addr_15021_7;

Selector_2 s15021_7(wires_3755_6[1], addr_3755_6, addr_positional[60087:60084], addr_15021_7);

wire[31:0] addr_15022_7;

Selector_2 s15022_7(wires_3755_6[2], addr_3755_6, addr_positional[60091:60088], addr_15022_7);

wire[31:0] addr_15023_7;

Selector_2 s15023_7(wires_3755_6[3], addr_3755_6, addr_positional[60095:60092], addr_15023_7);

wire[31:0] addr_15024_7;

Selector_2 s15024_7(wires_3756_6[0], addr_3756_6, addr_positional[60099:60096], addr_15024_7);

wire[31:0] addr_15025_7;

Selector_2 s15025_7(wires_3756_6[1], addr_3756_6, addr_positional[60103:60100], addr_15025_7);

wire[31:0] addr_15026_7;

Selector_2 s15026_7(wires_3756_6[2], addr_3756_6, addr_positional[60107:60104], addr_15026_7);

wire[31:0] addr_15027_7;

Selector_2 s15027_7(wires_3756_6[3], addr_3756_6, addr_positional[60111:60108], addr_15027_7);

wire[31:0] addr_15028_7;

Selector_2 s15028_7(wires_3757_6[0], addr_3757_6, addr_positional[60115:60112], addr_15028_7);

wire[31:0] addr_15029_7;

Selector_2 s15029_7(wires_3757_6[1], addr_3757_6, addr_positional[60119:60116], addr_15029_7);

wire[31:0] addr_15030_7;

Selector_2 s15030_7(wires_3757_6[2], addr_3757_6, addr_positional[60123:60120], addr_15030_7);

wire[31:0] addr_15031_7;

Selector_2 s15031_7(wires_3757_6[3], addr_3757_6, addr_positional[60127:60124], addr_15031_7);

wire[31:0] addr_15032_7;

Selector_2 s15032_7(wires_3758_6[0], addr_3758_6, addr_positional[60131:60128], addr_15032_7);

wire[31:0] addr_15033_7;

Selector_2 s15033_7(wires_3758_6[1], addr_3758_6, addr_positional[60135:60132], addr_15033_7);

wire[31:0] addr_15034_7;

Selector_2 s15034_7(wires_3758_6[2], addr_3758_6, addr_positional[60139:60136], addr_15034_7);

wire[31:0] addr_15035_7;

Selector_2 s15035_7(wires_3758_6[3], addr_3758_6, addr_positional[60143:60140], addr_15035_7);

wire[31:0] addr_15036_7;

Selector_2 s15036_7(wires_3759_6[0], addr_3759_6, addr_positional[60147:60144], addr_15036_7);

wire[31:0] addr_15037_7;

Selector_2 s15037_7(wires_3759_6[1], addr_3759_6, addr_positional[60151:60148], addr_15037_7);

wire[31:0] addr_15038_7;

Selector_2 s15038_7(wires_3759_6[2], addr_3759_6, addr_positional[60155:60152], addr_15038_7);

wire[31:0] addr_15039_7;

Selector_2 s15039_7(wires_3759_6[3], addr_3759_6, addr_positional[60159:60156], addr_15039_7);

wire[31:0] addr_15040_7;

Selector_2 s15040_7(wires_3760_6[0], addr_3760_6, addr_positional[60163:60160], addr_15040_7);

wire[31:0] addr_15041_7;

Selector_2 s15041_7(wires_3760_6[1], addr_3760_6, addr_positional[60167:60164], addr_15041_7);

wire[31:0] addr_15042_7;

Selector_2 s15042_7(wires_3760_6[2], addr_3760_6, addr_positional[60171:60168], addr_15042_7);

wire[31:0] addr_15043_7;

Selector_2 s15043_7(wires_3760_6[3], addr_3760_6, addr_positional[60175:60172], addr_15043_7);

wire[31:0] addr_15044_7;

Selector_2 s15044_7(wires_3761_6[0], addr_3761_6, addr_positional[60179:60176], addr_15044_7);

wire[31:0] addr_15045_7;

Selector_2 s15045_7(wires_3761_6[1], addr_3761_6, addr_positional[60183:60180], addr_15045_7);

wire[31:0] addr_15046_7;

Selector_2 s15046_7(wires_3761_6[2], addr_3761_6, addr_positional[60187:60184], addr_15046_7);

wire[31:0] addr_15047_7;

Selector_2 s15047_7(wires_3761_6[3], addr_3761_6, addr_positional[60191:60188], addr_15047_7);

wire[31:0] addr_15048_7;

Selector_2 s15048_7(wires_3762_6[0], addr_3762_6, addr_positional[60195:60192], addr_15048_7);

wire[31:0] addr_15049_7;

Selector_2 s15049_7(wires_3762_6[1], addr_3762_6, addr_positional[60199:60196], addr_15049_7);

wire[31:0] addr_15050_7;

Selector_2 s15050_7(wires_3762_6[2], addr_3762_6, addr_positional[60203:60200], addr_15050_7);

wire[31:0] addr_15051_7;

Selector_2 s15051_7(wires_3762_6[3], addr_3762_6, addr_positional[60207:60204], addr_15051_7);

wire[31:0] addr_15052_7;

Selector_2 s15052_7(wires_3763_6[0], addr_3763_6, addr_positional[60211:60208], addr_15052_7);

wire[31:0] addr_15053_7;

Selector_2 s15053_7(wires_3763_6[1], addr_3763_6, addr_positional[60215:60212], addr_15053_7);

wire[31:0] addr_15054_7;

Selector_2 s15054_7(wires_3763_6[2], addr_3763_6, addr_positional[60219:60216], addr_15054_7);

wire[31:0] addr_15055_7;

Selector_2 s15055_7(wires_3763_6[3], addr_3763_6, addr_positional[60223:60220], addr_15055_7);

wire[31:0] addr_15056_7;

Selector_2 s15056_7(wires_3764_6[0], addr_3764_6, addr_positional[60227:60224], addr_15056_7);

wire[31:0] addr_15057_7;

Selector_2 s15057_7(wires_3764_6[1], addr_3764_6, addr_positional[60231:60228], addr_15057_7);

wire[31:0] addr_15058_7;

Selector_2 s15058_7(wires_3764_6[2], addr_3764_6, addr_positional[60235:60232], addr_15058_7);

wire[31:0] addr_15059_7;

Selector_2 s15059_7(wires_3764_6[3], addr_3764_6, addr_positional[60239:60236], addr_15059_7);

wire[31:0] addr_15060_7;

Selector_2 s15060_7(wires_3765_6[0], addr_3765_6, addr_positional[60243:60240], addr_15060_7);

wire[31:0] addr_15061_7;

Selector_2 s15061_7(wires_3765_6[1], addr_3765_6, addr_positional[60247:60244], addr_15061_7);

wire[31:0] addr_15062_7;

Selector_2 s15062_7(wires_3765_6[2], addr_3765_6, addr_positional[60251:60248], addr_15062_7);

wire[31:0] addr_15063_7;

Selector_2 s15063_7(wires_3765_6[3], addr_3765_6, addr_positional[60255:60252], addr_15063_7);

wire[31:0] addr_15064_7;

Selector_2 s15064_7(wires_3766_6[0], addr_3766_6, addr_positional[60259:60256], addr_15064_7);

wire[31:0] addr_15065_7;

Selector_2 s15065_7(wires_3766_6[1], addr_3766_6, addr_positional[60263:60260], addr_15065_7);

wire[31:0] addr_15066_7;

Selector_2 s15066_7(wires_3766_6[2], addr_3766_6, addr_positional[60267:60264], addr_15066_7);

wire[31:0] addr_15067_7;

Selector_2 s15067_7(wires_3766_6[3], addr_3766_6, addr_positional[60271:60268], addr_15067_7);

wire[31:0] addr_15068_7;

Selector_2 s15068_7(wires_3767_6[0], addr_3767_6, addr_positional[60275:60272], addr_15068_7);

wire[31:0] addr_15069_7;

Selector_2 s15069_7(wires_3767_6[1], addr_3767_6, addr_positional[60279:60276], addr_15069_7);

wire[31:0] addr_15070_7;

Selector_2 s15070_7(wires_3767_6[2], addr_3767_6, addr_positional[60283:60280], addr_15070_7);

wire[31:0] addr_15071_7;

Selector_2 s15071_7(wires_3767_6[3], addr_3767_6, addr_positional[60287:60284], addr_15071_7);

wire[31:0] addr_15072_7;

Selector_2 s15072_7(wires_3768_6[0], addr_3768_6, addr_positional[60291:60288], addr_15072_7);

wire[31:0] addr_15073_7;

Selector_2 s15073_7(wires_3768_6[1], addr_3768_6, addr_positional[60295:60292], addr_15073_7);

wire[31:0] addr_15074_7;

Selector_2 s15074_7(wires_3768_6[2], addr_3768_6, addr_positional[60299:60296], addr_15074_7);

wire[31:0] addr_15075_7;

Selector_2 s15075_7(wires_3768_6[3], addr_3768_6, addr_positional[60303:60300], addr_15075_7);

wire[31:0] addr_15076_7;

Selector_2 s15076_7(wires_3769_6[0], addr_3769_6, addr_positional[60307:60304], addr_15076_7);

wire[31:0] addr_15077_7;

Selector_2 s15077_7(wires_3769_6[1], addr_3769_6, addr_positional[60311:60308], addr_15077_7);

wire[31:0] addr_15078_7;

Selector_2 s15078_7(wires_3769_6[2], addr_3769_6, addr_positional[60315:60312], addr_15078_7);

wire[31:0] addr_15079_7;

Selector_2 s15079_7(wires_3769_6[3], addr_3769_6, addr_positional[60319:60316], addr_15079_7);

wire[31:0] addr_15080_7;

Selector_2 s15080_7(wires_3770_6[0], addr_3770_6, addr_positional[60323:60320], addr_15080_7);

wire[31:0] addr_15081_7;

Selector_2 s15081_7(wires_3770_6[1], addr_3770_6, addr_positional[60327:60324], addr_15081_7);

wire[31:0] addr_15082_7;

Selector_2 s15082_7(wires_3770_6[2], addr_3770_6, addr_positional[60331:60328], addr_15082_7);

wire[31:0] addr_15083_7;

Selector_2 s15083_7(wires_3770_6[3], addr_3770_6, addr_positional[60335:60332], addr_15083_7);

wire[31:0] addr_15084_7;

Selector_2 s15084_7(wires_3771_6[0], addr_3771_6, addr_positional[60339:60336], addr_15084_7);

wire[31:0] addr_15085_7;

Selector_2 s15085_7(wires_3771_6[1], addr_3771_6, addr_positional[60343:60340], addr_15085_7);

wire[31:0] addr_15086_7;

Selector_2 s15086_7(wires_3771_6[2], addr_3771_6, addr_positional[60347:60344], addr_15086_7);

wire[31:0] addr_15087_7;

Selector_2 s15087_7(wires_3771_6[3], addr_3771_6, addr_positional[60351:60348], addr_15087_7);

wire[31:0] addr_15088_7;

Selector_2 s15088_7(wires_3772_6[0], addr_3772_6, addr_positional[60355:60352], addr_15088_7);

wire[31:0] addr_15089_7;

Selector_2 s15089_7(wires_3772_6[1], addr_3772_6, addr_positional[60359:60356], addr_15089_7);

wire[31:0] addr_15090_7;

Selector_2 s15090_7(wires_3772_6[2], addr_3772_6, addr_positional[60363:60360], addr_15090_7);

wire[31:0] addr_15091_7;

Selector_2 s15091_7(wires_3772_6[3], addr_3772_6, addr_positional[60367:60364], addr_15091_7);

wire[31:0] addr_15092_7;

Selector_2 s15092_7(wires_3773_6[0], addr_3773_6, addr_positional[60371:60368], addr_15092_7);

wire[31:0] addr_15093_7;

Selector_2 s15093_7(wires_3773_6[1], addr_3773_6, addr_positional[60375:60372], addr_15093_7);

wire[31:0] addr_15094_7;

Selector_2 s15094_7(wires_3773_6[2], addr_3773_6, addr_positional[60379:60376], addr_15094_7);

wire[31:0] addr_15095_7;

Selector_2 s15095_7(wires_3773_6[3], addr_3773_6, addr_positional[60383:60380], addr_15095_7);

wire[31:0] addr_15096_7;

Selector_2 s15096_7(wires_3774_6[0], addr_3774_6, addr_positional[60387:60384], addr_15096_7);

wire[31:0] addr_15097_7;

Selector_2 s15097_7(wires_3774_6[1], addr_3774_6, addr_positional[60391:60388], addr_15097_7);

wire[31:0] addr_15098_7;

Selector_2 s15098_7(wires_3774_6[2], addr_3774_6, addr_positional[60395:60392], addr_15098_7);

wire[31:0] addr_15099_7;

Selector_2 s15099_7(wires_3774_6[3], addr_3774_6, addr_positional[60399:60396], addr_15099_7);

wire[31:0] addr_15100_7;

Selector_2 s15100_7(wires_3775_6[0], addr_3775_6, addr_positional[60403:60400], addr_15100_7);

wire[31:0] addr_15101_7;

Selector_2 s15101_7(wires_3775_6[1], addr_3775_6, addr_positional[60407:60404], addr_15101_7);

wire[31:0] addr_15102_7;

Selector_2 s15102_7(wires_3775_6[2], addr_3775_6, addr_positional[60411:60408], addr_15102_7);

wire[31:0] addr_15103_7;

Selector_2 s15103_7(wires_3775_6[3], addr_3775_6, addr_positional[60415:60412], addr_15103_7);

wire[31:0] addr_15104_7;

Selector_2 s15104_7(wires_3776_6[0], addr_3776_6, addr_positional[60419:60416], addr_15104_7);

wire[31:0] addr_15105_7;

Selector_2 s15105_7(wires_3776_6[1], addr_3776_6, addr_positional[60423:60420], addr_15105_7);

wire[31:0] addr_15106_7;

Selector_2 s15106_7(wires_3776_6[2], addr_3776_6, addr_positional[60427:60424], addr_15106_7);

wire[31:0] addr_15107_7;

Selector_2 s15107_7(wires_3776_6[3], addr_3776_6, addr_positional[60431:60428], addr_15107_7);

wire[31:0] addr_15108_7;

Selector_2 s15108_7(wires_3777_6[0], addr_3777_6, addr_positional[60435:60432], addr_15108_7);

wire[31:0] addr_15109_7;

Selector_2 s15109_7(wires_3777_6[1], addr_3777_6, addr_positional[60439:60436], addr_15109_7);

wire[31:0] addr_15110_7;

Selector_2 s15110_7(wires_3777_6[2], addr_3777_6, addr_positional[60443:60440], addr_15110_7);

wire[31:0] addr_15111_7;

Selector_2 s15111_7(wires_3777_6[3], addr_3777_6, addr_positional[60447:60444], addr_15111_7);

wire[31:0] addr_15112_7;

Selector_2 s15112_7(wires_3778_6[0], addr_3778_6, addr_positional[60451:60448], addr_15112_7);

wire[31:0] addr_15113_7;

Selector_2 s15113_7(wires_3778_6[1], addr_3778_6, addr_positional[60455:60452], addr_15113_7);

wire[31:0] addr_15114_7;

Selector_2 s15114_7(wires_3778_6[2], addr_3778_6, addr_positional[60459:60456], addr_15114_7);

wire[31:0] addr_15115_7;

Selector_2 s15115_7(wires_3778_6[3], addr_3778_6, addr_positional[60463:60460], addr_15115_7);

wire[31:0] addr_15116_7;

Selector_2 s15116_7(wires_3779_6[0], addr_3779_6, addr_positional[60467:60464], addr_15116_7);

wire[31:0] addr_15117_7;

Selector_2 s15117_7(wires_3779_6[1], addr_3779_6, addr_positional[60471:60468], addr_15117_7);

wire[31:0] addr_15118_7;

Selector_2 s15118_7(wires_3779_6[2], addr_3779_6, addr_positional[60475:60472], addr_15118_7);

wire[31:0] addr_15119_7;

Selector_2 s15119_7(wires_3779_6[3], addr_3779_6, addr_positional[60479:60476], addr_15119_7);

wire[31:0] addr_15120_7;

Selector_2 s15120_7(wires_3780_6[0], addr_3780_6, addr_positional[60483:60480], addr_15120_7);

wire[31:0] addr_15121_7;

Selector_2 s15121_7(wires_3780_6[1], addr_3780_6, addr_positional[60487:60484], addr_15121_7);

wire[31:0] addr_15122_7;

Selector_2 s15122_7(wires_3780_6[2], addr_3780_6, addr_positional[60491:60488], addr_15122_7);

wire[31:0] addr_15123_7;

Selector_2 s15123_7(wires_3780_6[3], addr_3780_6, addr_positional[60495:60492], addr_15123_7);

wire[31:0] addr_15124_7;

Selector_2 s15124_7(wires_3781_6[0], addr_3781_6, addr_positional[60499:60496], addr_15124_7);

wire[31:0] addr_15125_7;

Selector_2 s15125_7(wires_3781_6[1], addr_3781_6, addr_positional[60503:60500], addr_15125_7);

wire[31:0] addr_15126_7;

Selector_2 s15126_7(wires_3781_6[2], addr_3781_6, addr_positional[60507:60504], addr_15126_7);

wire[31:0] addr_15127_7;

Selector_2 s15127_7(wires_3781_6[3], addr_3781_6, addr_positional[60511:60508], addr_15127_7);

wire[31:0] addr_15128_7;

Selector_2 s15128_7(wires_3782_6[0], addr_3782_6, addr_positional[60515:60512], addr_15128_7);

wire[31:0] addr_15129_7;

Selector_2 s15129_7(wires_3782_6[1], addr_3782_6, addr_positional[60519:60516], addr_15129_7);

wire[31:0] addr_15130_7;

Selector_2 s15130_7(wires_3782_6[2], addr_3782_6, addr_positional[60523:60520], addr_15130_7);

wire[31:0] addr_15131_7;

Selector_2 s15131_7(wires_3782_6[3], addr_3782_6, addr_positional[60527:60524], addr_15131_7);

wire[31:0] addr_15132_7;

Selector_2 s15132_7(wires_3783_6[0], addr_3783_6, addr_positional[60531:60528], addr_15132_7);

wire[31:0] addr_15133_7;

Selector_2 s15133_7(wires_3783_6[1], addr_3783_6, addr_positional[60535:60532], addr_15133_7);

wire[31:0] addr_15134_7;

Selector_2 s15134_7(wires_3783_6[2], addr_3783_6, addr_positional[60539:60536], addr_15134_7);

wire[31:0] addr_15135_7;

Selector_2 s15135_7(wires_3783_6[3], addr_3783_6, addr_positional[60543:60540], addr_15135_7);

wire[31:0] addr_15136_7;

Selector_2 s15136_7(wires_3784_6[0], addr_3784_6, addr_positional[60547:60544], addr_15136_7);

wire[31:0] addr_15137_7;

Selector_2 s15137_7(wires_3784_6[1], addr_3784_6, addr_positional[60551:60548], addr_15137_7);

wire[31:0] addr_15138_7;

Selector_2 s15138_7(wires_3784_6[2], addr_3784_6, addr_positional[60555:60552], addr_15138_7);

wire[31:0] addr_15139_7;

Selector_2 s15139_7(wires_3784_6[3], addr_3784_6, addr_positional[60559:60556], addr_15139_7);

wire[31:0] addr_15140_7;

Selector_2 s15140_7(wires_3785_6[0], addr_3785_6, addr_positional[60563:60560], addr_15140_7);

wire[31:0] addr_15141_7;

Selector_2 s15141_7(wires_3785_6[1], addr_3785_6, addr_positional[60567:60564], addr_15141_7);

wire[31:0] addr_15142_7;

Selector_2 s15142_7(wires_3785_6[2], addr_3785_6, addr_positional[60571:60568], addr_15142_7);

wire[31:0] addr_15143_7;

Selector_2 s15143_7(wires_3785_6[3], addr_3785_6, addr_positional[60575:60572], addr_15143_7);

wire[31:0] addr_15144_7;

Selector_2 s15144_7(wires_3786_6[0], addr_3786_6, addr_positional[60579:60576], addr_15144_7);

wire[31:0] addr_15145_7;

Selector_2 s15145_7(wires_3786_6[1], addr_3786_6, addr_positional[60583:60580], addr_15145_7);

wire[31:0] addr_15146_7;

Selector_2 s15146_7(wires_3786_6[2], addr_3786_6, addr_positional[60587:60584], addr_15146_7);

wire[31:0] addr_15147_7;

Selector_2 s15147_7(wires_3786_6[3], addr_3786_6, addr_positional[60591:60588], addr_15147_7);

wire[31:0] addr_15148_7;

Selector_2 s15148_7(wires_3787_6[0], addr_3787_6, addr_positional[60595:60592], addr_15148_7);

wire[31:0] addr_15149_7;

Selector_2 s15149_7(wires_3787_6[1], addr_3787_6, addr_positional[60599:60596], addr_15149_7);

wire[31:0] addr_15150_7;

Selector_2 s15150_7(wires_3787_6[2], addr_3787_6, addr_positional[60603:60600], addr_15150_7);

wire[31:0] addr_15151_7;

Selector_2 s15151_7(wires_3787_6[3], addr_3787_6, addr_positional[60607:60604], addr_15151_7);

wire[31:0] addr_15152_7;

Selector_2 s15152_7(wires_3788_6[0], addr_3788_6, addr_positional[60611:60608], addr_15152_7);

wire[31:0] addr_15153_7;

Selector_2 s15153_7(wires_3788_6[1], addr_3788_6, addr_positional[60615:60612], addr_15153_7);

wire[31:0] addr_15154_7;

Selector_2 s15154_7(wires_3788_6[2], addr_3788_6, addr_positional[60619:60616], addr_15154_7);

wire[31:0] addr_15155_7;

Selector_2 s15155_7(wires_3788_6[3], addr_3788_6, addr_positional[60623:60620], addr_15155_7);

wire[31:0] addr_15156_7;

Selector_2 s15156_7(wires_3789_6[0], addr_3789_6, addr_positional[60627:60624], addr_15156_7);

wire[31:0] addr_15157_7;

Selector_2 s15157_7(wires_3789_6[1], addr_3789_6, addr_positional[60631:60628], addr_15157_7);

wire[31:0] addr_15158_7;

Selector_2 s15158_7(wires_3789_6[2], addr_3789_6, addr_positional[60635:60632], addr_15158_7);

wire[31:0] addr_15159_7;

Selector_2 s15159_7(wires_3789_6[3], addr_3789_6, addr_positional[60639:60636], addr_15159_7);

wire[31:0] addr_15160_7;

Selector_2 s15160_7(wires_3790_6[0], addr_3790_6, addr_positional[60643:60640], addr_15160_7);

wire[31:0] addr_15161_7;

Selector_2 s15161_7(wires_3790_6[1], addr_3790_6, addr_positional[60647:60644], addr_15161_7);

wire[31:0] addr_15162_7;

Selector_2 s15162_7(wires_3790_6[2], addr_3790_6, addr_positional[60651:60648], addr_15162_7);

wire[31:0] addr_15163_7;

Selector_2 s15163_7(wires_3790_6[3], addr_3790_6, addr_positional[60655:60652], addr_15163_7);

wire[31:0] addr_15164_7;

Selector_2 s15164_7(wires_3791_6[0], addr_3791_6, addr_positional[60659:60656], addr_15164_7);

wire[31:0] addr_15165_7;

Selector_2 s15165_7(wires_3791_6[1], addr_3791_6, addr_positional[60663:60660], addr_15165_7);

wire[31:0] addr_15166_7;

Selector_2 s15166_7(wires_3791_6[2], addr_3791_6, addr_positional[60667:60664], addr_15166_7);

wire[31:0] addr_15167_7;

Selector_2 s15167_7(wires_3791_6[3], addr_3791_6, addr_positional[60671:60668], addr_15167_7);

wire[31:0] addr_15168_7;

Selector_2 s15168_7(wires_3792_6[0], addr_3792_6, addr_positional[60675:60672], addr_15168_7);

wire[31:0] addr_15169_7;

Selector_2 s15169_7(wires_3792_6[1], addr_3792_6, addr_positional[60679:60676], addr_15169_7);

wire[31:0] addr_15170_7;

Selector_2 s15170_7(wires_3792_6[2], addr_3792_6, addr_positional[60683:60680], addr_15170_7);

wire[31:0] addr_15171_7;

Selector_2 s15171_7(wires_3792_6[3], addr_3792_6, addr_positional[60687:60684], addr_15171_7);

wire[31:0] addr_15172_7;

Selector_2 s15172_7(wires_3793_6[0], addr_3793_6, addr_positional[60691:60688], addr_15172_7);

wire[31:0] addr_15173_7;

Selector_2 s15173_7(wires_3793_6[1], addr_3793_6, addr_positional[60695:60692], addr_15173_7);

wire[31:0] addr_15174_7;

Selector_2 s15174_7(wires_3793_6[2], addr_3793_6, addr_positional[60699:60696], addr_15174_7);

wire[31:0] addr_15175_7;

Selector_2 s15175_7(wires_3793_6[3], addr_3793_6, addr_positional[60703:60700], addr_15175_7);

wire[31:0] addr_15176_7;

Selector_2 s15176_7(wires_3794_6[0], addr_3794_6, addr_positional[60707:60704], addr_15176_7);

wire[31:0] addr_15177_7;

Selector_2 s15177_7(wires_3794_6[1], addr_3794_6, addr_positional[60711:60708], addr_15177_7);

wire[31:0] addr_15178_7;

Selector_2 s15178_7(wires_3794_6[2], addr_3794_6, addr_positional[60715:60712], addr_15178_7);

wire[31:0] addr_15179_7;

Selector_2 s15179_7(wires_3794_6[3], addr_3794_6, addr_positional[60719:60716], addr_15179_7);

wire[31:0] addr_15180_7;

Selector_2 s15180_7(wires_3795_6[0], addr_3795_6, addr_positional[60723:60720], addr_15180_7);

wire[31:0] addr_15181_7;

Selector_2 s15181_7(wires_3795_6[1], addr_3795_6, addr_positional[60727:60724], addr_15181_7);

wire[31:0] addr_15182_7;

Selector_2 s15182_7(wires_3795_6[2], addr_3795_6, addr_positional[60731:60728], addr_15182_7);

wire[31:0] addr_15183_7;

Selector_2 s15183_7(wires_3795_6[3], addr_3795_6, addr_positional[60735:60732], addr_15183_7);

wire[31:0] addr_15184_7;

Selector_2 s15184_7(wires_3796_6[0], addr_3796_6, addr_positional[60739:60736], addr_15184_7);

wire[31:0] addr_15185_7;

Selector_2 s15185_7(wires_3796_6[1], addr_3796_6, addr_positional[60743:60740], addr_15185_7);

wire[31:0] addr_15186_7;

Selector_2 s15186_7(wires_3796_6[2], addr_3796_6, addr_positional[60747:60744], addr_15186_7);

wire[31:0] addr_15187_7;

Selector_2 s15187_7(wires_3796_6[3], addr_3796_6, addr_positional[60751:60748], addr_15187_7);

wire[31:0] addr_15188_7;

Selector_2 s15188_7(wires_3797_6[0], addr_3797_6, addr_positional[60755:60752], addr_15188_7);

wire[31:0] addr_15189_7;

Selector_2 s15189_7(wires_3797_6[1], addr_3797_6, addr_positional[60759:60756], addr_15189_7);

wire[31:0] addr_15190_7;

Selector_2 s15190_7(wires_3797_6[2], addr_3797_6, addr_positional[60763:60760], addr_15190_7);

wire[31:0] addr_15191_7;

Selector_2 s15191_7(wires_3797_6[3], addr_3797_6, addr_positional[60767:60764], addr_15191_7);

wire[31:0] addr_15192_7;

Selector_2 s15192_7(wires_3798_6[0], addr_3798_6, addr_positional[60771:60768], addr_15192_7);

wire[31:0] addr_15193_7;

Selector_2 s15193_7(wires_3798_6[1], addr_3798_6, addr_positional[60775:60772], addr_15193_7);

wire[31:0] addr_15194_7;

Selector_2 s15194_7(wires_3798_6[2], addr_3798_6, addr_positional[60779:60776], addr_15194_7);

wire[31:0] addr_15195_7;

Selector_2 s15195_7(wires_3798_6[3], addr_3798_6, addr_positional[60783:60780], addr_15195_7);

wire[31:0] addr_15196_7;

Selector_2 s15196_7(wires_3799_6[0], addr_3799_6, addr_positional[60787:60784], addr_15196_7);

wire[31:0] addr_15197_7;

Selector_2 s15197_7(wires_3799_6[1], addr_3799_6, addr_positional[60791:60788], addr_15197_7);

wire[31:0] addr_15198_7;

Selector_2 s15198_7(wires_3799_6[2], addr_3799_6, addr_positional[60795:60792], addr_15198_7);

wire[31:0] addr_15199_7;

Selector_2 s15199_7(wires_3799_6[3], addr_3799_6, addr_positional[60799:60796], addr_15199_7);

wire[31:0] addr_15200_7;

Selector_2 s15200_7(wires_3800_6[0], addr_3800_6, addr_positional[60803:60800], addr_15200_7);

wire[31:0] addr_15201_7;

Selector_2 s15201_7(wires_3800_6[1], addr_3800_6, addr_positional[60807:60804], addr_15201_7);

wire[31:0] addr_15202_7;

Selector_2 s15202_7(wires_3800_6[2], addr_3800_6, addr_positional[60811:60808], addr_15202_7);

wire[31:0] addr_15203_7;

Selector_2 s15203_7(wires_3800_6[3], addr_3800_6, addr_positional[60815:60812], addr_15203_7);

wire[31:0] addr_15204_7;

Selector_2 s15204_7(wires_3801_6[0], addr_3801_6, addr_positional[60819:60816], addr_15204_7);

wire[31:0] addr_15205_7;

Selector_2 s15205_7(wires_3801_6[1], addr_3801_6, addr_positional[60823:60820], addr_15205_7);

wire[31:0] addr_15206_7;

Selector_2 s15206_7(wires_3801_6[2], addr_3801_6, addr_positional[60827:60824], addr_15206_7);

wire[31:0] addr_15207_7;

Selector_2 s15207_7(wires_3801_6[3], addr_3801_6, addr_positional[60831:60828], addr_15207_7);

wire[31:0] addr_15208_7;

Selector_2 s15208_7(wires_3802_6[0], addr_3802_6, addr_positional[60835:60832], addr_15208_7);

wire[31:0] addr_15209_7;

Selector_2 s15209_7(wires_3802_6[1], addr_3802_6, addr_positional[60839:60836], addr_15209_7);

wire[31:0] addr_15210_7;

Selector_2 s15210_7(wires_3802_6[2], addr_3802_6, addr_positional[60843:60840], addr_15210_7);

wire[31:0] addr_15211_7;

Selector_2 s15211_7(wires_3802_6[3], addr_3802_6, addr_positional[60847:60844], addr_15211_7);

wire[31:0] addr_15212_7;

Selector_2 s15212_7(wires_3803_6[0], addr_3803_6, addr_positional[60851:60848], addr_15212_7);

wire[31:0] addr_15213_7;

Selector_2 s15213_7(wires_3803_6[1], addr_3803_6, addr_positional[60855:60852], addr_15213_7);

wire[31:0] addr_15214_7;

Selector_2 s15214_7(wires_3803_6[2], addr_3803_6, addr_positional[60859:60856], addr_15214_7);

wire[31:0] addr_15215_7;

Selector_2 s15215_7(wires_3803_6[3], addr_3803_6, addr_positional[60863:60860], addr_15215_7);

wire[31:0] addr_15216_7;

Selector_2 s15216_7(wires_3804_6[0], addr_3804_6, addr_positional[60867:60864], addr_15216_7);

wire[31:0] addr_15217_7;

Selector_2 s15217_7(wires_3804_6[1], addr_3804_6, addr_positional[60871:60868], addr_15217_7);

wire[31:0] addr_15218_7;

Selector_2 s15218_7(wires_3804_6[2], addr_3804_6, addr_positional[60875:60872], addr_15218_7);

wire[31:0] addr_15219_7;

Selector_2 s15219_7(wires_3804_6[3], addr_3804_6, addr_positional[60879:60876], addr_15219_7);

wire[31:0] addr_15220_7;

Selector_2 s15220_7(wires_3805_6[0], addr_3805_6, addr_positional[60883:60880], addr_15220_7);

wire[31:0] addr_15221_7;

Selector_2 s15221_7(wires_3805_6[1], addr_3805_6, addr_positional[60887:60884], addr_15221_7);

wire[31:0] addr_15222_7;

Selector_2 s15222_7(wires_3805_6[2], addr_3805_6, addr_positional[60891:60888], addr_15222_7);

wire[31:0] addr_15223_7;

Selector_2 s15223_7(wires_3805_6[3], addr_3805_6, addr_positional[60895:60892], addr_15223_7);

wire[31:0] addr_15224_7;

Selector_2 s15224_7(wires_3806_6[0], addr_3806_6, addr_positional[60899:60896], addr_15224_7);

wire[31:0] addr_15225_7;

Selector_2 s15225_7(wires_3806_6[1], addr_3806_6, addr_positional[60903:60900], addr_15225_7);

wire[31:0] addr_15226_7;

Selector_2 s15226_7(wires_3806_6[2], addr_3806_6, addr_positional[60907:60904], addr_15226_7);

wire[31:0] addr_15227_7;

Selector_2 s15227_7(wires_3806_6[3], addr_3806_6, addr_positional[60911:60908], addr_15227_7);

wire[31:0] addr_15228_7;

Selector_2 s15228_7(wires_3807_6[0], addr_3807_6, addr_positional[60915:60912], addr_15228_7);

wire[31:0] addr_15229_7;

Selector_2 s15229_7(wires_3807_6[1], addr_3807_6, addr_positional[60919:60916], addr_15229_7);

wire[31:0] addr_15230_7;

Selector_2 s15230_7(wires_3807_6[2], addr_3807_6, addr_positional[60923:60920], addr_15230_7);

wire[31:0] addr_15231_7;

Selector_2 s15231_7(wires_3807_6[3], addr_3807_6, addr_positional[60927:60924], addr_15231_7);

wire[31:0] addr_15232_7;

Selector_2 s15232_7(wires_3808_6[0], addr_3808_6, addr_positional[60931:60928], addr_15232_7);

wire[31:0] addr_15233_7;

Selector_2 s15233_7(wires_3808_6[1], addr_3808_6, addr_positional[60935:60932], addr_15233_7);

wire[31:0] addr_15234_7;

Selector_2 s15234_7(wires_3808_6[2], addr_3808_6, addr_positional[60939:60936], addr_15234_7);

wire[31:0] addr_15235_7;

Selector_2 s15235_7(wires_3808_6[3], addr_3808_6, addr_positional[60943:60940], addr_15235_7);

wire[31:0] addr_15236_7;

Selector_2 s15236_7(wires_3809_6[0], addr_3809_6, addr_positional[60947:60944], addr_15236_7);

wire[31:0] addr_15237_7;

Selector_2 s15237_7(wires_3809_6[1], addr_3809_6, addr_positional[60951:60948], addr_15237_7);

wire[31:0] addr_15238_7;

Selector_2 s15238_7(wires_3809_6[2], addr_3809_6, addr_positional[60955:60952], addr_15238_7);

wire[31:0] addr_15239_7;

Selector_2 s15239_7(wires_3809_6[3], addr_3809_6, addr_positional[60959:60956], addr_15239_7);

wire[31:0] addr_15240_7;

Selector_2 s15240_7(wires_3810_6[0], addr_3810_6, addr_positional[60963:60960], addr_15240_7);

wire[31:0] addr_15241_7;

Selector_2 s15241_7(wires_3810_6[1], addr_3810_6, addr_positional[60967:60964], addr_15241_7);

wire[31:0] addr_15242_7;

Selector_2 s15242_7(wires_3810_6[2], addr_3810_6, addr_positional[60971:60968], addr_15242_7);

wire[31:0] addr_15243_7;

Selector_2 s15243_7(wires_3810_6[3], addr_3810_6, addr_positional[60975:60972], addr_15243_7);

wire[31:0] addr_15244_7;

Selector_2 s15244_7(wires_3811_6[0], addr_3811_6, addr_positional[60979:60976], addr_15244_7);

wire[31:0] addr_15245_7;

Selector_2 s15245_7(wires_3811_6[1], addr_3811_6, addr_positional[60983:60980], addr_15245_7);

wire[31:0] addr_15246_7;

Selector_2 s15246_7(wires_3811_6[2], addr_3811_6, addr_positional[60987:60984], addr_15246_7);

wire[31:0] addr_15247_7;

Selector_2 s15247_7(wires_3811_6[3], addr_3811_6, addr_positional[60991:60988], addr_15247_7);

wire[31:0] addr_15248_7;

Selector_2 s15248_7(wires_3812_6[0], addr_3812_6, addr_positional[60995:60992], addr_15248_7);

wire[31:0] addr_15249_7;

Selector_2 s15249_7(wires_3812_6[1], addr_3812_6, addr_positional[60999:60996], addr_15249_7);

wire[31:0] addr_15250_7;

Selector_2 s15250_7(wires_3812_6[2], addr_3812_6, addr_positional[61003:61000], addr_15250_7);

wire[31:0] addr_15251_7;

Selector_2 s15251_7(wires_3812_6[3], addr_3812_6, addr_positional[61007:61004], addr_15251_7);

wire[31:0] addr_15252_7;

Selector_2 s15252_7(wires_3813_6[0], addr_3813_6, addr_positional[61011:61008], addr_15252_7);

wire[31:0] addr_15253_7;

Selector_2 s15253_7(wires_3813_6[1], addr_3813_6, addr_positional[61015:61012], addr_15253_7);

wire[31:0] addr_15254_7;

Selector_2 s15254_7(wires_3813_6[2], addr_3813_6, addr_positional[61019:61016], addr_15254_7);

wire[31:0] addr_15255_7;

Selector_2 s15255_7(wires_3813_6[3], addr_3813_6, addr_positional[61023:61020], addr_15255_7);

wire[31:0] addr_15256_7;

Selector_2 s15256_7(wires_3814_6[0], addr_3814_6, addr_positional[61027:61024], addr_15256_7);

wire[31:0] addr_15257_7;

Selector_2 s15257_7(wires_3814_6[1], addr_3814_6, addr_positional[61031:61028], addr_15257_7);

wire[31:0] addr_15258_7;

Selector_2 s15258_7(wires_3814_6[2], addr_3814_6, addr_positional[61035:61032], addr_15258_7);

wire[31:0] addr_15259_7;

Selector_2 s15259_7(wires_3814_6[3], addr_3814_6, addr_positional[61039:61036], addr_15259_7);

wire[31:0] addr_15260_7;

Selector_2 s15260_7(wires_3815_6[0], addr_3815_6, addr_positional[61043:61040], addr_15260_7);

wire[31:0] addr_15261_7;

Selector_2 s15261_7(wires_3815_6[1], addr_3815_6, addr_positional[61047:61044], addr_15261_7);

wire[31:0] addr_15262_7;

Selector_2 s15262_7(wires_3815_6[2], addr_3815_6, addr_positional[61051:61048], addr_15262_7);

wire[31:0] addr_15263_7;

Selector_2 s15263_7(wires_3815_6[3], addr_3815_6, addr_positional[61055:61052], addr_15263_7);

wire[31:0] addr_15264_7;

Selector_2 s15264_7(wires_3816_6[0], addr_3816_6, addr_positional[61059:61056], addr_15264_7);

wire[31:0] addr_15265_7;

Selector_2 s15265_7(wires_3816_6[1], addr_3816_6, addr_positional[61063:61060], addr_15265_7);

wire[31:0] addr_15266_7;

Selector_2 s15266_7(wires_3816_6[2], addr_3816_6, addr_positional[61067:61064], addr_15266_7);

wire[31:0] addr_15267_7;

Selector_2 s15267_7(wires_3816_6[3], addr_3816_6, addr_positional[61071:61068], addr_15267_7);

wire[31:0] addr_15268_7;

Selector_2 s15268_7(wires_3817_6[0], addr_3817_6, addr_positional[61075:61072], addr_15268_7);

wire[31:0] addr_15269_7;

Selector_2 s15269_7(wires_3817_6[1], addr_3817_6, addr_positional[61079:61076], addr_15269_7);

wire[31:0] addr_15270_7;

Selector_2 s15270_7(wires_3817_6[2], addr_3817_6, addr_positional[61083:61080], addr_15270_7);

wire[31:0] addr_15271_7;

Selector_2 s15271_7(wires_3817_6[3], addr_3817_6, addr_positional[61087:61084], addr_15271_7);

wire[31:0] addr_15272_7;

Selector_2 s15272_7(wires_3818_6[0], addr_3818_6, addr_positional[61091:61088], addr_15272_7);

wire[31:0] addr_15273_7;

Selector_2 s15273_7(wires_3818_6[1], addr_3818_6, addr_positional[61095:61092], addr_15273_7);

wire[31:0] addr_15274_7;

Selector_2 s15274_7(wires_3818_6[2], addr_3818_6, addr_positional[61099:61096], addr_15274_7);

wire[31:0] addr_15275_7;

Selector_2 s15275_7(wires_3818_6[3], addr_3818_6, addr_positional[61103:61100], addr_15275_7);

wire[31:0] addr_15276_7;

Selector_2 s15276_7(wires_3819_6[0], addr_3819_6, addr_positional[61107:61104], addr_15276_7);

wire[31:0] addr_15277_7;

Selector_2 s15277_7(wires_3819_6[1], addr_3819_6, addr_positional[61111:61108], addr_15277_7);

wire[31:0] addr_15278_7;

Selector_2 s15278_7(wires_3819_6[2], addr_3819_6, addr_positional[61115:61112], addr_15278_7);

wire[31:0] addr_15279_7;

Selector_2 s15279_7(wires_3819_6[3], addr_3819_6, addr_positional[61119:61116], addr_15279_7);

wire[31:0] addr_15280_7;

Selector_2 s15280_7(wires_3820_6[0], addr_3820_6, addr_positional[61123:61120], addr_15280_7);

wire[31:0] addr_15281_7;

Selector_2 s15281_7(wires_3820_6[1], addr_3820_6, addr_positional[61127:61124], addr_15281_7);

wire[31:0] addr_15282_7;

Selector_2 s15282_7(wires_3820_6[2], addr_3820_6, addr_positional[61131:61128], addr_15282_7);

wire[31:0] addr_15283_7;

Selector_2 s15283_7(wires_3820_6[3], addr_3820_6, addr_positional[61135:61132], addr_15283_7);

wire[31:0] addr_15284_7;

Selector_2 s15284_7(wires_3821_6[0], addr_3821_6, addr_positional[61139:61136], addr_15284_7);

wire[31:0] addr_15285_7;

Selector_2 s15285_7(wires_3821_6[1], addr_3821_6, addr_positional[61143:61140], addr_15285_7);

wire[31:0] addr_15286_7;

Selector_2 s15286_7(wires_3821_6[2], addr_3821_6, addr_positional[61147:61144], addr_15286_7);

wire[31:0] addr_15287_7;

Selector_2 s15287_7(wires_3821_6[3], addr_3821_6, addr_positional[61151:61148], addr_15287_7);

wire[31:0] addr_15288_7;

Selector_2 s15288_7(wires_3822_6[0], addr_3822_6, addr_positional[61155:61152], addr_15288_7);

wire[31:0] addr_15289_7;

Selector_2 s15289_7(wires_3822_6[1], addr_3822_6, addr_positional[61159:61156], addr_15289_7);

wire[31:0] addr_15290_7;

Selector_2 s15290_7(wires_3822_6[2], addr_3822_6, addr_positional[61163:61160], addr_15290_7);

wire[31:0] addr_15291_7;

Selector_2 s15291_7(wires_3822_6[3], addr_3822_6, addr_positional[61167:61164], addr_15291_7);

wire[31:0] addr_15292_7;

Selector_2 s15292_7(wires_3823_6[0], addr_3823_6, addr_positional[61171:61168], addr_15292_7);

wire[31:0] addr_15293_7;

Selector_2 s15293_7(wires_3823_6[1], addr_3823_6, addr_positional[61175:61172], addr_15293_7);

wire[31:0] addr_15294_7;

Selector_2 s15294_7(wires_3823_6[2], addr_3823_6, addr_positional[61179:61176], addr_15294_7);

wire[31:0] addr_15295_7;

Selector_2 s15295_7(wires_3823_6[3], addr_3823_6, addr_positional[61183:61180], addr_15295_7);

wire[31:0] addr_15296_7;

Selector_2 s15296_7(wires_3824_6[0], addr_3824_6, addr_positional[61187:61184], addr_15296_7);

wire[31:0] addr_15297_7;

Selector_2 s15297_7(wires_3824_6[1], addr_3824_6, addr_positional[61191:61188], addr_15297_7);

wire[31:0] addr_15298_7;

Selector_2 s15298_7(wires_3824_6[2], addr_3824_6, addr_positional[61195:61192], addr_15298_7);

wire[31:0] addr_15299_7;

Selector_2 s15299_7(wires_3824_6[3], addr_3824_6, addr_positional[61199:61196], addr_15299_7);

wire[31:0] addr_15300_7;

Selector_2 s15300_7(wires_3825_6[0], addr_3825_6, addr_positional[61203:61200], addr_15300_7);

wire[31:0] addr_15301_7;

Selector_2 s15301_7(wires_3825_6[1], addr_3825_6, addr_positional[61207:61204], addr_15301_7);

wire[31:0] addr_15302_7;

Selector_2 s15302_7(wires_3825_6[2], addr_3825_6, addr_positional[61211:61208], addr_15302_7);

wire[31:0] addr_15303_7;

Selector_2 s15303_7(wires_3825_6[3], addr_3825_6, addr_positional[61215:61212], addr_15303_7);

wire[31:0] addr_15304_7;

Selector_2 s15304_7(wires_3826_6[0], addr_3826_6, addr_positional[61219:61216], addr_15304_7);

wire[31:0] addr_15305_7;

Selector_2 s15305_7(wires_3826_6[1], addr_3826_6, addr_positional[61223:61220], addr_15305_7);

wire[31:0] addr_15306_7;

Selector_2 s15306_7(wires_3826_6[2], addr_3826_6, addr_positional[61227:61224], addr_15306_7);

wire[31:0] addr_15307_7;

Selector_2 s15307_7(wires_3826_6[3], addr_3826_6, addr_positional[61231:61228], addr_15307_7);

wire[31:0] addr_15308_7;

Selector_2 s15308_7(wires_3827_6[0], addr_3827_6, addr_positional[61235:61232], addr_15308_7);

wire[31:0] addr_15309_7;

Selector_2 s15309_7(wires_3827_6[1], addr_3827_6, addr_positional[61239:61236], addr_15309_7);

wire[31:0] addr_15310_7;

Selector_2 s15310_7(wires_3827_6[2], addr_3827_6, addr_positional[61243:61240], addr_15310_7);

wire[31:0] addr_15311_7;

Selector_2 s15311_7(wires_3827_6[3], addr_3827_6, addr_positional[61247:61244], addr_15311_7);

wire[31:0] addr_15312_7;

Selector_2 s15312_7(wires_3828_6[0], addr_3828_6, addr_positional[61251:61248], addr_15312_7);

wire[31:0] addr_15313_7;

Selector_2 s15313_7(wires_3828_6[1], addr_3828_6, addr_positional[61255:61252], addr_15313_7);

wire[31:0] addr_15314_7;

Selector_2 s15314_7(wires_3828_6[2], addr_3828_6, addr_positional[61259:61256], addr_15314_7);

wire[31:0] addr_15315_7;

Selector_2 s15315_7(wires_3828_6[3], addr_3828_6, addr_positional[61263:61260], addr_15315_7);

wire[31:0] addr_15316_7;

Selector_2 s15316_7(wires_3829_6[0], addr_3829_6, addr_positional[61267:61264], addr_15316_7);

wire[31:0] addr_15317_7;

Selector_2 s15317_7(wires_3829_6[1], addr_3829_6, addr_positional[61271:61268], addr_15317_7);

wire[31:0] addr_15318_7;

Selector_2 s15318_7(wires_3829_6[2], addr_3829_6, addr_positional[61275:61272], addr_15318_7);

wire[31:0] addr_15319_7;

Selector_2 s15319_7(wires_3829_6[3], addr_3829_6, addr_positional[61279:61276], addr_15319_7);

wire[31:0] addr_15320_7;

Selector_2 s15320_7(wires_3830_6[0], addr_3830_6, addr_positional[61283:61280], addr_15320_7);

wire[31:0] addr_15321_7;

Selector_2 s15321_7(wires_3830_6[1], addr_3830_6, addr_positional[61287:61284], addr_15321_7);

wire[31:0] addr_15322_7;

Selector_2 s15322_7(wires_3830_6[2], addr_3830_6, addr_positional[61291:61288], addr_15322_7);

wire[31:0] addr_15323_7;

Selector_2 s15323_7(wires_3830_6[3], addr_3830_6, addr_positional[61295:61292], addr_15323_7);

wire[31:0] addr_15324_7;

Selector_2 s15324_7(wires_3831_6[0], addr_3831_6, addr_positional[61299:61296], addr_15324_7);

wire[31:0] addr_15325_7;

Selector_2 s15325_7(wires_3831_6[1], addr_3831_6, addr_positional[61303:61300], addr_15325_7);

wire[31:0] addr_15326_7;

Selector_2 s15326_7(wires_3831_6[2], addr_3831_6, addr_positional[61307:61304], addr_15326_7);

wire[31:0] addr_15327_7;

Selector_2 s15327_7(wires_3831_6[3], addr_3831_6, addr_positional[61311:61308], addr_15327_7);

wire[31:0] addr_15328_7;

Selector_2 s15328_7(wires_3832_6[0], addr_3832_6, addr_positional[61315:61312], addr_15328_7);

wire[31:0] addr_15329_7;

Selector_2 s15329_7(wires_3832_6[1], addr_3832_6, addr_positional[61319:61316], addr_15329_7);

wire[31:0] addr_15330_7;

Selector_2 s15330_7(wires_3832_6[2], addr_3832_6, addr_positional[61323:61320], addr_15330_7);

wire[31:0] addr_15331_7;

Selector_2 s15331_7(wires_3832_6[3], addr_3832_6, addr_positional[61327:61324], addr_15331_7);

wire[31:0] addr_15332_7;

Selector_2 s15332_7(wires_3833_6[0], addr_3833_6, addr_positional[61331:61328], addr_15332_7);

wire[31:0] addr_15333_7;

Selector_2 s15333_7(wires_3833_6[1], addr_3833_6, addr_positional[61335:61332], addr_15333_7);

wire[31:0] addr_15334_7;

Selector_2 s15334_7(wires_3833_6[2], addr_3833_6, addr_positional[61339:61336], addr_15334_7);

wire[31:0] addr_15335_7;

Selector_2 s15335_7(wires_3833_6[3], addr_3833_6, addr_positional[61343:61340], addr_15335_7);

wire[31:0] addr_15336_7;

Selector_2 s15336_7(wires_3834_6[0], addr_3834_6, addr_positional[61347:61344], addr_15336_7);

wire[31:0] addr_15337_7;

Selector_2 s15337_7(wires_3834_6[1], addr_3834_6, addr_positional[61351:61348], addr_15337_7);

wire[31:0] addr_15338_7;

Selector_2 s15338_7(wires_3834_6[2], addr_3834_6, addr_positional[61355:61352], addr_15338_7);

wire[31:0] addr_15339_7;

Selector_2 s15339_7(wires_3834_6[3], addr_3834_6, addr_positional[61359:61356], addr_15339_7);

wire[31:0] addr_15340_7;

Selector_2 s15340_7(wires_3835_6[0], addr_3835_6, addr_positional[61363:61360], addr_15340_7);

wire[31:0] addr_15341_7;

Selector_2 s15341_7(wires_3835_6[1], addr_3835_6, addr_positional[61367:61364], addr_15341_7);

wire[31:0] addr_15342_7;

Selector_2 s15342_7(wires_3835_6[2], addr_3835_6, addr_positional[61371:61368], addr_15342_7);

wire[31:0] addr_15343_7;

Selector_2 s15343_7(wires_3835_6[3], addr_3835_6, addr_positional[61375:61372], addr_15343_7);

wire[31:0] addr_15344_7;

Selector_2 s15344_7(wires_3836_6[0], addr_3836_6, addr_positional[61379:61376], addr_15344_7);

wire[31:0] addr_15345_7;

Selector_2 s15345_7(wires_3836_6[1], addr_3836_6, addr_positional[61383:61380], addr_15345_7);

wire[31:0] addr_15346_7;

Selector_2 s15346_7(wires_3836_6[2], addr_3836_6, addr_positional[61387:61384], addr_15346_7);

wire[31:0] addr_15347_7;

Selector_2 s15347_7(wires_3836_6[3], addr_3836_6, addr_positional[61391:61388], addr_15347_7);

wire[31:0] addr_15348_7;

Selector_2 s15348_7(wires_3837_6[0], addr_3837_6, addr_positional[61395:61392], addr_15348_7);

wire[31:0] addr_15349_7;

Selector_2 s15349_7(wires_3837_6[1], addr_3837_6, addr_positional[61399:61396], addr_15349_7);

wire[31:0] addr_15350_7;

Selector_2 s15350_7(wires_3837_6[2], addr_3837_6, addr_positional[61403:61400], addr_15350_7);

wire[31:0] addr_15351_7;

Selector_2 s15351_7(wires_3837_6[3], addr_3837_6, addr_positional[61407:61404], addr_15351_7);

wire[31:0] addr_15352_7;

Selector_2 s15352_7(wires_3838_6[0], addr_3838_6, addr_positional[61411:61408], addr_15352_7);

wire[31:0] addr_15353_7;

Selector_2 s15353_7(wires_3838_6[1], addr_3838_6, addr_positional[61415:61412], addr_15353_7);

wire[31:0] addr_15354_7;

Selector_2 s15354_7(wires_3838_6[2], addr_3838_6, addr_positional[61419:61416], addr_15354_7);

wire[31:0] addr_15355_7;

Selector_2 s15355_7(wires_3838_6[3], addr_3838_6, addr_positional[61423:61420], addr_15355_7);

wire[31:0] addr_15356_7;

Selector_2 s15356_7(wires_3839_6[0], addr_3839_6, addr_positional[61427:61424], addr_15356_7);

wire[31:0] addr_15357_7;

Selector_2 s15357_7(wires_3839_6[1], addr_3839_6, addr_positional[61431:61428], addr_15357_7);

wire[31:0] addr_15358_7;

Selector_2 s15358_7(wires_3839_6[2], addr_3839_6, addr_positional[61435:61432], addr_15358_7);

wire[31:0] addr_15359_7;

Selector_2 s15359_7(wires_3839_6[3], addr_3839_6, addr_positional[61439:61436], addr_15359_7);

wire[31:0] addr_15360_7;

Selector_2 s15360_7(wires_3840_6[0], addr_3840_6, addr_positional[61443:61440], addr_15360_7);

wire[31:0] addr_15361_7;

Selector_2 s15361_7(wires_3840_6[1], addr_3840_6, addr_positional[61447:61444], addr_15361_7);

wire[31:0] addr_15362_7;

Selector_2 s15362_7(wires_3840_6[2], addr_3840_6, addr_positional[61451:61448], addr_15362_7);

wire[31:0] addr_15363_7;

Selector_2 s15363_7(wires_3840_6[3], addr_3840_6, addr_positional[61455:61452], addr_15363_7);

wire[31:0] addr_15364_7;

Selector_2 s15364_7(wires_3841_6[0], addr_3841_6, addr_positional[61459:61456], addr_15364_7);

wire[31:0] addr_15365_7;

Selector_2 s15365_7(wires_3841_6[1], addr_3841_6, addr_positional[61463:61460], addr_15365_7);

wire[31:0] addr_15366_7;

Selector_2 s15366_7(wires_3841_6[2], addr_3841_6, addr_positional[61467:61464], addr_15366_7);

wire[31:0] addr_15367_7;

Selector_2 s15367_7(wires_3841_6[3], addr_3841_6, addr_positional[61471:61468], addr_15367_7);

wire[31:0] addr_15368_7;

Selector_2 s15368_7(wires_3842_6[0], addr_3842_6, addr_positional[61475:61472], addr_15368_7);

wire[31:0] addr_15369_7;

Selector_2 s15369_7(wires_3842_6[1], addr_3842_6, addr_positional[61479:61476], addr_15369_7);

wire[31:0] addr_15370_7;

Selector_2 s15370_7(wires_3842_6[2], addr_3842_6, addr_positional[61483:61480], addr_15370_7);

wire[31:0] addr_15371_7;

Selector_2 s15371_7(wires_3842_6[3], addr_3842_6, addr_positional[61487:61484], addr_15371_7);

wire[31:0] addr_15372_7;

Selector_2 s15372_7(wires_3843_6[0], addr_3843_6, addr_positional[61491:61488], addr_15372_7);

wire[31:0] addr_15373_7;

Selector_2 s15373_7(wires_3843_6[1], addr_3843_6, addr_positional[61495:61492], addr_15373_7);

wire[31:0] addr_15374_7;

Selector_2 s15374_7(wires_3843_6[2], addr_3843_6, addr_positional[61499:61496], addr_15374_7);

wire[31:0] addr_15375_7;

Selector_2 s15375_7(wires_3843_6[3], addr_3843_6, addr_positional[61503:61500], addr_15375_7);

wire[31:0] addr_15376_7;

Selector_2 s15376_7(wires_3844_6[0], addr_3844_6, addr_positional[61507:61504], addr_15376_7);

wire[31:0] addr_15377_7;

Selector_2 s15377_7(wires_3844_6[1], addr_3844_6, addr_positional[61511:61508], addr_15377_7);

wire[31:0] addr_15378_7;

Selector_2 s15378_7(wires_3844_6[2], addr_3844_6, addr_positional[61515:61512], addr_15378_7);

wire[31:0] addr_15379_7;

Selector_2 s15379_7(wires_3844_6[3], addr_3844_6, addr_positional[61519:61516], addr_15379_7);

wire[31:0] addr_15380_7;

Selector_2 s15380_7(wires_3845_6[0], addr_3845_6, addr_positional[61523:61520], addr_15380_7);

wire[31:0] addr_15381_7;

Selector_2 s15381_7(wires_3845_6[1], addr_3845_6, addr_positional[61527:61524], addr_15381_7);

wire[31:0] addr_15382_7;

Selector_2 s15382_7(wires_3845_6[2], addr_3845_6, addr_positional[61531:61528], addr_15382_7);

wire[31:0] addr_15383_7;

Selector_2 s15383_7(wires_3845_6[3], addr_3845_6, addr_positional[61535:61532], addr_15383_7);

wire[31:0] addr_15384_7;

Selector_2 s15384_7(wires_3846_6[0], addr_3846_6, addr_positional[61539:61536], addr_15384_7);

wire[31:0] addr_15385_7;

Selector_2 s15385_7(wires_3846_6[1], addr_3846_6, addr_positional[61543:61540], addr_15385_7);

wire[31:0] addr_15386_7;

Selector_2 s15386_7(wires_3846_6[2], addr_3846_6, addr_positional[61547:61544], addr_15386_7);

wire[31:0] addr_15387_7;

Selector_2 s15387_7(wires_3846_6[3], addr_3846_6, addr_positional[61551:61548], addr_15387_7);

wire[31:0] addr_15388_7;

Selector_2 s15388_7(wires_3847_6[0], addr_3847_6, addr_positional[61555:61552], addr_15388_7);

wire[31:0] addr_15389_7;

Selector_2 s15389_7(wires_3847_6[1], addr_3847_6, addr_positional[61559:61556], addr_15389_7);

wire[31:0] addr_15390_7;

Selector_2 s15390_7(wires_3847_6[2], addr_3847_6, addr_positional[61563:61560], addr_15390_7);

wire[31:0] addr_15391_7;

Selector_2 s15391_7(wires_3847_6[3], addr_3847_6, addr_positional[61567:61564], addr_15391_7);

wire[31:0] addr_15392_7;

Selector_2 s15392_7(wires_3848_6[0], addr_3848_6, addr_positional[61571:61568], addr_15392_7);

wire[31:0] addr_15393_7;

Selector_2 s15393_7(wires_3848_6[1], addr_3848_6, addr_positional[61575:61572], addr_15393_7);

wire[31:0] addr_15394_7;

Selector_2 s15394_7(wires_3848_6[2], addr_3848_6, addr_positional[61579:61576], addr_15394_7);

wire[31:0] addr_15395_7;

Selector_2 s15395_7(wires_3848_6[3], addr_3848_6, addr_positional[61583:61580], addr_15395_7);

wire[31:0] addr_15396_7;

Selector_2 s15396_7(wires_3849_6[0], addr_3849_6, addr_positional[61587:61584], addr_15396_7);

wire[31:0] addr_15397_7;

Selector_2 s15397_7(wires_3849_6[1], addr_3849_6, addr_positional[61591:61588], addr_15397_7);

wire[31:0] addr_15398_7;

Selector_2 s15398_7(wires_3849_6[2], addr_3849_6, addr_positional[61595:61592], addr_15398_7);

wire[31:0] addr_15399_7;

Selector_2 s15399_7(wires_3849_6[3], addr_3849_6, addr_positional[61599:61596], addr_15399_7);

wire[31:0] addr_15400_7;

Selector_2 s15400_7(wires_3850_6[0], addr_3850_6, addr_positional[61603:61600], addr_15400_7);

wire[31:0] addr_15401_7;

Selector_2 s15401_7(wires_3850_6[1], addr_3850_6, addr_positional[61607:61604], addr_15401_7);

wire[31:0] addr_15402_7;

Selector_2 s15402_7(wires_3850_6[2], addr_3850_6, addr_positional[61611:61608], addr_15402_7);

wire[31:0] addr_15403_7;

Selector_2 s15403_7(wires_3850_6[3], addr_3850_6, addr_positional[61615:61612], addr_15403_7);

wire[31:0] addr_15404_7;

Selector_2 s15404_7(wires_3851_6[0], addr_3851_6, addr_positional[61619:61616], addr_15404_7);

wire[31:0] addr_15405_7;

Selector_2 s15405_7(wires_3851_6[1], addr_3851_6, addr_positional[61623:61620], addr_15405_7);

wire[31:0] addr_15406_7;

Selector_2 s15406_7(wires_3851_6[2], addr_3851_6, addr_positional[61627:61624], addr_15406_7);

wire[31:0] addr_15407_7;

Selector_2 s15407_7(wires_3851_6[3], addr_3851_6, addr_positional[61631:61628], addr_15407_7);

wire[31:0] addr_15408_7;

Selector_2 s15408_7(wires_3852_6[0], addr_3852_6, addr_positional[61635:61632], addr_15408_7);

wire[31:0] addr_15409_7;

Selector_2 s15409_7(wires_3852_6[1], addr_3852_6, addr_positional[61639:61636], addr_15409_7);

wire[31:0] addr_15410_7;

Selector_2 s15410_7(wires_3852_6[2], addr_3852_6, addr_positional[61643:61640], addr_15410_7);

wire[31:0] addr_15411_7;

Selector_2 s15411_7(wires_3852_6[3], addr_3852_6, addr_positional[61647:61644], addr_15411_7);

wire[31:0] addr_15412_7;

Selector_2 s15412_7(wires_3853_6[0], addr_3853_6, addr_positional[61651:61648], addr_15412_7);

wire[31:0] addr_15413_7;

Selector_2 s15413_7(wires_3853_6[1], addr_3853_6, addr_positional[61655:61652], addr_15413_7);

wire[31:0] addr_15414_7;

Selector_2 s15414_7(wires_3853_6[2], addr_3853_6, addr_positional[61659:61656], addr_15414_7);

wire[31:0] addr_15415_7;

Selector_2 s15415_7(wires_3853_6[3], addr_3853_6, addr_positional[61663:61660], addr_15415_7);

wire[31:0] addr_15416_7;

Selector_2 s15416_7(wires_3854_6[0], addr_3854_6, addr_positional[61667:61664], addr_15416_7);

wire[31:0] addr_15417_7;

Selector_2 s15417_7(wires_3854_6[1], addr_3854_6, addr_positional[61671:61668], addr_15417_7);

wire[31:0] addr_15418_7;

Selector_2 s15418_7(wires_3854_6[2], addr_3854_6, addr_positional[61675:61672], addr_15418_7);

wire[31:0] addr_15419_7;

Selector_2 s15419_7(wires_3854_6[3], addr_3854_6, addr_positional[61679:61676], addr_15419_7);

wire[31:0] addr_15420_7;

Selector_2 s15420_7(wires_3855_6[0], addr_3855_6, addr_positional[61683:61680], addr_15420_7);

wire[31:0] addr_15421_7;

Selector_2 s15421_7(wires_3855_6[1], addr_3855_6, addr_positional[61687:61684], addr_15421_7);

wire[31:0] addr_15422_7;

Selector_2 s15422_7(wires_3855_6[2], addr_3855_6, addr_positional[61691:61688], addr_15422_7);

wire[31:0] addr_15423_7;

Selector_2 s15423_7(wires_3855_6[3], addr_3855_6, addr_positional[61695:61692], addr_15423_7);

wire[31:0] addr_15424_7;

Selector_2 s15424_7(wires_3856_6[0], addr_3856_6, addr_positional[61699:61696], addr_15424_7);

wire[31:0] addr_15425_7;

Selector_2 s15425_7(wires_3856_6[1], addr_3856_6, addr_positional[61703:61700], addr_15425_7);

wire[31:0] addr_15426_7;

Selector_2 s15426_7(wires_3856_6[2], addr_3856_6, addr_positional[61707:61704], addr_15426_7);

wire[31:0] addr_15427_7;

Selector_2 s15427_7(wires_3856_6[3], addr_3856_6, addr_positional[61711:61708], addr_15427_7);

wire[31:0] addr_15428_7;

Selector_2 s15428_7(wires_3857_6[0], addr_3857_6, addr_positional[61715:61712], addr_15428_7);

wire[31:0] addr_15429_7;

Selector_2 s15429_7(wires_3857_6[1], addr_3857_6, addr_positional[61719:61716], addr_15429_7);

wire[31:0] addr_15430_7;

Selector_2 s15430_7(wires_3857_6[2], addr_3857_6, addr_positional[61723:61720], addr_15430_7);

wire[31:0] addr_15431_7;

Selector_2 s15431_7(wires_3857_6[3], addr_3857_6, addr_positional[61727:61724], addr_15431_7);

wire[31:0] addr_15432_7;

Selector_2 s15432_7(wires_3858_6[0], addr_3858_6, addr_positional[61731:61728], addr_15432_7);

wire[31:0] addr_15433_7;

Selector_2 s15433_7(wires_3858_6[1], addr_3858_6, addr_positional[61735:61732], addr_15433_7);

wire[31:0] addr_15434_7;

Selector_2 s15434_7(wires_3858_6[2], addr_3858_6, addr_positional[61739:61736], addr_15434_7);

wire[31:0] addr_15435_7;

Selector_2 s15435_7(wires_3858_6[3], addr_3858_6, addr_positional[61743:61740], addr_15435_7);

wire[31:0] addr_15436_7;

Selector_2 s15436_7(wires_3859_6[0], addr_3859_6, addr_positional[61747:61744], addr_15436_7);

wire[31:0] addr_15437_7;

Selector_2 s15437_7(wires_3859_6[1], addr_3859_6, addr_positional[61751:61748], addr_15437_7);

wire[31:0] addr_15438_7;

Selector_2 s15438_7(wires_3859_6[2], addr_3859_6, addr_positional[61755:61752], addr_15438_7);

wire[31:0] addr_15439_7;

Selector_2 s15439_7(wires_3859_6[3], addr_3859_6, addr_positional[61759:61756], addr_15439_7);

wire[31:0] addr_15440_7;

Selector_2 s15440_7(wires_3860_6[0], addr_3860_6, addr_positional[61763:61760], addr_15440_7);

wire[31:0] addr_15441_7;

Selector_2 s15441_7(wires_3860_6[1], addr_3860_6, addr_positional[61767:61764], addr_15441_7);

wire[31:0] addr_15442_7;

Selector_2 s15442_7(wires_3860_6[2], addr_3860_6, addr_positional[61771:61768], addr_15442_7);

wire[31:0] addr_15443_7;

Selector_2 s15443_7(wires_3860_6[3], addr_3860_6, addr_positional[61775:61772], addr_15443_7);

wire[31:0] addr_15444_7;

Selector_2 s15444_7(wires_3861_6[0], addr_3861_6, addr_positional[61779:61776], addr_15444_7);

wire[31:0] addr_15445_7;

Selector_2 s15445_7(wires_3861_6[1], addr_3861_6, addr_positional[61783:61780], addr_15445_7);

wire[31:0] addr_15446_7;

Selector_2 s15446_7(wires_3861_6[2], addr_3861_6, addr_positional[61787:61784], addr_15446_7);

wire[31:0] addr_15447_7;

Selector_2 s15447_7(wires_3861_6[3], addr_3861_6, addr_positional[61791:61788], addr_15447_7);

wire[31:0] addr_15448_7;

Selector_2 s15448_7(wires_3862_6[0], addr_3862_6, addr_positional[61795:61792], addr_15448_7);

wire[31:0] addr_15449_7;

Selector_2 s15449_7(wires_3862_6[1], addr_3862_6, addr_positional[61799:61796], addr_15449_7);

wire[31:0] addr_15450_7;

Selector_2 s15450_7(wires_3862_6[2], addr_3862_6, addr_positional[61803:61800], addr_15450_7);

wire[31:0] addr_15451_7;

Selector_2 s15451_7(wires_3862_6[3], addr_3862_6, addr_positional[61807:61804], addr_15451_7);

wire[31:0] addr_15452_7;

Selector_2 s15452_7(wires_3863_6[0], addr_3863_6, addr_positional[61811:61808], addr_15452_7);

wire[31:0] addr_15453_7;

Selector_2 s15453_7(wires_3863_6[1], addr_3863_6, addr_positional[61815:61812], addr_15453_7);

wire[31:0] addr_15454_7;

Selector_2 s15454_7(wires_3863_6[2], addr_3863_6, addr_positional[61819:61816], addr_15454_7);

wire[31:0] addr_15455_7;

Selector_2 s15455_7(wires_3863_6[3], addr_3863_6, addr_positional[61823:61820], addr_15455_7);

wire[31:0] addr_15456_7;

Selector_2 s15456_7(wires_3864_6[0], addr_3864_6, addr_positional[61827:61824], addr_15456_7);

wire[31:0] addr_15457_7;

Selector_2 s15457_7(wires_3864_6[1], addr_3864_6, addr_positional[61831:61828], addr_15457_7);

wire[31:0] addr_15458_7;

Selector_2 s15458_7(wires_3864_6[2], addr_3864_6, addr_positional[61835:61832], addr_15458_7);

wire[31:0] addr_15459_7;

Selector_2 s15459_7(wires_3864_6[3], addr_3864_6, addr_positional[61839:61836], addr_15459_7);

wire[31:0] addr_15460_7;

Selector_2 s15460_7(wires_3865_6[0], addr_3865_6, addr_positional[61843:61840], addr_15460_7);

wire[31:0] addr_15461_7;

Selector_2 s15461_7(wires_3865_6[1], addr_3865_6, addr_positional[61847:61844], addr_15461_7);

wire[31:0] addr_15462_7;

Selector_2 s15462_7(wires_3865_6[2], addr_3865_6, addr_positional[61851:61848], addr_15462_7);

wire[31:0] addr_15463_7;

Selector_2 s15463_7(wires_3865_6[3], addr_3865_6, addr_positional[61855:61852], addr_15463_7);

wire[31:0] addr_15464_7;

Selector_2 s15464_7(wires_3866_6[0], addr_3866_6, addr_positional[61859:61856], addr_15464_7);

wire[31:0] addr_15465_7;

Selector_2 s15465_7(wires_3866_6[1], addr_3866_6, addr_positional[61863:61860], addr_15465_7);

wire[31:0] addr_15466_7;

Selector_2 s15466_7(wires_3866_6[2], addr_3866_6, addr_positional[61867:61864], addr_15466_7);

wire[31:0] addr_15467_7;

Selector_2 s15467_7(wires_3866_6[3], addr_3866_6, addr_positional[61871:61868], addr_15467_7);

wire[31:0] addr_15468_7;

Selector_2 s15468_7(wires_3867_6[0], addr_3867_6, addr_positional[61875:61872], addr_15468_7);

wire[31:0] addr_15469_7;

Selector_2 s15469_7(wires_3867_6[1], addr_3867_6, addr_positional[61879:61876], addr_15469_7);

wire[31:0] addr_15470_7;

Selector_2 s15470_7(wires_3867_6[2], addr_3867_6, addr_positional[61883:61880], addr_15470_7);

wire[31:0] addr_15471_7;

Selector_2 s15471_7(wires_3867_6[3], addr_3867_6, addr_positional[61887:61884], addr_15471_7);

wire[31:0] addr_15472_7;

Selector_2 s15472_7(wires_3868_6[0], addr_3868_6, addr_positional[61891:61888], addr_15472_7);

wire[31:0] addr_15473_7;

Selector_2 s15473_7(wires_3868_6[1], addr_3868_6, addr_positional[61895:61892], addr_15473_7);

wire[31:0] addr_15474_7;

Selector_2 s15474_7(wires_3868_6[2], addr_3868_6, addr_positional[61899:61896], addr_15474_7);

wire[31:0] addr_15475_7;

Selector_2 s15475_7(wires_3868_6[3], addr_3868_6, addr_positional[61903:61900], addr_15475_7);

wire[31:0] addr_15476_7;

Selector_2 s15476_7(wires_3869_6[0], addr_3869_6, addr_positional[61907:61904], addr_15476_7);

wire[31:0] addr_15477_7;

Selector_2 s15477_7(wires_3869_6[1], addr_3869_6, addr_positional[61911:61908], addr_15477_7);

wire[31:0] addr_15478_7;

Selector_2 s15478_7(wires_3869_6[2], addr_3869_6, addr_positional[61915:61912], addr_15478_7);

wire[31:0] addr_15479_7;

Selector_2 s15479_7(wires_3869_6[3], addr_3869_6, addr_positional[61919:61916], addr_15479_7);

wire[31:0] addr_15480_7;

Selector_2 s15480_7(wires_3870_6[0], addr_3870_6, addr_positional[61923:61920], addr_15480_7);

wire[31:0] addr_15481_7;

Selector_2 s15481_7(wires_3870_6[1], addr_3870_6, addr_positional[61927:61924], addr_15481_7);

wire[31:0] addr_15482_7;

Selector_2 s15482_7(wires_3870_6[2], addr_3870_6, addr_positional[61931:61928], addr_15482_7);

wire[31:0] addr_15483_7;

Selector_2 s15483_7(wires_3870_6[3], addr_3870_6, addr_positional[61935:61932], addr_15483_7);

wire[31:0] addr_15484_7;

Selector_2 s15484_7(wires_3871_6[0], addr_3871_6, addr_positional[61939:61936], addr_15484_7);

wire[31:0] addr_15485_7;

Selector_2 s15485_7(wires_3871_6[1], addr_3871_6, addr_positional[61943:61940], addr_15485_7);

wire[31:0] addr_15486_7;

Selector_2 s15486_7(wires_3871_6[2], addr_3871_6, addr_positional[61947:61944], addr_15486_7);

wire[31:0] addr_15487_7;

Selector_2 s15487_7(wires_3871_6[3], addr_3871_6, addr_positional[61951:61948], addr_15487_7);

wire[31:0] addr_15488_7;

Selector_2 s15488_7(wires_3872_6[0], addr_3872_6, addr_positional[61955:61952], addr_15488_7);

wire[31:0] addr_15489_7;

Selector_2 s15489_7(wires_3872_6[1], addr_3872_6, addr_positional[61959:61956], addr_15489_7);

wire[31:0] addr_15490_7;

Selector_2 s15490_7(wires_3872_6[2], addr_3872_6, addr_positional[61963:61960], addr_15490_7);

wire[31:0] addr_15491_7;

Selector_2 s15491_7(wires_3872_6[3], addr_3872_6, addr_positional[61967:61964], addr_15491_7);

wire[31:0] addr_15492_7;

Selector_2 s15492_7(wires_3873_6[0], addr_3873_6, addr_positional[61971:61968], addr_15492_7);

wire[31:0] addr_15493_7;

Selector_2 s15493_7(wires_3873_6[1], addr_3873_6, addr_positional[61975:61972], addr_15493_7);

wire[31:0] addr_15494_7;

Selector_2 s15494_7(wires_3873_6[2], addr_3873_6, addr_positional[61979:61976], addr_15494_7);

wire[31:0] addr_15495_7;

Selector_2 s15495_7(wires_3873_6[3], addr_3873_6, addr_positional[61983:61980], addr_15495_7);

wire[31:0] addr_15496_7;

Selector_2 s15496_7(wires_3874_6[0], addr_3874_6, addr_positional[61987:61984], addr_15496_7);

wire[31:0] addr_15497_7;

Selector_2 s15497_7(wires_3874_6[1], addr_3874_6, addr_positional[61991:61988], addr_15497_7);

wire[31:0] addr_15498_7;

Selector_2 s15498_7(wires_3874_6[2], addr_3874_6, addr_positional[61995:61992], addr_15498_7);

wire[31:0] addr_15499_7;

Selector_2 s15499_7(wires_3874_6[3], addr_3874_6, addr_positional[61999:61996], addr_15499_7);

wire[31:0] addr_15500_7;

Selector_2 s15500_7(wires_3875_6[0], addr_3875_6, addr_positional[62003:62000], addr_15500_7);

wire[31:0] addr_15501_7;

Selector_2 s15501_7(wires_3875_6[1], addr_3875_6, addr_positional[62007:62004], addr_15501_7);

wire[31:0] addr_15502_7;

Selector_2 s15502_7(wires_3875_6[2], addr_3875_6, addr_positional[62011:62008], addr_15502_7);

wire[31:0] addr_15503_7;

Selector_2 s15503_7(wires_3875_6[3], addr_3875_6, addr_positional[62015:62012], addr_15503_7);

wire[31:0] addr_15504_7;

Selector_2 s15504_7(wires_3876_6[0], addr_3876_6, addr_positional[62019:62016], addr_15504_7);

wire[31:0] addr_15505_7;

Selector_2 s15505_7(wires_3876_6[1], addr_3876_6, addr_positional[62023:62020], addr_15505_7);

wire[31:0] addr_15506_7;

Selector_2 s15506_7(wires_3876_6[2], addr_3876_6, addr_positional[62027:62024], addr_15506_7);

wire[31:0] addr_15507_7;

Selector_2 s15507_7(wires_3876_6[3], addr_3876_6, addr_positional[62031:62028], addr_15507_7);

wire[31:0] addr_15508_7;

Selector_2 s15508_7(wires_3877_6[0], addr_3877_6, addr_positional[62035:62032], addr_15508_7);

wire[31:0] addr_15509_7;

Selector_2 s15509_7(wires_3877_6[1], addr_3877_6, addr_positional[62039:62036], addr_15509_7);

wire[31:0] addr_15510_7;

Selector_2 s15510_7(wires_3877_6[2], addr_3877_6, addr_positional[62043:62040], addr_15510_7);

wire[31:0] addr_15511_7;

Selector_2 s15511_7(wires_3877_6[3], addr_3877_6, addr_positional[62047:62044], addr_15511_7);

wire[31:0] addr_15512_7;

Selector_2 s15512_7(wires_3878_6[0], addr_3878_6, addr_positional[62051:62048], addr_15512_7);

wire[31:0] addr_15513_7;

Selector_2 s15513_7(wires_3878_6[1], addr_3878_6, addr_positional[62055:62052], addr_15513_7);

wire[31:0] addr_15514_7;

Selector_2 s15514_7(wires_3878_6[2], addr_3878_6, addr_positional[62059:62056], addr_15514_7);

wire[31:0] addr_15515_7;

Selector_2 s15515_7(wires_3878_6[3], addr_3878_6, addr_positional[62063:62060], addr_15515_7);

wire[31:0] addr_15516_7;

Selector_2 s15516_7(wires_3879_6[0], addr_3879_6, addr_positional[62067:62064], addr_15516_7);

wire[31:0] addr_15517_7;

Selector_2 s15517_7(wires_3879_6[1], addr_3879_6, addr_positional[62071:62068], addr_15517_7);

wire[31:0] addr_15518_7;

Selector_2 s15518_7(wires_3879_6[2], addr_3879_6, addr_positional[62075:62072], addr_15518_7);

wire[31:0] addr_15519_7;

Selector_2 s15519_7(wires_3879_6[3], addr_3879_6, addr_positional[62079:62076], addr_15519_7);

wire[31:0] addr_15520_7;

Selector_2 s15520_7(wires_3880_6[0], addr_3880_6, addr_positional[62083:62080], addr_15520_7);

wire[31:0] addr_15521_7;

Selector_2 s15521_7(wires_3880_6[1], addr_3880_6, addr_positional[62087:62084], addr_15521_7);

wire[31:0] addr_15522_7;

Selector_2 s15522_7(wires_3880_6[2], addr_3880_6, addr_positional[62091:62088], addr_15522_7);

wire[31:0] addr_15523_7;

Selector_2 s15523_7(wires_3880_6[3], addr_3880_6, addr_positional[62095:62092], addr_15523_7);

wire[31:0] addr_15524_7;

Selector_2 s15524_7(wires_3881_6[0], addr_3881_6, addr_positional[62099:62096], addr_15524_7);

wire[31:0] addr_15525_7;

Selector_2 s15525_7(wires_3881_6[1], addr_3881_6, addr_positional[62103:62100], addr_15525_7);

wire[31:0] addr_15526_7;

Selector_2 s15526_7(wires_3881_6[2], addr_3881_6, addr_positional[62107:62104], addr_15526_7);

wire[31:0] addr_15527_7;

Selector_2 s15527_7(wires_3881_6[3], addr_3881_6, addr_positional[62111:62108], addr_15527_7);

wire[31:0] addr_15528_7;

Selector_2 s15528_7(wires_3882_6[0], addr_3882_6, addr_positional[62115:62112], addr_15528_7);

wire[31:0] addr_15529_7;

Selector_2 s15529_7(wires_3882_6[1], addr_3882_6, addr_positional[62119:62116], addr_15529_7);

wire[31:0] addr_15530_7;

Selector_2 s15530_7(wires_3882_6[2], addr_3882_6, addr_positional[62123:62120], addr_15530_7);

wire[31:0] addr_15531_7;

Selector_2 s15531_7(wires_3882_6[3], addr_3882_6, addr_positional[62127:62124], addr_15531_7);

wire[31:0] addr_15532_7;

Selector_2 s15532_7(wires_3883_6[0], addr_3883_6, addr_positional[62131:62128], addr_15532_7);

wire[31:0] addr_15533_7;

Selector_2 s15533_7(wires_3883_6[1], addr_3883_6, addr_positional[62135:62132], addr_15533_7);

wire[31:0] addr_15534_7;

Selector_2 s15534_7(wires_3883_6[2], addr_3883_6, addr_positional[62139:62136], addr_15534_7);

wire[31:0] addr_15535_7;

Selector_2 s15535_7(wires_3883_6[3], addr_3883_6, addr_positional[62143:62140], addr_15535_7);

wire[31:0] addr_15536_7;

Selector_2 s15536_7(wires_3884_6[0], addr_3884_6, addr_positional[62147:62144], addr_15536_7);

wire[31:0] addr_15537_7;

Selector_2 s15537_7(wires_3884_6[1], addr_3884_6, addr_positional[62151:62148], addr_15537_7);

wire[31:0] addr_15538_7;

Selector_2 s15538_7(wires_3884_6[2], addr_3884_6, addr_positional[62155:62152], addr_15538_7);

wire[31:0] addr_15539_7;

Selector_2 s15539_7(wires_3884_6[3], addr_3884_6, addr_positional[62159:62156], addr_15539_7);

wire[31:0] addr_15540_7;

Selector_2 s15540_7(wires_3885_6[0], addr_3885_6, addr_positional[62163:62160], addr_15540_7);

wire[31:0] addr_15541_7;

Selector_2 s15541_7(wires_3885_6[1], addr_3885_6, addr_positional[62167:62164], addr_15541_7);

wire[31:0] addr_15542_7;

Selector_2 s15542_7(wires_3885_6[2], addr_3885_6, addr_positional[62171:62168], addr_15542_7);

wire[31:0] addr_15543_7;

Selector_2 s15543_7(wires_3885_6[3], addr_3885_6, addr_positional[62175:62172], addr_15543_7);

wire[31:0] addr_15544_7;

Selector_2 s15544_7(wires_3886_6[0], addr_3886_6, addr_positional[62179:62176], addr_15544_7);

wire[31:0] addr_15545_7;

Selector_2 s15545_7(wires_3886_6[1], addr_3886_6, addr_positional[62183:62180], addr_15545_7);

wire[31:0] addr_15546_7;

Selector_2 s15546_7(wires_3886_6[2], addr_3886_6, addr_positional[62187:62184], addr_15546_7);

wire[31:0] addr_15547_7;

Selector_2 s15547_7(wires_3886_6[3], addr_3886_6, addr_positional[62191:62188], addr_15547_7);

wire[31:0] addr_15548_7;

Selector_2 s15548_7(wires_3887_6[0], addr_3887_6, addr_positional[62195:62192], addr_15548_7);

wire[31:0] addr_15549_7;

Selector_2 s15549_7(wires_3887_6[1], addr_3887_6, addr_positional[62199:62196], addr_15549_7);

wire[31:0] addr_15550_7;

Selector_2 s15550_7(wires_3887_6[2], addr_3887_6, addr_positional[62203:62200], addr_15550_7);

wire[31:0] addr_15551_7;

Selector_2 s15551_7(wires_3887_6[3], addr_3887_6, addr_positional[62207:62204], addr_15551_7);

wire[31:0] addr_15552_7;

Selector_2 s15552_7(wires_3888_6[0], addr_3888_6, addr_positional[62211:62208], addr_15552_7);

wire[31:0] addr_15553_7;

Selector_2 s15553_7(wires_3888_6[1], addr_3888_6, addr_positional[62215:62212], addr_15553_7);

wire[31:0] addr_15554_7;

Selector_2 s15554_7(wires_3888_6[2], addr_3888_6, addr_positional[62219:62216], addr_15554_7);

wire[31:0] addr_15555_7;

Selector_2 s15555_7(wires_3888_6[3], addr_3888_6, addr_positional[62223:62220], addr_15555_7);

wire[31:0] addr_15556_7;

Selector_2 s15556_7(wires_3889_6[0], addr_3889_6, addr_positional[62227:62224], addr_15556_7);

wire[31:0] addr_15557_7;

Selector_2 s15557_7(wires_3889_6[1], addr_3889_6, addr_positional[62231:62228], addr_15557_7);

wire[31:0] addr_15558_7;

Selector_2 s15558_7(wires_3889_6[2], addr_3889_6, addr_positional[62235:62232], addr_15558_7);

wire[31:0] addr_15559_7;

Selector_2 s15559_7(wires_3889_6[3], addr_3889_6, addr_positional[62239:62236], addr_15559_7);

wire[31:0] addr_15560_7;

Selector_2 s15560_7(wires_3890_6[0], addr_3890_6, addr_positional[62243:62240], addr_15560_7);

wire[31:0] addr_15561_7;

Selector_2 s15561_7(wires_3890_6[1], addr_3890_6, addr_positional[62247:62244], addr_15561_7);

wire[31:0] addr_15562_7;

Selector_2 s15562_7(wires_3890_6[2], addr_3890_6, addr_positional[62251:62248], addr_15562_7);

wire[31:0] addr_15563_7;

Selector_2 s15563_7(wires_3890_6[3], addr_3890_6, addr_positional[62255:62252], addr_15563_7);

wire[31:0] addr_15564_7;

Selector_2 s15564_7(wires_3891_6[0], addr_3891_6, addr_positional[62259:62256], addr_15564_7);

wire[31:0] addr_15565_7;

Selector_2 s15565_7(wires_3891_6[1], addr_3891_6, addr_positional[62263:62260], addr_15565_7);

wire[31:0] addr_15566_7;

Selector_2 s15566_7(wires_3891_6[2], addr_3891_6, addr_positional[62267:62264], addr_15566_7);

wire[31:0] addr_15567_7;

Selector_2 s15567_7(wires_3891_6[3], addr_3891_6, addr_positional[62271:62268], addr_15567_7);

wire[31:0] addr_15568_7;

Selector_2 s15568_7(wires_3892_6[0], addr_3892_6, addr_positional[62275:62272], addr_15568_7);

wire[31:0] addr_15569_7;

Selector_2 s15569_7(wires_3892_6[1], addr_3892_6, addr_positional[62279:62276], addr_15569_7);

wire[31:0] addr_15570_7;

Selector_2 s15570_7(wires_3892_6[2], addr_3892_6, addr_positional[62283:62280], addr_15570_7);

wire[31:0] addr_15571_7;

Selector_2 s15571_7(wires_3892_6[3], addr_3892_6, addr_positional[62287:62284], addr_15571_7);

wire[31:0] addr_15572_7;

Selector_2 s15572_7(wires_3893_6[0], addr_3893_6, addr_positional[62291:62288], addr_15572_7);

wire[31:0] addr_15573_7;

Selector_2 s15573_7(wires_3893_6[1], addr_3893_6, addr_positional[62295:62292], addr_15573_7);

wire[31:0] addr_15574_7;

Selector_2 s15574_7(wires_3893_6[2], addr_3893_6, addr_positional[62299:62296], addr_15574_7);

wire[31:0] addr_15575_7;

Selector_2 s15575_7(wires_3893_6[3], addr_3893_6, addr_positional[62303:62300], addr_15575_7);

wire[31:0] addr_15576_7;

Selector_2 s15576_7(wires_3894_6[0], addr_3894_6, addr_positional[62307:62304], addr_15576_7);

wire[31:0] addr_15577_7;

Selector_2 s15577_7(wires_3894_6[1], addr_3894_6, addr_positional[62311:62308], addr_15577_7);

wire[31:0] addr_15578_7;

Selector_2 s15578_7(wires_3894_6[2], addr_3894_6, addr_positional[62315:62312], addr_15578_7);

wire[31:0] addr_15579_7;

Selector_2 s15579_7(wires_3894_6[3], addr_3894_6, addr_positional[62319:62316], addr_15579_7);

wire[31:0] addr_15580_7;

Selector_2 s15580_7(wires_3895_6[0], addr_3895_6, addr_positional[62323:62320], addr_15580_7);

wire[31:0] addr_15581_7;

Selector_2 s15581_7(wires_3895_6[1], addr_3895_6, addr_positional[62327:62324], addr_15581_7);

wire[31:0] addr_15582_7;

Selector_2 s15582_7(wires_3895_6[2], addr_3895_6, addr_positional[62331:62328], addr_15582_7);

wire[31:0] addr_15583_7;

Selector_2 s15583_7(wires_3895_6[3], addr_3895_6, addr_positional[62335:62332], addr_15583_7);

wire[31:0] addr_15584_7;

Selector_2 s15584_7(wires_3896_6[0], addr_3896_6, addr_positional[62339:62336], addr_15584_7);

wire[31:0] addr_15585_7;

Selector_2 s15585_7(wires_3896_6[1], addr_3896_6, addr_positional[62343:62340], addr_15585_7);

wire[31:0] addr_15586_7;

Selector_2 s15586_7(wires_3896_6[2], addr_3896_6, addr_positional[62347:62344], addr_15586_7);

wire[31:0] addr_15587_7;

Selector_2 s15587_7(wires_3896_6[3], addr_3896_6, addr_positional[62351:62348], addr_15587_7);

wire[31:0] addr_15588_7;

Selector_2 s15588_7(wires_3897_6[0], addr_3897_6, addr_positional[62355:62352], addr_15588_7);

wire[31:0] addr_15589_7;

Selector_2 s15589_7(wires_3897_6[1], addr_3897_6, addr_positional[62359:62356], addr_15589_7);

wire[31:0] addr_15590_7;

Selector_2 s15590_7(wires_3897_6[2], addr_3897_6, addr_positional[62363:62360], addr_15590_7);

wire[31:0] addr_15591_7;

Selector_2 s15591_7(wires_3897_6[3], addr_3897_6, addr_positional[62367:62364], addr_15591_7);

wire[31:0] addr_15592_7;

Selector_2 s15592_7(wires_3898_6[0], addr_3898_6, addr_positional[62371:62368], addr_15592_7);

wire[31:0] addr_15593_7;

Selector_2 s15593_7(wires_3898_6[1], addr_3898_6, addr_positional[62375:62372], addr_15593_7);

wire[31:0] addr_15594_7;

Selector_2 s15594_7(wires_3898_6[2], addr_3898_6, addr_positional[62379:62376], addr_15594_7);

wire[31:0] addr_15595_7;

Selector_2 s15595_7(wires_3898_6[3], addr_3898_6, addr_positional[62383:62380], addr_15595_7);

wire[31:0] addr_15596_7;

Selector_2 s15596_7(wires_3899_6[0], addr_3899_6, addr_positional[62387:62384], addr_15596_7);

wire[31:0] addr_15597_7;

Selector_2 s15597_7(wires_3899_6[1], addr_3899_6, addr_positional[62391:62388], addr_15597_7);

wire[31:0] addr_15598_7;

Selector_2 s15598_7(wires_3899_6[2], addr_3899_6, addr_positional[62395:62392], addr_15598_7);

wire[31:0] addr_15599_7;

Selector_2 s15599_7(wires_3899_6[3], addr_3899_6, addr_positional[62399:62396], addr_15599_7);

wire[31:0] addr_15600_7;

Selector_2 s15600_7(wires_3900_6[0], addr_3900_6, addr_positional[62403:62400], addr_15600_7);

wire[31:0] addr_15601_7;

Selector_2 s15601_7(wires_3900_6[1], addr_3900_6, addr_positional[62407:62404], addr_15601_7);

wire[31:0] addr_15602_7;

Selector_2 s15602_7(wires_3900_6[2], addr_3900_6, addr_positional[62411:62408], addr_15602_7);

wire[31:0] addr_15603_7;

Selector_2 s15603_7(wires_3900_6[3], addr_3900_6, addr_positional[62415:62412], addr_15603_7);

wire[31:0] addr_15604_7;

Selector_2 s15604_7(wires_3901_6[0], addr_3901_6, addr_positional[62419:62416], addr_15604_7);

wire[31:0] addr_15605_7;

Selector_2 s15605_7(wires_3901_6[1], addr_3901_6, addr_positional[62423:62420], addr_15605_7);

wire[31:0] addr_15606_7;

Selector_2 s15606_7(wires_3901_6[2], addr_3901_6, addr_positional[62427:62424], addr_15606_7);

wire[31:0] addr_15607_7;

Selector_2 s15607_7(wires_3901_6[3], addr_3901_6, addr_positional[62431:62428], addr_15607_7);

wire[31:0] addr_15608_7;

Selector_2 s15608_7(wires_3902_6[0], addr_3902_6, addr_positional[62435:62432], addr_15608_7);

wire[31:0] addr_15609_7;

Selector_2 s15609_7(wires_3902_6[1], addr_3902_6, addr_positional[62439:62436], addr_15609_7);

wire[31:0] addr_15610_7;

Selector_2 s15610_7(wires_3902_6[2], addr_3902_6, addr_positional[62443:62440], addr_15610_7);

wire[31:0] addr_15611_7;

Selector_2 s15611_7(wires_3902_6[3], addr_3902_6, addr_positional[62447:62444], addr_15611_7);

wire[31:0] addr_15612_7;

Selector_2 s15612_7(wires_3903_6[0], addr_3903_6, addr_positional[62451:62448], addr_15612_7);

wire[31:0] addr_15613_7;

Selector_2 s15613_7(wires_3903_6[1], addr_3903_6, addr_positional[62455:62452], addr_15613_7);

wire[31:0] addr_15614_7;

Selector_2 s15614_7(wires_3903_6[2], addr_3903_6, addr_positional[62459:62456], addr_15614_7);

wire[31:0] addr_15615_7;

Selector_2 s15615_7(wires_3903_6[3], addr_3903_6, addr_positional[62463:62460], addr_15615_7);

wire[31:0] addr_15616_7;

Selector_2 s15616_7(wires_3904_6[0], addr_3904_6, addr_positional[62467:62464], addr_15616_7);

wire[31:0] addr_15617_7;

Selector_2 s15617_7(wires_3904_6[1], addr_3904_6, addr_positional[62471:62468], addr_15617_7);

wire[31:0] addr_15618_7;

Selector_2 s15618_7(wires_3904_6[2], addr_3904_6, addr_positional[62475:62472], addr_15618_7);

wire[31:0] addr_15619_7;

Selector_2 s15619_7(wires_3904_6[3], addr_3904_6, addr_positional[62479:62476], addr_15619_7);

wire[31:0] addr_15620_7;

Selector_2 s15620_7(wires_3905_6[0], addr_3905_6, addr_positional[62483:62480], addr_15620_7);

wire[31:0] addr_15621_7;

Selector_2 s15621_7(wires_3905_6[1], addr_3905_6, addr_positional[62487:62484], addr_15621_7);

wire[31:0] addr_15622_7;

Selector_2 s15622_7(wires_3905_6[2], addr_3905_6, addr_positional[62491:62488], addr_15622_7);

wire[31:0] addr_15623_7;

Selector_2 s15623_7(wires_3905_6[3], addr_3905_6, addr_positional[62495:62492], addr_15623_7);

wire[31:0] addr_15624_7;

Selector_2 s15624_7(wires_3906_6[0], addr_3906_6, addr_positional[62499:62496], addr_15624_7);

wire[31:0] addr_15625_7;

Selector_2 s15625_7(wires_3906_6[1], addr_3906_6, addr_positional[62503:62500], addr_15625_7);

wire[31:0] addr_15626_7;

Selector_2 s15626_7(wires_3906_6[2], addr_3906_6, addr_positional[62507:62504], addr_15626_7);

wire[31:0] addr_15627_7;

Selector_2 s15627_7(wires_3906_6[3], addr_3906_6, addr_positional[62511:62508], addr_15627_7);

wire[31:0] addr_15628_7;

Selector_2 s15628_7(wires_3907_6[0], addr_3907_6, addr_positional[62515:62512], addr_15628_7);

wire[31:0] addr_15629_7;

Selector_2 s15629_7(wires_3907_6[1], addr_3907_6, addr_positional[62519:62516], addr_15629_7);

wire[31:0] addr_15630_7;

Selector_2 s15630_7(wires_3907_6[2], addr_3907_6, addr_positional[62523:62520], addr_15630_7);

wire[31:0] addr_15631_7;

Selector_2 s15631_7(wires_3907_6[3], addr_3907_6, addr_positional[62527:62524], addr_15631_7);

wire[31:0] addr_15632_7;

Selector_2 s15632_7(wires_3908_6[0], addr_3908_6, addr_positional[62531:62528], addr_15632_7);

wire[31:0] addr_15633_7;

Selector_2 s15633_7(wires_3908_6[1], addr_3908_6, addr_positional[62535:62532], addr_15633_7);

wire[31:0] addr_15634_7;

Selector_2 s15634_7(wires_3908_6[2], addr_3908_6, addr_positional[62539:62536], addr_15634_7);

wire[31:0] addr_15635_7;

Selector_2 s15635_7(wires_3908_6[3], addr_3908_6, addr_positional[62543:62540], addr_15635_7);

wire[31:0] addr_15636_7;

Selector_2 s15636_7(wires_3909_6[0], addr_3909_6, addr_positional[62547:62544], addr_15636_7);

wire[31:0] addr_15637_7;

Selector_2 s15637_7(wires_3909_6[1], addr_3909_6, addr_positional[62551:62548], addr_15637_7);

wire[31:0] addr_15638_7;

Selector_2 s15638_7(wires_3909_6[2], addr_3909_6, addr_positional[62555:62552], addr_15638_7);

wire[31:0] addr_15639_7;

Selector_2 s15639_7(wires_3909_6[3], addr_3909_6, addr_positional[62559:62556], addr_15639_7);

wire[31:0] addr_15640_7;

Selector_2 s15640_7(wires_3910_6[0], addr_3910_6, addr_positional[62563:62560], addr_15640_7);

wire[31:0] addr_15641_7;

Selector_2 s15641_7(wires_3910_6[1], addr_3910_6, addr_positional[62567:62564], addr_15641_7);

wire[31:0] addr_15642_7;

Selector_2 s15642_7(wires_3910_6[2], addr_3910_6, addr_positional[62571:62568], addr_15642_7);

wire[31:0] addr_15643_7;

Selector_2 s15643_7(wires_3910_6[3], addr_3910_6, addr_positional[62575:62572], addr_15643_7);

wire[31:0] addr_15644_7;

Selector_2 s15644_7(wires_3911_6[0], addr_3911_6, addr_positional[62579:62576], addr_15644_7);

wire[31:0] addr_15645_7;

Selector_2 s15645_7(wires_3911_6[1], addr_3911_6, addr_positional[62583:62580], addr_15645_7);

wire[31:0] addr_15646_7;

Selector_2 s15646_7(wires_3911_6[2], addr_3911_6, addr_positional[62587:62584], addr_15646_7);

wire[31:0] addr_15647_7;

Selector_2 s15647_7(wires_3911_6[3], addr_3911_6, addr_positional[62591:62588], addr_15647_7);

wire[31:0] addr_15648_7;

Selector_2 s15648_7(wires_3912_6[0], addr_3912_6, addr_positional[62595:62592], addr_15648_7);

wire[31:0] addr_15649_7;

Selector_2 s15649_7(wires_3912_6[1], addr_3912_6, addr_positional[62599:62596], addr_15649_7);

wire[31:0] addr_15650_7;

Selector_2 s15650_7(wires_3912_6[2], addr_3912_6, addr_positional[62603:62600], addr_15650_7);

wire[31:0] addr_15651_7;

Selector_2 s15651_7(wires_3912_6[3], addr_3912_6, addr_positional[62607:62604], addr_15651_7);

wire[31:0] addr_15652_7;

Selector_2 s15652_7(wires_3913_6[0], addr_3913_6, addr_positional[62611:62608], addr_15652_7);

wire[31:0] addr_15653_7;

Selector_2 s15653_7(wires_3913_6[1], addr_3913_6, addr_positional[62615:62612], addr_15653_7);

wire[31:0] addr_15654_7;

Selector_2 s15654_7(wires_3913_6[2], addr_3913_6, addr_positional[62619:62616], addr_15654_7);

wire[31:0] addr_15655_7;

Selector_2 s15655_7(wires_3913_6[3], addr_3913_6, addr_positional[62623:62620], addr_15655_7);

wire[31:0] addr_15656_7;

Selector_2 s15656_7(wires_3914_6[0], addr_3914_6, addr_positional[62627:62624], addr_15656_7);

wire[31:0] addr_15657_7;

Selector_2 s15657_7(wires_3914_6[1], addr_3914_6, addr_positional[62631:62628], addr_15657_7);

wire[31:0] addr_15658_7;

Selector_2 s15658_7(wires_3914_6[2], addr_3914_6, addr_positional[62635:62632], addr_15658_7);

wire[31:0] addr_15659_7;

Selector_2 s15659_7(wires_3914_6[3], addr_3914_6, addr_positional[62639:62636], addr_15659_7);

wire[31:0] addr_15660_7;

Selector_2 s15660_7(wires_3915_6[0], addr_3915_6, addr_positional[62643:62640], addr_15660_7);

wire[31:0] addr_15661_7;

Selector_2 s15661_7(wires_3915_6[1], addr_3915_6, addr_positional[62647:62644], addr_15661_7);

wire[31:0] addr_15662_7;

Selector_2 s15662_7(wires_3915_6[2], addr_3915_6, addr_positional[62651:62648], addr_15662_7);

wire[31:0] addr_15663_7;

Selector_2 s15663_7(wires_3915_6[3], addr_3915_6, addr_positional[62655:62652], addr_15663_7);

wire[31:0] addr_15664_7;

Selector_2 s15664_7(wires_3916_6[0], addr_3916_6, addr_positional[62659:62656], addr_15664_7);

wire[31:0] addr_15665_7;

Selector_2 s15665_7(wires_3916_6[1], addr_3916_6, addr_positional[62663:62660], addr_15665_7);

wire[31:0] addr_15666_7;

Selector_2 s15666_7(wires_3916_6[2], addr_3916_6, addr_positional[62667:62664], addr_15666_7);

wire[31:0] addr_15667_7;

Selector_2 s15667_7(wires_3916_6[3], addr_3916_6, addr_positional[62671:62668], addr_15667_7);

wire[31:0] addr_15668_7;

Selector_2 s15668_7(wires_3917_6[0], addr_3917_6, addr_positional[62675:62672], addr_15668_7);

wire[31:0] addr_15669_7;

Selector_2 s15669_7(wires_3917_6[1], addr_3917_6, addr_positional[62679:62676], addr_15669_7);

wire[31:0] addr_15670_7;

Selector_2 s15670_7(wires_3917_6[2], addr_3917_6, addr_positional[62683:62680], addr_15670_7);

wire[31:0] addr_15671_7;

Selector_2 s15671_7(wires_3917_6[3], addr_3917_6, addr_positional[62687:62684], addr_15671_7);

wire[31:0] addr_15672_7;

Selector_2 s15672_7(wires_3918_6[0], addr_3918_6, addr_positional[62691:62688], addr_15672_7);

wire[31:0] addr_15673_7;

Selector_2 s15673_7(wires_3918_6[1], addr_3918_6, addr_positional[62695:62692], addr_15673_7);

wire[31:0] addr_15674_7;

Selector_2 s15674_7(wires_3918_6[2], addr_3918_6, addr_positional[62699:62696], addr_15674_7);

wire[31:0] addr_15675_7;

Selector_2 s15675_7(wires_3918_6[3], addr_3918_6, addr_positional[62703:62700], addr_15675_7);

wire[31:0] addr_15676_7;

Selector_2 s15676_7(wires_3919_6[0], addr_3919_6, addr_positional[62707:62704], addr_15676_7);

wire[31:0] addr_15677_7;

Selector_2 s15677_7(wires_3919_6[1], addr_3919_6, addr_positional[62711:62708], addr_15677_7);

wire[31:0] addr_15678_7;

Selector_2 s15678_7(wires_3919_6[2], addr_3919_6, addr_positional[62715:62712], addr_15678_7);

wire[31:0] addr_15679_7;

Selector_2 s15679_7(wires_3919_6[3], addr_3919_6, addr_positional[62719:62716], addr_15679_7);

wire[31:0] addr_15680_7;

Selector_2 s15680_7(wires_3920_6[0], addr_3920_6, addr_positional[62723:62720], addr_15680_7);

wire[31:0] addr_15681_7;

Selector_2 s15681_7(wires_3920_6[1], addr_3920_6, addr_positional[62727:62724], addr_15681_7);

wire[31:0] addr_15682_7;

Selector_2 s15682_7(wires_3920_6[2], addr_3920_6, addr_positional[62731:62728], addr_15682_7);

wire[31:0] addr_15683_7;

Selector_2 s15683_7(wires_3920_6[3], addr_3920_6, addr_positional[62735:62732], addr_15683_7);

wire[31:0] addr_15684_7;

Selector_2 s15684_7(wires_3921_6[0], addr_3921_6, addr_positional[62739:62736], addr_15684_7);

wire[31:0] addr_15685_7;

Selector_2 s15685_7(wires_3921_6[1], addr_3921_6, addr_positional[62743:62740], addr_15685_7);

wire[31:0] addr_15686_7;

Selector_2 s15686_7(wires_3921_6[2], addr_3921_6, addr_positional[62747:62744], addr_15686_7);

wire[31:0] addr_15687_7;

Selector_2 s15687_7(wires_3921_6[3], addr_3921_6, addr_positional[62751:62748], addr_15687_7);

wire[31:0] addr_15688_7;

Selector_2 s15688_7(wires_3922_6[0], addr_3922_6, addr_positional[62755:62752], addr_15688_7);

wire[31:0] addr_15689_7;

Selector_2 s15689_7(wires_3922_6[1], addr_3922_6, addr_positional[62759:62756], addr_15689_7);

wire[31:0] addr_15690_7;

Selector_2 s15690_7(wires_3922_6[2], addr_3922_6, addr_positional[62763:62760], addr_15690_7);

wire[31:0] addr_15691_7;

Selector_2 s15691_7(wires_3922_6[3], addr_3922_6, addr_positional[62767:62764], addr_15691_7);

wire[31:0] addr_15692_7;

Selector_2 s15692_7(wires_3923_6[0], addr_3923_6, addr_positional[62771:62768], addr_15692_7);

wire[31:0] addr_15693_7;

Selector_2 s15693_7(wires_3923_6[1], addr_3923_6, addr_positional[62775:62772], addr_15693_7);

wire[31:0] addr_15694_7;

Selector_2 s15694_7(wires_3923_6[2], addr_3923_6, addr_positional[62779:62776], addr_15694_7);

wire[31:0] addr_15695_7;

Selector_2 s15695_7(wires_3923_6[3], addr_3923_6, addr_positional[62783:62780], addr_15695_7);

wire[31:0] addr_15696_7;

Selector_2 s15696_7(wires_3924_6[0], addr_3924_6, addr_positional[62787:62784], addr_15696_7);

wire[31:0] addr_15697_7;

Selector_2 s15697_7(wires_3924_6[1], addr_3924_6, addr_positional[62791:62788], addr_15697_7);

wire[31:0] addr_15698_7;

Selector_2 s15698_7(wires_3924_6[2], addr_3924_6, addr_positional[62795:62792], addr_15698_7);

wire[31:0] addr_15699_7;

Selector_2 s15699_7(wires_3924_6[3], addr_3924_6, addr_positional[62799:62796], addr_15699_7);

wire[31:0] addr_15700_7;

Selector_2 s15700_7(wires_3925_6[0], addr_3925_6, addr_positional[62803:62800], addr_15700_7);

wire[31:0] addr_15701_7;

Selector_2 s15701_7(wires_3925_6[1], addr_3925_6, addr_positional[62807:62804], addr_15701_7);

wire[31:0] addr_15702_7;

Selector_2 s15702_7(wires_3925_6[2], addr_3925_6, addr_positional[62811:62808], addr_15702_7);

wire[31:0] addr_15703_7;

Selector_2 s15703_7(wires_3925_6[3], addr_3925_6, addr_positional[62815:62812], addr_15703_7);

wire[31:0] addr_15704_7;

Selector_2 s15704_7(wires_3926_6[0], addr_3926_6, addr_positional[62819:62816], addr_15704_7);

wire[31:0] addr_15705_7;

Selector_2 s15705_7(wires_3926_6[1], addr_3926_6, addr_positional[62823:62820], addr_15705_7);

wire[31:0] addr_15706_7;

Selector_2 s15706_7(wires_3926_6[2], addr_3926_6, addr_positional[62827:62824], addr_15706_7);

wire[31:0] addr_15707_7;

Selector_2 s15707_7(wires_3926_6[3], addr_3926_6, addr_positional[62831:62828], addr_15707_7);

wire[31:0] addr_15708_7;

Selector_2 s15708_7(wires_3927_6[0], addr_3927_6, addr_positional[62835:62832], addr_15708_7);

wire[31:0] addr_15709_7;

Selector_2 s15709_7(wires_3927_6[1], addr_3927_6, addr_positional[62839:62836], addr_15709_7);

wire[31:0] addr_15710_7;

Selector_2 s15710_7(wires_3927_6[2], addr_3927_6, addr_positional[62843:62840], addr_15710_7);

wire[31:0] addr_15711_7;

Selector_2 s15711_7(wires_3927_6[3], addr_3927_6, addr_positional[62847:62844], addr_15711_7);

wire[31:0] addr_15712_7;

Selector_2 s15712_7(wires_3928_6[0], addr_3928_6, addr_positional[62851:62848], addr_15712_7);

wire[31:0] addr_15713_7;

Selector_2 s15713_7(wires_3928_6[1], addr_3928_6, addr_positional[62855:62852], addr_15713_7);

wire[31:0] addr_15714_7;

Selector_2 s15714_7(wires_3928_6[2], addr_3928_6, addr_positional[62859:62856], addr_15714_7);

wire[31:0] addr_15715_7;

Selector_2 s15715_7(wires_3928_6[3], addr_3928_6, addr_positional[62863:62860], addr_15715_7);

wire[31:0] addr_15716_7;

Selector_2 s15716_7(wires_3929_6[0], addr_3929_6, addr_positional[62867:62864], addr_15716_7);

wire[31:0] addr_15717_7;

Selector_2 s15717_7(wires_3929_6[1], addr_3929_6, addr_positional[62871:62868], addr_15717_7);

wire[31:0] addr_15718_7;

Selector_2 s15718_7(wires_3929_6[2], addr_3929_6, addr_positional[62875:62872], addr_15718_7);

wire[31:0] addr_15719_7;

Selector_2 s15719_7(wires_3929_6[3], addr_3929_6, addr_positional[62879:62876], addr_15719_7);

wire[31:0] addr_15720_7;

Selector_2 s15720_7(wires_3930_6[0], addr_3930_6, addr_positional[62883:62880], addr_15720_7);

wire[31:0] addr_15721_7;

Selector_2 s15721_7(wires_3930_6[1], addr_3930_6, addr_positional[62887:62884], addr_15721_7);

wire[31:0] addr_15722_7;

Selector_2 s15722_7(wires_3930_6[2], addr_3930_6, addr_positional[62891:62888], addr_15722_7);

wire[31:0] addr_15723_7;

Selector_2 s15723_7(wires_3930_6[3], addr_3930_6, addr_positional[62895:62892], addr_15723_7);

wire[31:0] addr_15724_7;

Selector_2 s15724_7(wires_3931_6[0], addr_3931_6, addr_positional[62899:62896], addr_15724_7);

wire[31:0] addr_15725_7;

Selector_2 s15725_7(wires_3931_6[1], addr_3931_6, addr_positional[62903:62900], addr_15725_7);

wire[31:0] addr_15726_7;

Selector_2 s15726_7(wires_3931_6[2], addr_3931_6, addr_positional[62907:62904], addr_15726_7);

wire[31:0] addr_15727_7;

Selector_2 s15727_7(wires_3931_6[3], addr_3931_6, addr_positional[62911:62908], addr_15727_7);

wire[31:0] addr_15728_7;

Selector_2 s15728_7(wires_3932_6[0], addr_3932_6, addr_positional[62915:62912], addr_15728_7);

wire[31:0] addr_15729_7;

Selector_2 s15729_7(wires_3932_6[1], addr_3932_6, addr_positional[62919:62916], addr_15729_7);

wire[31:0] addr_15730_7;

Selector_2 s15730_7(wires_3932_6[2], addr_3932_6, addr_positional[62923:62920], addr_15730_7);

wire[31:0] addr_15731_7;

Selector_2 s15731_7(wires_3932_6[3], addr_3932_6, addr_positional[62927:62924], addr_15731_7);

wire[31:0] addr_15732_7;

Selector_2 s15732_7(wires_3933_6[0], addr_3933_6, addr_positional[62931:62928], addr_15732_7);

wire[31:0] addr_15733_7;

Selector_2 s15733_7(wires_3933_6[1], addr_3933_6, addr_positional[62935:62932], addr_15733_7);

wire[31:0] addr_15734_7;

Selector_2 s15734_7(wires_3933_6[2], addr_3933_6, addr_positional[62939:62936], addr_15734_7);

wire[31:0] addr_15735_7;

Selector_2 s15735_7(wires_3933_6[3], addr_3933_6, addr_positional[62943:62940], addr_15735_7);

wire[31:0] addr_15736_7;

Selector_2 s15736_7(wires_3934_6[0], addr_3934_6, addr_positional[62947:62944], addr_15736_7);

wire[31:0] addr_15737_7;

Selector_2 s15737_7(wires_3934_6[1], addr_3934_6, addr_positional[62951:62948], addr_15737_7);

wire[31:0] addr_15738_7;

Selector_2 s15738_7(wires_3934_6[2], addr_3934_6, addr_positional[62955:62952], addr_15738_7);

wire[31:0] addr_15739_7;

Selector_2 s15739_7(wires_3934_6[3], addr_3934_6, addr_positional[62959:62956], addr_15739_7);

wire[31:0] addr_15740_7;

Selector_2 s15740_7(wires_3935_6[0], addr_3935_6, addr_positional[62963:62960], addr_15740_7);

wire[31:0] addr_15741_7;

Selector_2 s15741_7(wires_3935_6[1], addr_3935_6, addr_positional[62967:62964], addr_15741_7);

wire[31:0] addr_15742_7;

Selector_2 s15742_7(wires_3935_6[2], addr_3935_6, addr_positional[62971:62968], addr_15742_7);

wire[31:0] addr_15743_7;

Selector_2 s15743_7(wires_3935_6[3], addr_3935_6, addr_positional[62975:62972], addr_15743_7);

wire[31:0] addr_15744_7;

Selector_2 s15744_7(wires_3936_6[0], addr_3936_6, addr_positional[62979:62976], addr_15744_7);

wire[31:0] addr_15745_7;

Selector_2 s15745_7(wires_3936_6[1], addr_3936_6, addr_positional[62983:62980], addr_15745_7);

wire[31:0] addr_15746_7;

Selector_2 s15746_7(wires_3936_6[2], addr_3936_6, addr_positional[62987:62984], addr_15746_7);

wire[31:0] addr_15747_7;

Selector_2 s15747_7(wires_3936_6[3], addr_3936_6, addr_positional[62991:62988], addr_15747_7);

wire[31:0] addr_15748_7;

Selector_2 s15748_7(wires_3937_6[0], addr_3937_6, addr_positional[62995:62992], addr_15748_7);

wire[31:0] addr_15749_7;

Selector_2 s15749_7(wires_3937_6[1], addr_3937_6, addr_positional[62999:62996], addr_15749_7);

wire[31:0] addr_15750_7;

Selector_2 s15750_7(wires_3937_6[2], addr_3937_6, addr_positional[63003:63000], addr_15750_7);

wire[31:0] addr_15751_7;

Selector_2 s15751_7(wires_3937_6[3], addr_3937_6, addr_positional[63007:63004], addr_15751_7);

wire[31:0] addr_15752_7;

Selector_2 s15752_7(wires_3938_6[0], addr_3938_6, addr_positional[63011:63008], addr_15752_7);

wire[31:0] addr_15753_7;

Selector_2 s15753_7(wires_3938_6[1], addr_3938_6, addr_positional[63015:63012], addr_15753_7);

wire[31:0] addr_15754_7;

Selector_2 s15754_7(wires_3938_6[2], addr_3938_6, addr_positional[63019:63016], addr_15754_7);

wire[31:0] addr_15755_7;

Selector_2 s15755_7(wires_3938_6[3], addr_3938_6, addr_positional[63023:63020], addr_15755_7);

wire[31:0] addr_15756_7;

Selector_2 s15756_7(wires_3939_6[0], addr_3939_6, addr_positional[63027:63024], addr_15756_7);

wire[31:0] addr_15757_7;

Selector_2 s15757_7(wires_3939_6[1], addr_3939_6, addr_positional[63031:63028], addr_15757_7);

wire[31:0] addr_15758_7;

Selector_2 s15758_7(wires_3939_6[2], addr_3939_6, addr_positional[63035:63032], addr_15758_7);

wire[31:0] addr_15759_7;

Selector_2 s15759_7(wires_3939_6[3], addr_3939_6, addr_positional[63039:63036], addr_15759_7);

wire[31:0] addr_15760_7;

Selector_2 s15760_7(wires_3940_6[0], addr_3940_6, addr_positional[63043:63040], addr_15760_7);

wire[31:0] addr_15761_7;

Selector_2 s15761_7(wires_3940_6[1], addr_3940_6, addr_positional[63047:63044], addr_15761_7);

wire[31:0] addr_15762_7;

Selector_2 s15762_7(wires_3940_6[2], addr_3940_6, addr_positional[63051:63048], addr_15762_7);

wire[31:0] addr_15763_7;

Selector_2 s15763_7(wires_3940_6[3], addr_3940_6, addr_positional[63055:63052], addr_15763_7);

wire[31:0] addr_15764_7;

Selector_2 s15764_7(wires_3941_6[0], addr_3941_6, addr_positional[63059:63056], addr_15764_7);

wire[31:0] addr_15765_7;

Selector_2 s15765_7(wires_3941_6[1], addr_3941_6, addr_positional[63063:63060], addr_15765_7);

wire[31:0] addr_15766_7;

Selector_2 s15766_7(wires_3941_6[2], addr_3941_6, addr_positional[63067:63064], addr_15766_7);

wire[31:0] addr_15767_7;

Selector_2 s15767_7(wires_3941_6[3], addr_3941_6, addr_positional[63071:63068], addr_15767_7);

wire[31:0] addr_15768_7;

Selector_2 s15768_7(wires_3942_6[0], addr_3942_6, addr_positional[63075:63072], addr_15768_7);

wire[31:0] addr_15769_7;

Selector_2 s15769_7(wires_3942_6[1], addr_3942_6, addr_positional[63079:63076], addr_15769_7);

wire[31:0] addr_15770_7;

Selector_2 s15770_7(wires_3942_6[2], addr_3942_6, addr_positional[63083:63080], addr_15770_7);

wire[31:0] addr_15771_7;

Selector_2 s15771_7(wires_3942_6[3], addr_3942_6, addr_positional[63087:63084], addr_15771_7);

wire[31:0] addr_15772_7;

Selector_2 s15772_7(wires_3943_6[0], addr_3943_6, addr_positional[63091:63088], addr_15772_7);

wire[31:0] addr_15773_7;

Selector_2 s15773_7(wires_3943_6[1], addr_3943_6, addr_positional[63095:63092], addr_15773_7);

wire[31:0] addr_15774_7;

Selector_2 s15774_7(wires_3943_6[2], addr_3943_6, addr_positional[63099:63096], addr_15774_7);

wire[31:0] addr_15775_7;

Selector_2 s15775_7(wires_3943_6[3], addr_3943_6, addr_positional[63103:63100], addr_15775_7);

wire[31:0] addr_15776_7;

Selector_2 s15776_7(wires_3944_6[0], addr_3944_6, addr_positional[63107:63104], addr_15776_7);

wire[31:0] addr_15777_7;

Selector_2 s15777_7(wires_3944_6[1], addr_3944_6, addr_positional[63111:63108], addr_15777_7);

wire[31:0] addr_15778_7;

Selector_2 s15778_7(wires_3944_6[2], addr_3944_6, addr_positional[63115:63112], addr_15778_7);

wire[31:0] addr_15779_7;

Selector_2 s15779_7(wires_3944_6[3], addr_3944_6, addr_positional[63119:63116], addr_15779_7);

wire[31:0] addr_15780_7;

Selector_2 s15780_7(wires_3945_6[0], addr_3945_6, addr_positional[63123:63120], addr_15780_7);

wire[31:0] addr_15781_7;

Selector_2 s15781_7(wires_3945_6[1], addr_3945_6, addr_positional[63127:63124], addr_15781_7);

wire[31:0] addr_15782_7;

Selector_2 s15782_7(wires_3945_6[2], addr_3945_6, addr_positional[63131:63128], addr_15782_7);

wire[31:0] addr_15783_7;

Selector_2 s15783_7(wires_3945_6[3], addr_3945_6, addr_positional[63135:63132], addr_15783_7);

wire[31:0] addr_15784_7;

Selector_2 s15784_7(wires_3946_6[0], addr_3946_6, addr_positional[63139:63136], addr_15784_7);

wire[31:0] addr_15785_7;

Selector_2 s15785_7(wires_3946_6[1], addr_3946_6, addr_positional[63143:63140], addr_15785_7);

wire[31:0] addr_15786_7;

Selector_2 s15786_7(wires_3946_6[2], addr_3946_6, addr_positional[63147:63144], addr_15786_7);

wire[31:0] addr_15787_7;

Selector_2 s15787_7(wires_3946_6[3], addr_3946_6, addr_positional[63151:63148], addr_15787_7);

wire[31:0] addr_15788_7;

Selector_2 s15788_7(wires_3947_6[0], addr_3947_6, addr_positional[63155:63152], addr_15788_7);

wire[31:0] addr_15789_7;

Selector_2 s15789_7(wires_3947_6[1], addr_3947_6, addr_positional[63159:63156], addr_15789_7);

wire[31:0] addr_15790_7;

Selector_2 s15790_7(wires_3947_6[2], addr_3947_6, addr_positional[63163:63160], addr_15790_7);

wire[31:0] addr_15791_7;

Selector_2 s15791_7(wires_3947_6[3], addr_3947_6, addr_positional[63167:63164], addr_15791_7);

wire[31:0] addr_15792_7;

Selector_2 s15792_7(wires_3948_6[0], addr_3948_6, addr_positional[63171:63168], addr_15792_7);

wire[31:0] addr_15793_7;

Selector_2 s15793_7(wires_3948_6[1], addr_3948_6, addr_positional[63175:63172], addr_15793_7);

wire[31:0] addr_15794_7;

Selector_2 s15794_7(wires_3948_6[2], addr_3948_6, addr_positional[63179:63176], addr_15794_7);

wire[31:0] addr_15795_7;

Selector_2 s15795_7(wires_3948_6[3], addr_3948_6, addr_positional[63183:63180], addr_15795_7);

wire[31:0] addr_15796_7;

Selector_2 s15796_7(wires_3949_6[0], addr_3949_6, addr_positional[63187:63184], addr_15796_7);

wire[31:0] addr_15797_7;

Selector_2 s15797_7(wires_3949_6[1], addr_3949_6, addr_positional[63191:63188], addr_15797_7);

wire[31:0] addr_15798_7;

Selector_2 s15798_7(wires_3949_6[2], addr_3949_6, addr_positional[63195:63192], addr_15798_7);

wire[31:0] addr_15799_7;

Selector_2 s15799_7(wires_3949_6[3], addr_3949_6, addr_positional[63199:63196], addr_15799_7);

wire[31:0] addr_15800_7;

Selector_2 s15800_7(wires_3950_6[0], addr_3950_6, addr_positional[63203:63200], addr_15800_7);

wire[31:0] addr_15801_7;

Selector_2 s15801_7(wires_3950_6[1], addr_3950_6, addr_positional[63207:63204], addr_15801_7);

wire[31:0] addr_15802_7;

Selector_2 s15802_7(wires_3950_6[2], addr_3950_6, addr_positional[63211:63208], addr_15802_7);

wire[31:0] addr_15803_7;

Selector_2 s15803_7(wires_3950_6[3], addr_3950_6, addr_positional[63215:63212], addr_15803_7);

wire[31:0] addr_15804_7;

Selector_2 s15804_7(wires_3951_6[0], addr_3951_6, addr_positional[63219:63216], addr_15804_7);

wire[31:0] addr_15805_7;

Selector_2 s15805_7(wires_3951_6[1], addr_3951_6, addr_positional[63223:63220], addr_15805_7);

wire[31:0] addr_15806_7;

Selector_2 s15806_7(wires_3951_6[2], addr_3951_6, addr_positional[63227:63224], addr_15806_7);

wire[31:0] addr_15807_7;

Selector_2 s15807_7(wires_3951_6[3], addr_3951_6, addr_positional[63231:63228], addr_15807_7);

wire[31:0] addr_15808_7;

Selector_2 s15808_7(wires_3952_6[0], addr_3952_6, addr_positional[63235:63232], addr_15808_7);

wire[31:0] addr_15809_7;

Selector_2 s15809_7(wires_3952_6[1], addr_3952_6, addr_positional[63239:63236], addr_15809_7);

wire[31:0] addr_15810_7;

Selector_2 s15810_7(wires_3952_6[2], addr_3952_6, addr_positional[63243:63240], addr_15810_7);

wire[31:0] addr_15811_7;

Selector_2 s15811_7(wires_3952_6[3], addr_3952_6, addr_positional[63247:63244], addr_15811_7);

wire[31:0] addr_15812_7;

Selector_2 s15812_7(wires_3953_6[0], addr_3953_6, addr_positional[63251:63248], addr_15812_7);

wire[31:0] addr_15813_7;

Selector_2 s15813_7(wires_3953_6[1], addr_3953_6, addr_positional[63255:63252], addr_15813_7);

wire[31:0] addr_15814_7;

Selector_2 s15814_7(wires_3953_6[2], addr_3953_6, addr_positional[63259:63256], addr_15814_7);

wire[31:0] addr_15815_7;

Selector_2 s15815_7(wires_3953_6[3], addr_3953_6, addr_positional[63263:63260], addr_15815_7);

wire[31:0] addr_15816_7;

Selector_2 s15816_7(wires_3954_6[0], addr_3954_6, addr_positional[63267:63264], addr_15816_7);

wire[31:0] addr_15817_7;

Selector_2 s15817_7(wires_3954_6[1], addr_3954_6, addr_positional[63271:63268], addr_15817_7);

wire[31:0] addr_15818_7;

Selector_2 s15818_7(wires_3954_6[2], addr_3954_6, addr_positional[63275:63272], addr_15818_7);

wire[31:0] addr_15819_7;

Selector_2 s15819_7(wires_3954_6[3], addr_3954_6, addr_positional[63279:63276], addr_15819_7);

wire[31:0] addr_15820_7;

Selector_2 s15820_7(wires_3955_6[0], addr_3955_6, addr_positional[63283:63280], addr_15820_7);

wire[31:0] addr_15821_7;

Selector_2 s15821_7(wires_3955_6[1], addr_3955_6, addr_positional[63287:63284], addr_15821_7);

wire[31:0] addr_15822_7;

Selector_2 s15822_7(wires_3955_6[2], addr_3955_6, addr_positional[63291:63288], addr_15822_7);

wire[31:0] addr_15823_7;

Selector_2 s15823_7(wires_3955_6[3], addr_3955_6, addr_positional[63295:63292], addr_15823_7);

wire[31:0] addr_15824_7;

Selector_2 s15824_7(wires_3956_6[0], addr_3956_6, addr_positional[63299:63296], addr_15824_7);

wire[31:0] addr_15825_7;

Selector_2 s15825_7(wires_3956_6[1], addr_3956_6, addr_positional[63303:63300], addr_15825_7);

wire[31:0] addr_15826_7;

Selector_2 s15826_7(wires_3956_6[2], addr_3956_6, addr_positional[63307:63304], addr_15826_7);

wire[31:0] addr_15827_7;

Selector_2 s15827_7(wires_3956_6[3], addr_3956_6, addr_positional[63311:63308], addr_15827_7);

wire[31:0] addr_15828_7;

Selector_2 s15828_7(wires_3957_6[0], addr_3957_6, addr_positional[63315:63312], addr_15828_7);

wire[31:0] addr_15829_7;

Selector_2 s15829_7(wires_3957_6[1], addr_3957_6, addr_positional[63319:63316], addr_15829_7);

wire[31:0] addr_15830_7;

Selector_2 s15830_7(wires_3957_6[2], addr_3957_6, addr_positional[63323:63320], addr_15830_7);

wire[31:0] addr_15831_7;

Selector_2 s15831_7(wires_3957_6[3], addr_3957_6, addr_positional[63327:63324], addr_15831_7);

wire[31:0] addr_15832_7;

Selector_2 s15832_7(wires_3958_6[0], addr_3958_6, addr_positional[63331:63328], addr_15832_7);

wire[31:0] addr_15833_7;

Selector_2 s15833_7(wires_3958_6[1], addr_3958_6, addr_positional[63335:63332], addr_15833_7);

wire[31:0] addr_15834_7;

Selector_2 s15834_7(wires_3958_6[2], addr_3958_6, addr_positional[63339:63336], addr_15834_7);

wire[31:0] addr_15835_7;

Selector_2 s15835_7(wires_3958_6[3], addr_3958_6, addr_positional[63343:63340], addr_15835_7);

wire[31:0] addr_15836_7;

Selector_2 s15836_7(wires_3959_6[0], addr_3959_6, addr_positional[63347:63344], addr_15836_7);

wire[31:0] addr_15837_7;

Selector_2 s15837_7(wires_3959_6[1], addr_3959_6, addr_positional[63351:63348], addr_15837_7);

wire[31:0] addr_15838_7;

Selector_2 s15838_7(wires_3959_6[2], addr_3959_6, addr_positional[63355:63352], addr_15838_7);

wire[31:0] addr_15839_7;

Selector_2 s15839_7(wires_3959_6[3], addr_3959_6, addr_positional[63359:63356], addr_15839_7);

wire[31:0] addr_15840_7;

Selector_2 s15840_7(wires_3960_6[0], addr_3960_6, addr_positional[63363:63360], addr_15840_7);

wire[31:0] addr_15841_7;

Selector_2 s15841_7(wires_3960_6[1], addr_3960_6, addr_positional[63367:63364], addr_15841_7);

wire[31:0] addr_15842_7;

Selector_2 s15842_7(wires_3960_6[2], addr_3960_6, addr_positional[63371:63368], addr_15842_7);

wire[31:0] addr_15843_7;

Selector_2 s15843_7(wires_3960_6[3], addr_3960_6, addr_positional[63375:63372], addr_15843_7);

wire[31:0] addr_15844_7;

Selector_2 s15844_7(wires_3961_6[0], addr_3961_6, addr_positional[63379:63376], addr_15844_7);

wire[31:0] addr_15845_7;

Selector_2 s15845_7(wires_3961_6[1], addr_3961_6, addr_positional[63383:63380], addr_15845_7);

wire[31:0] addr_15846_7;

Selector_2 s15846_7(wires_3961_6[2], addr_3961_6, addr_positional[63387:63384], addr_15846_7);

wire[31:0] addr_15847_7;

Selector_2 s15847_7(wires_3961_6[3], addr_3961_6, addr_positional[63391:63388], addr_15847_7);

wire[31:0] addr_15848_7;

Selector_2 s15848_7(wires_3962_6[0], addr_3962_6, addr_positional[63395:63392], addr_15848_7);

wire[31:0] addr_15849_7;

Selector_2 s15849_7(wires_3962_6[1], addr_3962_6, addr_positional[63399:63396], addr_15849_7);

wire[31:0] addr_15850_7;

Selector_2 s15850_7(wires_3962_6[2], addr_3962_6, addr_positional[63403:63400], addr_15850_7);

wire[31:0] addr_15851_7;

Selector_2 s15851_7(wires_3962_6[3], addr_3962_6, addr_positional[63407:63404], addr_15851_7);

wire[31:0] addr_15852_7;

Selector_2 s15852_7(wires_3963_6[0], addr_3963_6, addr_positional[63411:63408], addr_15852_7);

wire[31:0] addr_15853_7;

Selector_2 s15853_7(wires_3963_6[1], addr_3963_6, addr_positional[63415:63412], addr_15853_7);

wire[31:0] addr_15854_7;

Selector_2 s15854_7(wires_3963_6[2], addr_3963_6, addr_positional[63419:63416], addr_15854_7);

wire[31:0] addr_15855_7;

Selector_2 s15855_7(wires_3963_6[3], addr_3963_6, addr_positional[63423:63420], addr_15855_7);

wire[31:0] addr_15856_7;

Selector_2 s15856_7(wires_3964_6[0], addr_3964_6, addr_positional[63427:63424], addr_15856_7);

wire[31:0] addr_15857_7;

Selector_2 s15857_7(wires_3964_6[1], addr_3964_6, addr_positional[63431:63428], addr_15857_7);

wire[31:0] addr_15858_7;

Selector_2 s15858_7(wires_3964_6[2], addr_3964_6, addr_positional[63435:63432], addr_15858_7);

wire[31:0] addr_15859_7;

Selector_2 s15859_7(wires_3964_6[3], addr_3964_6, addr_positional[63439:63436], addr_15859_7);

wire[31:0] addr_15860_7;

Selector_2 s15860_7(wires_3965_6[0], addr_3965_6, addr_positional[63443:63440], addr_15860_7);

wire[31:0] addr_15861_7;

Selector_2 s15861_7(wires_3965_6[1], addr_3965_6, addr_positional[63447:63444], addr_15861_7);

wire[31:0] addr_15862_7;

Selector_2 s15862_7(wires_3965_6[2], addr_3965_6, addr_positional[63451:63448], addr_15862_7);

wire[31:0] addr_15863_7;

Selector_2 s15863_7(wires_3965_6[3], addr_3965_6, addr_positional[63455:63452], addr_15863_7);

wire[31:0] addr_15864_7;

Selector_2 s15864_7(wires_3966_6[0], addr_3966_6, addr_positional[63459:63456], addr_15864_7);

wire[31:0] addr_15865_7;

Selector_2 s15865_7(wires_3966_6[1], addr_3966_6, addr_positional[63463:63460], addr_15865_7);

wire[31:0] addr_15866_7;

Selector_2 s15866_7(wires_3966_6[2], addr_3966_6, addr_positional[63467:63464], addr_15866_7);

wire[31:0] addr_15867_7;

Selector_2 s15867_7(wires_3966_6[3], addr_3966_6, addr_positional[63471:63468], addr_15867_7);

wire[31:0] addr_15868_7;

Selector_2 s15868_7(wires_3967_6[0], addr_3967_6, addr_positional[63475:63472], addr_15868_7);

wire[31:0] addr_15869_7;

Selector_2 s15869_7(wires_3967_6[1], addr_3967_6, addr_positional[63479:63476], addr_15869_7);

wire[31:0] addr_15870_7;

Selector_2 s15870_7(wires_3967_6[2], addr_3967_6, addr_positional[63483:63480], addr_15870_7);

wire[31:0] addr_15871_7;

Selector_2 s15871_7(wires_3967_6[3], addr_3967_6, addr_positional[63487:63484], addr_15871_7);

wire[31:0] addr_15872_7;

Selector_2 s15872_7(wires_3968_6[0], addr_3968_6, addr_positional[63491:63488], addr_15872_7);

wire[31:0] addr_15873_7;

Selector_2 s15873_7(wires_3968_6[1], addr_3968_6, addr_positional[63495:63492], addr_15873_7);

wire[31:0] addr_15874_7;

Selector_2 s15874_7(wires_3968_6[2], addr_3968_6, addr_positional[63499:63496], addr_15874_7);

wire[31:0] addr_15875_7;

Selector_2 s15875_7(wires_3968_6[3], addr_3968_6, addr_positional[63503:63500], addr_15875_7);

wire[31:0] addr_15876_7;

Selector_2 s15876_7(wires_3969_6[0], addr_3969_6, addr_positional[63507:63504], addr_15876_7);

wire[31:0] addr_15877_7;

Selector_2 s15877_7(wires_3969_6[1], addr_3969_6, addr_positional[63511:63508], addr_15877_7);

wire[31:0] addr_15878_7;

Selector_2 s15878_7(wires_3969_6[2], addr_3969_6, addr_positional[63515:63512], addr_15878_7);

wire[31:0] addr_15879_7;

Selector_2 s15879_7(wires_3969_6[3], addr_3969_6, addr_positional[63519:63516], addr_15879_7);

wire[31:0] addr_15880_7;

Selector_2 s15880_7(wires_3970_6[0], addr_3970_6, addr_positional[63523:63520], addr_15880_7);

wire[31:0] addr_15881_7;

Selector_2 s15881_7(wires_3970_6[1], addr_3970_6, addr_positional[63527:63524], addr_15881_7);

wire[31:0] addr_15882_7;

Selector_2 s15882_7(wires_3970_6[2], addr_3970_6, addr_positional[63531:63528], addr_15882_7);

wire[31:0] addr_15883_7;

Selector_2 s15883_7(wires_3970_6[3], addr_3970_6, addr_positional[63535:63532], addr_15883_7);

wire[31:0] addr_15884_7;

Selector_2 s15884_7(wires_3971_6[0], addr_3971_6, addr_positional[63539:63536], addr_15884_7);

wire[31:0] addr_15885_7;

Selector_2 s15885_7(wires_3971_6[1], addr_3971_6, addr_positional[63543:63540], addr_15885_7);

wire[31:0] addr_15886_7;

Selector_2 s15886_7(wires_3971_6[2], addr_3971_6, addr_positional[63547:63544], addr_15886_7);

wire[31:0] addr_15887_7;

Selector_2 s15887_7(wires_3971_6[3], addr_3971_6, addr_positional[63551:63548], addr_15887_7);

wire[31:0] addr_15888_7;

Selector_2 s15888_7(wires_3972_6[0], addr_3972_6, addr_positional[63555:63552], addr_15888_7);

wire[31:0] addr_15889_7;

Selector_2 s15889_7(wires_3972_6[1], addr_3972_6, addr_positional[63559:63556], addr_15889_7);

wire[31:0] addr_15890_7;

Selector_2 s15890_7(wires_3972_6[2], addr_3972_6, addr_positional[63563:63560], addr_15890_7);

wire[31:0] addr_15891_7;

Selector_2 s15891_7(wires_3972_6[3], addr_3972_6, addr_positional[63567:63564], addr_15891_7);

wire[31:0] addr_15892_7;

Selector_2 s15892_7(wires_3973_6[0], addr_3973_6, addr_positional[63571:63568], addr_15892_7);

wire[31:0] addr_15893_7;

Selector_2 s15893_7(wires_3973_6[1], addr_3973_6, addr_positional[63575:63572], addr_15893_7);

wire[31:0] addr_15894_7;

Selector_2 s15894_7(wires_3973_6[2], addr_3973_6, addr_positional[63579:63576], addr_15894_7);

wire[31:0] addr_15895_7;

Selector_2 s15895_7(wires_3973_6[3], addr_3973_6, addr_positional[63583:63580], addr_15895_7);

wire[31:0] addr_15896_7;

Selector_2 s15896_7(wires_3974_6[0], addr_3974_6, addr_positional[63587:63584], addr_15896_7);

wire[31:0] addr_15897_7;

Selector_2 s15897_7(wires_3974_6[1], addr_3974_6, addr_positional[63591:63588], addr_15897_7);

wire[31:0] addr_15898_7;

Selector_2 s15898_7(wires_3974_6[2], addr_3974_6, addr_positional[63595:63592], addr_15898_7);

wire[31:0] addr_15899_7;

Selector_2 s15899_7(wires_3974_6[3], addr_3974_6, addr_positional[63599:63596], addr_15899_7);

wire[31:0] addr_15900_7;

Selector_2 s15900_7(wires_3975_6[0], addr_3975_6, addr_positional[63603:63600], addr_15900_7);

wire[31:0] addr_15901_7;

Selector_2 s15901_7(wires_3975_6[1], addr_3975_6, addr_positional[63607:63604], addr_15901_7);

wire[31:0] addr_15902_7;

Selector_2 s15902_7(wires_3975_6[2], addr_3975_6, addr_positional[63611:63608], addr_15902_7);

wire[31:0] addr_15903_7;

Selector_2 s15903_7(wires_3975_6[3], addr_3975_6, addr_positional[63615:63612], addr_15903_7);

wire[31:0] addr_15904_7;

Selector_2 s15904_7(wires_3976_6[0], addr_3976_6, addr_positional[63619:63616], addr_15904_7);

wire[31:0] addr_15905_7;

Selector_2 s15905_7(wires_3976_6[1], addr_3976_6, addr_positional[63623:63620], addr_15905_7);

wire[31:0] addr_15906_7;

Selector_2 s15906_7(wires_3976_6[2], addr_3976_6, addr_positional[63627:63624], addr_15906_7);

wire[31:0] addr_15907_7;

Selector_2 s15907_7(wires_3976_6[3], addr_3976_6, addr_positional[63631:63628], addr_15907_7);

wire[31:0] addr_15908_7;

Selector_2 s15908_7(wires_3977_6[0], addr_3977_6, addr_positional[63635:63632], addr_15908_7);

wire[31:0] addr_15909_7;

Selector_2 s15909_7(wires_3977_6[1], addr_3977_6, addr_positional[63639:63636], addr_15909_7);

wire[31:0] addr_15910_7;

Selector_2 s15910_7(wires_3977_6[2], addr_3977_6, addr_positional[63643:63640], addr_15910_7);

wire[31:0] addr_15911_7;

Selector_2 s15911_7(wires_3977_6[3], addr_3977_6, addr_positional[63647:63644], addr_15911_7);

wire[31:0] addr_15912_7;

Selector_2 s15912_7(wires_3978_6[0], addr_3978_6, addr_positional[63651:63648], addr_15912_7);

wire[31:0] addr_15913_7;

Selector_2 s15913_7(wires_3978_6[1], addr_3978_6, addr_positional[63655:63652], addr_15913_7);

wire[31:0] addr_15914_7;

Selector_2 s15914_7(wires_3978_6[2], addr_3978_6, addr_positional[63659:63656], addr_15914_7);

wire[31:0] addr_15915_7;

Selector_2 s15915_7(wires_3978_6[3], addr_3978_6, addr_positional[63663:63660], addr_15915_7);

wire[31:0] addr_15916_7;

Selector_2 s15916_7(wires_3979_6[0], addr_3979_6, addr_positional[63667:63664], addr_15916_7);

wire[31:0] addr_15917_7;

Selector_2 s15917_7(wires_3979_6[1], addr_3979_6, addr_positional[63671:63668], addr_15917_7);

wire[31:0] addr_15918_7;

Selector_2 s15918_7(wires_3979_6[2], addr_3979_6, addr_positional[63675:63672], addr_15918_7);

wire[31:0] addr_15919_7;

Selector_2 s15919_7(wires_3979_6[3], addr_3979_6, addr_positional[63679:63676], addr_15919_7);

wire[31:0] addr_15920_7;

Selector_2 s15920_7(wires_3980_6[0], addr_3980_6, addr_positional[63683:63680], addr_15920_7);

wire[31:0] addr_15921_7;

Selector_2 s15921_7(wires_3980_6[1], addr_3980_6, addr_positional[63687:63684], addr_15921_7);

wire[31:0] addr_15922_7;

Selector_2 s15922_7(wires_3980_6[2], addr_3980_6, addr_positional[63691:63688], addr_15922_7);

wire[31:0] addr_15923_7;

Selector_2 s15923_7(wires_3980_6[3], addr_3980_6, addr_positional[63695:63692], addr_15923_7);

wire[31:0] addr_15924_7;

Selector_2 s15924_7(wires_3981_6[0], addr_3981_6, addr_positional[63699:63696], addr_15924_7);

wire[31:0] addr_15925_7;

Selector_2 s15925_7(wires_3981_6[1], addr_3981_6, addr_positional[63703:63700], addr_15925_7);

wire[31:0] addr_15926_7;

Selector_2 s15926_7(wires_3981_6[2], addr_3981_6, addr_positional[63707:63704], addr_15926_7);

wire[31:0] addr_15927_7;

Selector_2 s15927_7(wires_3981_6[3], addr_3981_6, addr_positional[63711:63708], addr_15927_7);

wire[31:0] addr_15928_7;

Selector_2 s15928_7(wires_3982_6[0], addr_3982_6, addr_positional[63715:63712], addr_15928_7);

wire[31:0] addr_15929_7;

Selector_2 s15929_7(wires_3982_6[1], addr_3982_6, addr_positional[63719:63716], addr_15929_7);

wire[31:0] addr_15930_7;

Selector_2 s15930_7(wires_3982_6[2], addr_3982_6, addr_positional[63723:63720], addr_15930_7);

wire[31:0] addr_15931_7;

Selector_2 s15931_7(wires_3982_6[3], addr_3982_6, addr_positional[63727:63724], addr_15931_7);

wire[31:0] addr_15932_7;

Selector_2 s15932_7(wires_3983_6[0], addr_3983_6, addr_positional[63731:63728], addr_15932_7);

wire[31:0] addr_15933_7;

Selector_2 s15933_7(wires_3983_6[1], addr_3983_6, addr_positional[63735:63732], addr_15933_7);

wire[31:0] addr_15934_7;

Selector_2 s15934_7(wires_3983_6[2], addr_3983_6, addr_positional[63739:63736], addr_15934_7);

wire[31:0] addr_15935_7;

Selector_2 s15935_7(wires_3983_6[3], addr_3983_6, addr_positional[63743:63740], addr_15935_7);

wire[31:0] addr_15936_7;

Selector_2 s15936_7(wires_3984_6[0], addr_3984_6, addr_positional[63747:63744], addr_15936_7);

wire[31:0] addr_15937_7;

Selector_2 s15937_7(wires_3984_6[1], addr_3984_6, addr_positional[63751:63748], addr_15937_7);

wire[31:0] addr_15938_7;

Selector_2 s15938_7(wires_3984_6[2], addr_3984_6, addr_positional[63755:63752], addr_15938_7);

wire[31:0] addr_15939_7;

Selector_2 s15939_7(wires_3984_6[3], addr_3984_6, addr_positional[63759:63756], addr_15939_7);

wire[31:0] addr_15940_7;

Selector_2 s15940_7(wires_3985_6[0], addr_3985_6, addr_positional[63763:63760], addr_15940_7);

wire[31:0] addr_15941_7;

Selector_2 s15941_7(wires_3985_6[1], addr_3985_6, addr_positional[63767:63764], addr_15941_7);

wire[31:0] addr_15942_7;

Selector_2 s15942_7(wires_3985_6[2], addr_3985_6, addr_positional[63771:63768], addr_15942_7);

wire[31:0] addr_15943_7;

Selector_2 s15943_7(wires_3985_6[3], addr_3985_6, addr_positional[63775:63772], addr_15943_7);

wire[31:0] addr_15944_7;

Selector_2 s15944_7(wires_3986_6[0], addr_3986_6, addr_positional[63779:63776], addr_15944_7);

wire[31:0] addr_15945_7;

Selector_2 s15945_7(wires_3986_6[1], addr_3986_6, addr_positional[63783:63780], addr_15945_7);

wire[31:0] addr_15946_7;

Selector_2 s15946_7(wires_3986_6[2], addr_3986_6, addr_positional[63787:63784], addr_15946_7);

wire[31:0] addr_15947_7;

Selector_2 s15947_7(wires_3986_6[3], addr_3986_6, addr_positional[63791:63788], addr_15947_7);

wire[31:0] addr_15948_7;

Selector_2 s15948_7(wires_3987_6[0], addr_3987_6, addr_positional[63795:63792], addr_15948_7);

wire[31:0] addr_15949_7;

Selector_2 s15949_7(wires_3987_6[1], addr_3987_6, addr_positional[63799:63796], addr_15949_7);

wire[31:0] addr_15950_7;

Selector_2 s15950_7(wires_3987_6[2], addr_3987_6, addr_positional[63803:63800], addr_15950_7);

wire[31:0] addr_15951_7;

Selector_2 s15951_7(wires_3987_6[3], addr_3987_6, addr_positional[63807:63804], addr_15951_7);

wire[31:0] addr_15952_7;

Selector_2 s15952_7(wires_3988_6[0], addr_3988_6, addr_positional[63811:63808], addr_15952_7);

wire[31:0] addr_15953_7;

Selector_2 s15953_7(wires_3988_6[1], addr_3988_6, addr_positional[63815:63812], addr_15953_7);

wire[31:0] addr_15954_7;

Selector_2 s15954_7(wires_3988_6[2], addr_3988_6, addr_positional[63819:63816], addr_15954_7);

wire[31:0] addr_15955_7;

Selector_2 s15955_7(wires_3988_6[3], addr_3988_6, addr_positional[63823:63820], addr_15955_7);

wire[31:0] addr_15956_7;

Selector_2 s15956_7(wires_3989_6[0], addr_3989_6, addr_positional[63827:63824], addr_15956_7);

wire[31:0] addr_15957_7;

Selector_2 s15957_7(wires_3989_6[1], addr_3989_6, addr_positional[63831:63828], addr_15957_7);

wire[31:0] addr_15958_7;

Selector_2 s15958_7(wires_3989_6[2], addr_3989_6, addr_positional[63835:63832], addr_15958_7);

wire[31:0] addr_15959_7;

Selector_2 s15959_7(wires_3989_6[3], addr_3989_6, addr_positional[63839:63836], addr_15959_7);

wire[31:0] addr_15960_7;

Selector_2 s15960_7(wires_3990_6[0], addr_3990_6, addr_positional[63843:63840], addr_15960_7);

wire[31:0] addr_15961_7;

Selector_2 s15961_7(wires_3990_6[1], addr_3990_6, addr_positional[63847:63844], addr_15961_7);

wire[31:0] addr_15962_7;

Selector_2 s15962_7(wires_3990_6[2], addr_3990_6, addr_positional[63851:63848], addr_15962_7);

wire[31:0] addr_15963_7;

Selector_2 s15963_7(wires_3990_6[3], addr_3990_6, addr_positional[63855:63852], addr_15963_7);

wire[31:0] addr_15964_7;

Selector_2 s15964_7(wires_3991_6[0], addr_3991_6, addr_positional[63859:63856], addr_15964_7);

wire[31:0] addr_15965_7;

Selector_2 s15965_7(wires_3991_6[1], addr_3991_6, addr_positional[63863:63860], addr_15965_7);

wire[31:0] addr_15966_7;

Selector_2 s15966_7(wires_3991_6[2], addr_3991_6, addr_positional[63867:63864], addr_15966_7);

wire[31:0] addr_15967_7;

Selector_2 s15967_7(wires_3991_6[3], addr_3991_6, addr_positional[63871:63868], addr_15967_7);

wire[31:0] addr_15968_7;

Selector_2 s15968_7(wires_3992_6[0], addr_3992_6, addr_positional[63875:63872], addr_15968_7);

wire[31:0] addr_15969_7;

Selector_2 s15969_7(wires_3992_6[1], addr_3992_6, addr_positional[63879:63876], addr_15969_7);

wire[31:0] addr_15970_7;

Selector_2 s15970_7(wires_3992_6[2], addr_3992_6, addr_positional[63883:63880], addr_15970_7);

wire[31:0] addr_15971_7;

Selector_2 s15971_7(wires_3992_6[3], addr_3992_6, addr_positional[63887:63884], addr_15971_7);

wire[31:0] addr_15972_7;

Selector_2 s15972_7(wires_3993_6[0], addr_3993_6, addr_positional[63891:63888], addr_15972_7);

wire[31:0] addr_15973_7;

Selector_2 s15973_7(wires_3993_6[1], addr_3993_6, addr_positional[63895:63892], addr_15973_7);

wire[31:0] addr_15974_7;

Selector_2 s15974_7(wires_3993_6[2], addr_3993_6, addr_positional[63899:63896], addr_15974_7);

wire[31:0] addr_15975_7;

Selector_2 s15975_7(wires_3993_6[3], addr_3993_6, addr_positional[63903:63900], addr_15975_7);

wire[31:0] addr_15976_7;

Selector_2 s15976_7(wires_3994_6[0], addr_3994_6, addr_positional[63907:63904], addr_15976_7);

wire[31:0] addr_15977_7;

Selector_2 s15977_7(wires_3994_6[1], addr_3994_6, addr_positional[63911:63908], addr_15977_7);

wire[31:0] addr_15978_7;

Selector_2 s15978_7(wires_3994_6[2], addr_3994_6, addr_positional[63915:63912], addr_15978_7);

wire[31:0] addr_15979_7;

Selector_2 s15979_7(wires_3994_6[3], addr_3994_6, addr_positional[63919:63916], addr_15979_7);

wire[31:0] addr_15980_7;

Selector_2 s15980_7(wires_3995_6[0], addr_3995_6, addr_positional[63923:63920], addr_15980_7);

wire[31:0] addr_15981_7;

Selector_2 s15981_7(wires_3995_6[1], addr_3995_6, addr_positional[63927:63924], addr_15981_7);

wire[31:0] addr_15982_7;

Selector_2 s15982_7(wires_3995_6[2], addr_3995_6, addr_positional[63931:63928], addr_15982_7);

wire[31:0] addr_15983_7;

Selector_2 s15983_7(wires_3995_6[3], addr_3995_6, addr_positional[63935:63932], addr_15983_7);

wire[31:0] addr_15984_7;

Selector_2 s15984_7(wires_3996_6[0], addr_3996_6, addr_positional[63939:63936], addr_15984_7);

wire[31:0] addr_15985_7;

Selector_2 s15985_7(wires_3996_6[1], addr_3996_6, addr_positional[63943:63940], addr_15985_7);

wire[31:0] addr_15986_7;

Selector_2 s15986_7(wires_3996_6[2], addr_3996_6, addr_positional[63947:63944], addr_15986_7);

wire[31:0] addr_15987_7;

Selector_2 s15987_7(wires_3996_6[3], addr_3996_6, addr_positional[63951:63948], addr_15987_7);

wire[31:0] addr_15988_7;

Selector_2 s15988_7(wires_3997_6[0], addr_3997_6, addr_positional[63955:63952], addr_15988_7);

wire[31:0] addr_15989_7;

Selector_2 s15989_7(wires_3997_6[1], addr_3997_6, addr_positional[63959:63956], addr_15989_7);

wire[31:0] addr_15990_7;

Selector_2 s15990_7(wires_3997_6[2], addr_3997_6, addr_positional[63963:63960], addr_15990_7);

wire[31:0] addr_15991_7;

Selector_2 s15991_7(wires_3997_6[3], addr_3997_6, addr_positional[63967:63964], addr_15991_7);

wire[31:0] addr_15992_7;

Selector_2 s15992_7(wires_3998_6[0], addr_3998_6, addr_positional[63971:63968], addr_15992_7);

wire[31:0] addr_15993_7;

Selector_2 s15993_7(wires_3998_6[1], addr_3998_6, addr_positional[63975:63972], addr_15993_7);

wire[31:0] addr_15994_7;

Selector_2 s15994_7(wires_3998_6[2], addr_3998_6, addr_positional[63979:63976], addr_15994_7);

wire[31:0] addr_15995_7;

Selector_2 s15995_7(wires_3998_6[3], addr_3998_6, addr_positional[63983:63980], addr_15995_7);

wire[31:0] addr_15996_7;

Selector_2 s15996_7(wires_3999_6[0], addr_3999_6, addr_positional[63987:63984], addr_15996_7);

wire[31:0] addr_15997_7;

Selector_2 s15997_7(wires_3999_6[1], addr_3999_6, addr_positional[63991:63988], addr_15997_7);

wire[31:0] addr_15998_7;

Selector_2 s15998_7(wires_3999_6[2], addr_3999_6, addr_positional[63995:63992], addr_15998_7);

wire[31:0] addr_15999_7;

Selector_2 s15999_7(wires_3999_6[3], addr_3999_6, addr_positional[63999:63996], addr_15999_7);

wire[31:0] addr_16000_7;

Selector_2 s16000_7(wires_4000_6[0], addr_4000_6, addr_positional[64003:64000], addr_16000_7);

wire[31:0] addr_16001_7;

Selector_2 s16001_7(wires_4000_6[1], addr_4000_6, addr_positional[64007:64004], addr_16001_7);

wire[31:0] addr_16002_7;

Selector_2 s16002_7(wires_4000_6[2], addr_4000_6, addr_positional[64011:64008], addr_16002_7);

wire[31:0] addr_16003_7;

Selector_2 s16003_7(wires_4000_6[3], addr_4000_6, addr_positional[64015:64012], addr_16003_7);

wire[31:0] addr_16004_7;

Selector_2 s16004_7(wires_4001_6[0], addr_4001_6, addr_positional[64019:64016], addr_16004_7);

wire[31:0] addr_16005_7;

Selector_2 s16005_7(wires_4001_6[1], addr_4001_6, addr_positional[64023:64020], addr_16005_7);

wire[31:0] addr_16006_7;

Selector_2 s16006_7(wires_4001_6[2], addr_4001_6, addr_positional[64027:64024], addr_16006_7);

wire[31:0] addr_16007_7;

Selector_2 s16007_7(wires_4001_6[3], addr_4001_6, addr_positional[64031:64028], addr_16007_7);

wire[31:0] addr_16008_7;

Selector_2 s16008_7(wires_4002_6[0], addr_4002_6, addr_positional[64035:64032], addr_16008_7);

wire[31:0] addr_16009_7;

Selector_2 s16009_7(wires_4002_6[1], addr_4002_6, addr_positional[64039:64036], addr_16009_7);

wire[31:0] addr_16010_7;

Selector_2 s16010_7(wires_4002_6[2], addr_4002_6, addr_positional[64043:64040], addr_16010_7);

wire[31:0] addr_16011_7;

Selector_2 s16011_7(wires_4002_6[3], addr_4002_6, addr_positional[64047:64044], addr_16011_7);

wire[31:0] addr_16012_7;

Selector_2 s16012_7(wires_4003_6[0], addr_4003_6, addr_positional[64051:64048], addr_16012_7);

wire[31:0] addr_16013_7;

Selector_2 s16013_7(wires_4003_6[1], addr_4003_6, addr_positional[64055:64052], addr_16013_7);

wire[31:0] addr_16014_7;

Selector_2 s16014_7(wires_4003_6[2], addr_4003_6, addr_positional[64059:64056], addr_16014_7);

wire[31:0] addr_16015_7;

Selector_2 s16015_7(wires_4003_6[3], addr_4003_6, addr_positional[64063:64060], addr_16015_7);

wire[31:0] addr_16016_7;

Selector_2 s16016_7(wires_4004_6[0], addr_4004_6, addr_positional[64067:64064], addr_16016_7);

wire[31:0] addr_16017_7;

Selector_2 s16017_7(wires_4004_6[1], addr_4004_6, addr_positional[64071:64068], addr_16017_7);

wire[31:0] addr_16018_7;

Selector_2 s16018_7(wires_4004_6[2], addr_4004_6, addr_positional[64075:64072], addr_16018_7);

wire[31:0] addr_16019_7;

Selector_2 s16019_7(wires_4004_6[3], addr_4004_6, addr_positional[64079:64076], addr_16019_7);

wire[31:0] addr_16020_7;

Selector_2 s16020_7(wires_4005_6[0], addr_4005_6, addr_positional[64083:64080], addr_16020_7);

wire[31:0] addr_16021_7;

Selector_2 s16021_7(wires_4005_6[1], addr_4005_6, addr_positional[64087:64084], addr_16021_7);

wire[31:0] addr_16022_7;

Selector_2 s16022_7(wires_4005_6[2], addr_4005_6, addr_positional[64091:64088], addr_16022_7);

wire[31:0] addr_16023_7;

Selector_2 s16023_7(wires_4005_6[3], addr_4005_6, addr_positional[64095:64092], addr_16023_7);

wire[31:0] addr_16024_7;

Selector_2 s16024_7(wires_4006_6[0], addr_4006_6, addr_positional[64099:64096], addr_16024_7);

wire[31:0] addr_16025_7;

Selector_2 s16025_7(wires_4006_6[1], addr_4006_6, addr_positional[64103:64100], addr_16025_7);

wire[31:0] addr_16026_7;

Selector_2 s16026_7(wires_4006_6[2], addr_4006_6, addr_positional[64107:64104], addr_16026_7);

wire[31:0] addr_16027_7;

Selector_2 s16027_7(wires_4006_6[3], addr_4006_6, addr_positional[64111:64108], addr_16027_7);

wire[31:0] addr_16028_7;

Selector_2 s16028_7(wires_4007_6[0], addr_4007_6, addr_positional[64115:64112], addr_16028_7);

wire[31:0] addr_16029_7;

Selector_2 s16029_7(wires_4007_6[1], addr_4007_6, addr_positional[64119:64116], addr_16029_7);

wire[31:0] addr_16030_7;

Selector_2 s16030_7(wires_4007_6[2], addr_4007_6, addr_positional[64123:64120], addr_16030_7);

wire[31:0] addr_16031_7;

Selector_2 s16031_7(wires_4007_6[3], addr_4007_6, addr_positional[64127:64124], addr_16031_7);

wire[31:0] addr_16032_7;

Selector_2 s16032_7(wires_4008_6[0], addr_4008_6, addr_positional[64131:64128], addr_16032_7);

wire[31:0] addr_16033_7;

Selector_2 s16033_7(wires_4008_6[1], addr_4008_6, addr_positional[64135:64132], addr_16033_7);

wire[31:0] addr_16034_7;

Selector_2 s16034_7(wires_4008_6[2], addr_4008_6, addr_positional[64139:64136], addr_16034_7);

wire[31:0] addr_16035_7;

Selector_2 s16035_7(wires_4008_6[3], addr_4008_6, addr_positional[64143:64140], addr_16035_7);

wire[31:0] addr_16036_7;

Selector_2 s16036_7(wires_4009_6[0], addr_4009_6, addr_positional[64147:64144], addr_16036_7);

wire[31:0] addr_16037_7;

Selector_2 s16037_7(wires_4009_6[1], addr_4009_6, addr_positional[64151:64148], addr_16037_7);

wire[31:0] addr_16038_7;

Selector_2 s16038_7(wires_4009_6[2], addr_4009_6, addr_positional[64155:64152], addr_16038_7);

wire[31:0] addr_16039_7;

Selector_2 s16039_7(wires_4009_6[3], addr_4009_6, addr_positional[64159:64156], addr_16039_7);

wire[31:0] addr_16040_7;

Selector_2 s16040_7(wires_4010_6[0], addr_4010_6, addr_positional[64163:64160], addr_16040_7);

wire[31:0] addr_16041_7;

Selector_2 s16041_7(wires_4010_6[1], addr_4010_6, addr_positional[64167:64164], addr_16041_7);

wire[31:0] addr_16042_7;

Selector_2 s16042_7(wires_4010_6[2], addr_4010_6, addr_positional[64171:64168], addr_16042_7);

wire[31:0] addr_16043_7;

Selector_2 s16043_7(wires_4010_6[3], addr_4010_6, addr_positional[64175:64172], addr_16043_7);

wire[31:0] addr_16044_7;

Selector_2 s16044_7(wires_4011_6[0], addr_4011_6, addr_positional[64179:64176], addr_16044_7);

wire[31:0] addr_16045_7;

Selector_2 s16045_7(wires_4011_6[1], addr_4011_6, addr_positional[64183:64180], addr_16045_7);

wire[31:0] addr_16046_7;

Selector_2 s16046_7(wires_4011_6[2], addr_4011_6, addr_positional[64187:64184], addr_16046_7);

wire[31:0] addr_16047_7;

Selector_2 s16047_7(wires_4011_6[3], addr_4011_6, addr_positional[64191:64188], addr_16047_7);

wire[31:0] addr_16048_7;

Selector_2 s16048_7(wires_4012_6[0], addr_4012_6, addr_positional[64195:64192], addr_16048_7);

wire[31:0] addr_16049_7;

Selector_2 s16049_7(wires_4012_6[1], addr_4012_6, addr_positional[64199:64196], addr_16049_7);

wire[31:0] addr_16050_7;

Selector_2 s16050_7(wires_4012_6[2], addr_4012_6, addr_positional[64203:64200], addr_16050_7);

wire[31:0] addr_16051_7;

Selector_2 s16051_7(wires_4012_6[3], addr_4012_6, addr_positional[64207:64204], addr_16051_7);

wire[31:0] addr_16052_7;

Selector_2 s16052_7(wires_4013_6[0], addr_4013_6, addr_positional[64211:64208], addr_16052_7);

wire[31:0] addr_16053_7;

Selector_2 s16053_7(wires_4013_6[1], addr_4013_6, addr_positional[64215:64212], addr_16053_7);

wire[31:0] addr_16054_7;

Selector_2 s16054_7(wires_4013_6[2], addr_4013_6, addr_positional[64219:64216], addr_16054_7);

wire[31:0] addr_16055_7;

Selector_2 s16055_7(wires_4013_6[3], addr_4013_6, addr_positional[64223:64220], addr_16055_7);

wire[31:0] addr_16056_7;

Selector_2 s16056_7(wires_4014_6[0], addr_4014_6, addr_positional[64227:64224], addr_16056_7);

wire[31:0] addr_16057_7;

Selector_2 s16057_7(wires_4014_6[1], addr_4014_6, addr_positional[64231:64228], addr_16057_7);

wire[31:0] addr_16058_7;

Selector_2 s16058_7(wires_4014_6[2], addr_4014_6, addr_positional[64235:64232], addr_16058_7);

wire[31:0] addr_16059_7;

Selector_2 s16059_7(wires_4014_6[3], addr_4014_6, addr_positional[64239:64236], addr_16059_7);

wire[31:0] addr_16060_7;

Selector_2 s16060_7(wires_4015_6[0], addr_4015_6, addr_positional[64243:64240], addr_16060_7);

wire[31:0] addr_16061_7;

Selector_2 s16061_7(wires_4015_6[1], addr_4015_6, addr_positional[64247:64244], addr_16061_7);

wire[31:0] addr_16062_7;

Selector_2 s16062_7(wires_4015_6[2], addr_4015_6, addr_positional[64251:64248], addr_16062_7);

wire[31:0] addr_16063_7;

Selector_2 s16063_7(wires_4015_6[3], addr_4015_6, addr_positional[64255:64252], addr_16063_7);

wire[31:0] addr_16064_7;

Selector_2 s16064_7(wires_4016_6[0], addr_4016_6, addr_positional[64259:64256], addr_16064_7);

wire[31:0] addr_16065_7;

Selector_2 s16065_7(wires_4016_6[1], addr_4016_6, addr_positional[64263:64260], addr_16065_7);

wire[31:0] addr_16066_7;

Selector_2 s16066_7(wires_4016_6[2], addr_4016_6, addr_positional[64267:64264], addr_16066_7);

wire[31:0] addr_16067_7;

Selector_2 s16067_7(wires_4016_6[3], addr_4016_6, addr_positional[64271:64268], addr_16067_7);

wire[31:0] addr_16068_7;

Selector_2 s16068_7(wires_4017_6[0], addr_4017_6, addr_positional[64275:64272], addr_16068_7);

wire[31:0] addr_16069_7;

Selector_2 s16069_7(wires_4017_6[1], addr_4017_6, addr_positional[64279:64276], addr_16069_7);

wire[31:0] addr_16070_7;

Selector_2 s16070_7(wires_4017_6[2], addr_4017_6, addr_positional[64283:64280], addr_16070_7);

wire[31:0] addr_16071_7;

Selector_2 s16071_7(wires_4017_6[3], addr_4017_6, addr_positional[64287:64284], addr_16071_7);

wire[31:0] addr_16072_7;

Selector_2 s16072_7(wires_4018_6[0], addr_4018_6, addr_positional[64291:64288], addr_16072_7);

wire[31:0] addr_16073_7;

Selector_2 s16073_7(wires_4018_6[1], addr_4018_6, addr_positional[64295:64292], addr_16073_7);

wire[31:0] addr_16074_7;

Selector_2 s16074_7(wires_4018_6[2], addr_4018_6, addr_positional[64299:64296], addr_16074_7);

wire[31:0] addr_16075_7;

Selector_2 s16075_7(wires_4018_6[3], addr_4018_6, addr_positional[64303:64300], addr_16075_7);

wire[31:0] addr_16076_7;

Selector_2 s16076_7(wires_4019_6[0], addr_4019_6, addr_positional[64307:64304], addr_16076_7);

wire[31:0] addr_16077_7;

Selector_2 s16077_7(wires_4019_6[1], addr_4019_6, addr_positional[64311:64308], addr_16077_7);

wire[31:0] addr_16078_7;

Selector_2 s16078_7(wires_4019_6[2], addr_4019_6, addr_positional[64315:64312], addr_16078_7);

wire[31:0] addr_16079_7;

Selector_2 s16079_7(wires_4019_6[3], addr_4019_6, addr_positional[64319:64316], addr_16079_7);

wire[31:0] addr_16080_7;

Selector_2 s16080_7(wires_4020_6[0], addr_4020_6, addr_positional[64323:64320], addr_16080_7);

wire[31:0] addr_16081_7;

Selector_2 s16081_7(wires_4020_6[1], addr_4020_6, addr_positional[64327:64324], addr_16081_7);

wire[31:0] addr_16082_7;

Selector_2 s16082_7(wires_4020_6[2], addr_4020_6, addr_positional[64331:64328], addr_16082_7);

wire[31:0] addr_16083_7;

Selector_2 s16083_7(wires_4020_6[3], addr_4020_6, addr_positional[64335:64332], addr_16083_7);

wire[31:0] addr_16084_7;

Selector_2 s16084_7(wires_4021_6[0], addr_4021_6, addr_positional[64339:64336], addr_16084_7);

wire[31:0] addr_16085_7;

Selector_2 s16085_7(wires_4021_6[1], addr_4021_6, addr_positional[64343:64340], addr_16085_7);

wire[31:0] addr_16086_7;

Selector_2 s16086_7(wires_4021_6[2], addr_4021_6, addr_positional[64347:64344], addr_16086_7);

wire[31:0] addr_16087_7;

Selector_2 s16087_7(wires_4021_6[3], addr_4021_6, addr_positional[64351:64348], addr_16087_7);

wire[31:0] addr_16088_7;

Selector_2 s16088_7(wires_4022_6[0], addr_4022_6, addr_positional[64355:64352], addr_16088_7);

wire[31:0] addr_16089_7;

Selector_2 s16089_7(wires_4022_6[1], addr_4022_6, addr_positional[64359:64356], addr_16089_7);

wire[31:0] addr_16090_7;

Selector_2 s16090_7(wires_4022_6[2], addr_4022_6, addr_positional[64363:64360], addr_16090_7);

wire[31:0] addr_16091_7;

Selector_2 s16091_7(wires_4022_6[3], addr_4022_6, addr_positional[64367:64364], addr_16091_7);

wire[31:0] addr_16092_7;

Selector_2 s16092_7(wires_4023_6[0], addr_4023_6, addr_positional[64371:64368], addr_16092_7);

wire[31:0] addr_16093_7;

Selector_2 s16093_7(wires_4023_6[1], addr_4023_6, addr_positional[64375:64372], addr_16093_7);

wire[31:0] addr_16094_7;

Selector_2 s16094_7(wires_4023_6[2], addr_4023_6, addr_positional[64379:64376], addr_16094_7);

wire[31:0] addr_16095_7;

Selector_2 s16095_7(wires_4023_6[3], addr_4023_6, addr_positional[64383:64380], addr_16095_7);

wire[31:0] addr_16096_7;

Selector_2 s16096_7(wires_4024_6[0], addr_4024_6, addr_positional[64387:64384], addr_16096_7);

wire[31:0] addr_16097_7;

Selector_2 s16097_7(wires_4024_6[1], addr_4024_6, addr_positional[64391:64388], addr_16097_7);

wire[31:0] addr_16098_7;

Selector_2 s16098_7(wires_4024_6[2], addr_4024_6, addr_positional[64395:64392], addr_16098_7);

wire[31:0] addr_16099_7;

Selector_2 s16099_7(wires_4024_6[3], addr_4024_6, addr_positional[64399:64396], addr_16099_7);

wire[31:0] addr_16100_7;

Selector_2 s16100_7(wires_4025_6[0], addr_4025_6, addr_positional[64403:64400], addr_16100_7);

wire[31:0] addr_16101_7;

Selector_2 s16101_7(wires_4025_6[1], addr_4025_6, addr_positional[64407:64404], addr_16101_7);

wire[31:0] addr_16102_7;

Selector_2 s16102_7(wires_4025_6[2], addr_4025_6, addr_positional[64411:64408], addr_16102_7);

wire[31:0] addr_16103_7;

Selector_2 s16103_7(wires_4025_6[3], addr_4025_6, addr_positional[64415:64412], addr_16103_7);

wire[31:0] addr_16104_7;

Selector_2 s16104_7(wires_4026_6[0], addr_4026_6, addr_positional[64419:64416], addr_16104_7);

wire[31:0] addr_16105_7;

Selector_2 s16105_7(wires_4026_6[1], addr_4026_6, addr_positional[64423:64420], addr_16105_7);

wire[31:0] addr_16106_7;

Selector_2 s16106_7(wires_4026_6[2], addr_4026_6, addr_positional[64427:64424], addr_16106_7);

wire[31:0] addr_16107_7;

Selector_2 s16107_7(wires_4026_6[3], addr_4026_6, addr_positional[64431:64428], addr_16107_7);

wire[31:0] addr_16108_7;

Selector_2 s16108_7(wires_4027_6[0], addr_4027_6, addr_positional[64435:64432], addr_16108_7);

wire[31:0] addr_16109_7;

Selector_2 s16109_7(wires_4027_6[1], addr_4027_6, addr_positional[64439:64436], addr_16109_7);

wire[31:0] addr_16110_7;

Selector_2 s16110_7(wires_4027_6[2], addr_4027_6, addr_positional[64443:64440], addr_16110_7);

wire[31:0] addr_16111_7;

Selector_2 s16111_7(wires_4027_6[3], addr_4027_6, addr_positional[64447:64444], addr_16111_7);

wire[31:0] addr_16112_7;

Selector_2 s16112_7(wires_4028_6[0], addr_4028_6, addr_positional[64451:64448], addr_16112_7);

wire[31:0] addr_16113_7;

Selector_2 s16113_7(wires_4028_6[1], addr_4028_6, addr_positional[64455:64452], addr_16113_7);

wire[31:0] addr_16114_7;

Selector_2 s16114_7(wires_4028_6[2], addr_4028_6, addr_positional[64459:64456], addr_16114_7);

wire[31:0] addr_16115_7;

Selector_2 s16115_7(wires_4028_6[3], addr_4028_6, addr_positional[64463:64460], addr_16115_7);

wire[31:0] addr_16116_7;

Selector_2 s16116_7(wires_4029_6[0], addr_4029_6, addr_positional[64467:64464], addr_16116_7);

wire[31:0] addr_16117_7;

Selector_2 s16117_7(wires_4029_6[1], addr_4029_6, addr_positional[64471:64468], addr_16117_7);

wire[31:0] addr_16118_7;

Selector_2 s16118_7(wires_4029_6[2], addr_4029_6, addr_positional[64475:64472], addr_16118_7);

wire[31:0] addr_16119_7;

Selector_2 s16119_7(wires_4029_6[3], addr_4029_6, addr_positional[64479:64476], addr_16119_7);

wire[31:0] addr_16120_7;

Selector_2 s16120_7(wires_4030_6[0], addr_4030_6, addr_positional[64483:64480], addr_16120_7);

wire[31:0] addr_16121_7;

Selector_2 s16121_7(wires_4030_6[1], addr_4030_6, addr_positional[64487:64484], addr_16121_7);

wire[31:0] addr_16122_7;

Selector_2 s16122_7(wires_4030_6[2], addr_4030_6, addr_positional[64491:64488], addr_16122_7);

wire[31:0] addr_16123_7;

Selector_2 s16123_7(wires_4030_6[3], addr_4030_6, addr_positional[64495:64492], addr_16123_7);

wire[31:0] addr_16124_7;

Selector_2 s16124_7(wires_4031_6[0], addr_4031_6, addr_positional[64499:64496], addr_16124_7);

wire[31:0] addr_16125_7;

Selector_2 s16125_7(wires_4031_6[1], addr_4031_6, addr_positional[64503:64500], addr_16125_7);

wire[31:0] addr_16126_7;

Selector_2 s16126_7(wires_4031_6[2], addr_4031_6, addr_positional[64507:64504], addr_16126_7);

wire[31:0] addr_16127_7;

Selector_2 s16127_7(wires_4031_6[3], addr_4031_6, addr_positional[64511:64508], addr_16127_7);

wire[31:0] addr_16128_7;

Selector_2 s16128_7(wires_4032_6[0], addr_4032_6, addr_positional[64515:64512], addr_16128_7);

wire[31:0] addr_16129_7;

Selector_2 s16129_7(wires_4032_6[1], addr_4032_6, addr_positional[64519:64516], addr_16129_7);

wire[31:0] addr_16130_7;

Selector_2 s16130_7(wires_4032_6[2], addr_4032_6, addr_positional[64523:64520], addr_16130_7);

wire[31:0] addr_16131_7;

Selector_2 s16131_7(wires_4032_6[3], addr_4032_6, addr_positional[64527:64524], addr_16131_7);

wire[31:0] addr_16132_7;

Selector_2 s16132_7(wires_4033_6[0], addr_4033_6, addr_positional[64531:64528], addr_16132_7);

wire[31:0] addr_16133_7;

Selector_2 s16133_7(wires_4033_6[1], addr_4033_6, addr_positional[64535:64532], addr_16133_7);

wire[31:0] addr_16134_7;

Selector_2 s16134_7(wires_4033_6[2], addr_4033_6, addr_positional[64539:64536], addr_16134_7);

wire[31:0] addr_16135_7;

Selector_2 s16135_7(wires_4033_6[3], addr_4033_6, addr_positional[64543:64540], addr_16135_7);

wire[31:0] addr_16136_7;

Selector_2 s16136_7(wires_4034_6[0], addr_4034_6, addr_positional[64547:64544], addr_16136_7);

wire[31:0] addr_16137_7;

Selector_2 s16137_7(wires_4034_6[1], addr_4034_6, addr_positional[64551:64548], addr_16137_7);

wire[31:0] addr_16138_7;

Selector_2 s16138_7(wires_4034_6[2], addr_4034_6, addr_positional[64555:64552], addr_16138_7);

wire[31:0] addr_16139_7;

Selector_2 s16139_7(wires_4034_6[3], addr_4034_6, addr_positional[64559:64556], addr_16139_7);

wire[31:0] addr_16140_7;

Selector_2 s16140_7(wires_4035_6[0], addr_4035_6, addr_positional[64563:64560], addr_16140_7);

wire[31:0] addr_16141_7;

Selector_2 s16141_7(wires_4035_6[1], addr_4035_6, addr_positional[64567:64564], addr_16141_7);

wire[31:0] addr_16142_7;

Selector_2 s16142_7(wires_4035_6[2], addr_4035_6, addr_positional[64571:64568], addr_16142_7);

wire[31:0] addr_16143_7;

Selector_2 s16143_7(wires_4035_6[3], addr_4035_6, addr_positional[64575:64572], addr_16143_7);

wire[31:0] addr_16144_7;

Selector_2 s16144_7(wires_4036_6[0], addr_4036_6, addr_positional[64579:64576], addr_16144_7);

wire[31:0] addr_16145_7;

Selector_2 s16145_7(wires_4036_6[1], addr_4036_6, addr_positional[64583:64580], addr_16145_7);

wire[31:0] addr_16146_7;

Selector_2 s16146_7(wires_4036_6[2], addr_4036_6, addr_positional[64587:64584], addr_16146_7);

wire[31:0] addr_16147_7;

Selector_2 s16147_7(wires_4036_6[3], addr_4036_6, addr_positional[64591:64588], addr_16147_7);

wire[31:0] addr_16148_7;

Selector_2 s16148_7(wires_4037_6[0], addr_4037_6, addr_positional[64595:64592], addr_16148_7);

wire[31:0] addr_16149_7;

Selector_2 s16149_7(wires_4037_6[1], addr_4037_6, addr_positional[64599:64596], addr_16149_7);

wire[31:0] addr_16150_7;

Selector_2 s16150_7(wires_4037_6[2], addr_4037_6, addr_positional[64603:64600], addr_16150_7);

wire[31:0] addr_16151_7;

Selector_2 s16151_7(wires_4037_6[3], addr_4037_6, addr_positional[64607:64604], addr_16151_7);

wire[31:0] addr_16152_7;

Selector_2 s16152_7(wires_4038_6[0], addr_4038_6, addr_positional[64611:64608], addr_16152_7);

wire[31:0] addr_16153_7;

Selector_2 s16153_7(wires_4038_6[1], addr_4038_6, addr_positional[64615:64612], addr_16153_7);

wire[31:0] addr_16154_7;

Selector_2 s16154_7(wires_4038_6[2], addr_4038_6, addr_positional[64619:64616], addr_16154_7);

wire[31:0] addr_16155_7;

Selector_2 s16155_7(wires_4038_6[3], addr_4038_6, addr_positional[64623:64620], addr_16155_7);

wire[31:0] addr_16156_7;

Selector_2 s16156_7(wires_4039_6[0], addr_4039_6, addr_positional[64627:64624], addr_16156_7);

wire[31:0] addr_16157_7;

Selector_2 s16157_7(wires_4039_6[1], addr_4039_6, addr_positional[64631:64628], addr_16157_7);

wire[31:0] addr_16158_7;

Selector_2 s16158_7(wires_4039_6[2], addr_4039_6, addr_positional[64635:64632], addr_16158_7);

wire[31:0] addr_16159_7;

Selector_2 s16159_7(wires_4039_6[3], addr_4039_6, addr_positional[64639:64636], addr_16159_7);

wire[31:0] addr_16160_7;

Selector_2 s16160_7(wires_4040_6[0], addr_4040_6, addr_positional[64643:64640], addr_16160_7);

wire[31:0] addr_16161_7;

Selector_2 s16161_7(wires_4040_6[1], addr_4040_6, addr_positional[64647:64644], addr_16161_7);

wire[31:0] addr_16162_7;

Selector_2 s16162_7(wires_4040_6[2], addr_4040_6, addr_positional[64651:64648], addr_16162_7);

wire[31:0] addr_16163_7;

Selector_2 s16163_7(wires_4040_6[3], addr_4040_6, addr_positional[64655:64652], addr_16163_7);

wire[31:0] addr_16164_7;

Selector_2 s16164_7(wires_4041_6[0], addr_4041_6, addr_positional[64659:64656], addr_16164_7);

wire[31:0] addr_16165_7;

Selector_2 s16165_7(wires_4041_6[1], addr_4041_6, addr_positional[64663:64660], addr_16165_7);

wire[31:0] addr_16166_7;

Selector_2 s16166_7(wires_4041_6[2], addr_4041_6, addr_positional[64667:64664], addr_16166_7);

wire[31:0] addr_16167_7;

Selector_2 s16167_7(wires_4041_6[3], addr_4041_6, addr_positional[64671:64668], addr_16167_7);

wire[31:0] addr_16168_7;

Selector_2 s16168_7(wires_4042_6[0], addr_4042_6, addr_positional[64675:64672], addr_16168_7);

wire[31:0] addr_16169_7;

Selector_2 s16169_7(wires_4042_6[1], addr_4042_6, addr_positional[64679:64676], addr_16169_7);

wire[31:0] addr_16170_7;

Selector_2 s16170_7(wires_4042_6[2], addr_4042_6, addr_positional[64683:64680], addr_16170_7);

wire[31:0] addr_16171_7;

Selector_2 s16171_7(wires_4042_6[3], addr_4042_6, addr_positional[64687:64684], addr_16171_7);

wire[31:0] addr_16172_7;

Selector_2 s16172_7(wires_4043_6[0], addr_4043_6, addr_positional[64691:64688], addr_16172_7);

wire[31:0] addr_16173_7;

Selector_2 s16173_7(wires_4043_6[1], addr_4043_6, addr_positional[64695:64692], addr_16173_7);

wire[31:0] addr_16174_7;

Selector_2 s16174_7(wires_4043_6[2], addr_4043_6, addr_positional[64699:64696], addr_16174_7);

wire[31:0] addr_16175_7;

Selector_2 s16175_7(wires_4043_6[3], addr_4043_6, addr_positional[64703:64700], addr_16175_7);

wire[31:0] addr_16176_7;

Selector_2 s16176_7(wires_4044_6[0], addr_4044_6, addr_positional[64707:64704], addr_16176_7);

wire[31:0] addr_16177_7;

Selector_2 s16177_7(wires_4044_6[1], addr_4044_6, addr_positional[64711:64708], addr_16177_7);

wire[31:0] addr_16178_7;

Selector_2 s16178_7(wires_4044_6[2], addr_4044_6, addr_positional[64715:64712], addr_16178_7);

wire[31:0] addr_16179_7;

Selector_2 s16179_7(wires_4044_6[3], addr_4044_6, addr_positional[64719:64716], addr_16179_7);

wire[31:0] addr_16180_7;

Selector_2 s16180_7(wires_4045_6[0], addr_4045_6, addr_positional[64723:64720], addr_16180_7);

wire[31:0] addr_16181_7;

Selector_2 s16181_7(wires_4045_6[1], addr_4045_6, addr_positional[64727:64724], addr_16181_7);

wire[31:0] addr_16182_7;

Selector_2 s16182_7(wires_4045_6[2], addr_4045_6, addr_positional[64731:64728], addr_16182_7);

wire[31:0] addr_16183_7;

Selector_2 s16183_7(wires_4045_6[3], addr_4045_6, addr_positional[64735:64732], addr_16183_7);

wire[31:0] addr_16184_7;

Selector_2 s16184_7(wires_4046_6[0], addr_4046_6, addr_positional[64739:64736], addr_16184_7);

wire[31:0] addr_16185_7;

Selector_2 s16185_7(wires_4046_6[1], addr_4046_6, addr_positional[64743:64740], addr_16185_7);

wire[31:0] addr_16186_7;

Selector_2 s16186_7(wires_4046_6[2], addr_4046_6, addr_positional[64747:64744], addr_16186_7);

wire[31:0] addr_16187_7;

Selector_2 s16187_7(wires_4046_6[3], addr_4046_6, addr_positional[64751:64748], addr_16187_7);

wire[31:0] addr_16188_7;

Selector_2 s16188_7(wires_4047_6[0], addr_4047_6, addr_positional[64755:64752], addr_16188_7);

wire[31:0] addr_16189_7;

Selector_2 s16189_7(wires_4047_6[1], addr_4047_6, addr_positional[64759:64756], addr_16189_7);

wire[31:0] addr_16190_7;

Selector_2 s16190_7(wires_4047_6[2], addr_4047_6, addr_positional[64763:64760], addr_16190_7);

wire[31:0] addr_16191_7;

Selector_2 s16191_7(wires_4047_6[3], addr_4047_6, addr_positional[64767:64764], addr_16191_7);

wire[31:0] addr_16192_7;

Selector_2 s16192_7(wires_4048_6[0], addr_4048_6, addr_positional[64771:64768], addr_16192_7);

wire[31:0] addr_16193_7;

Selector_2 s16193_7(wires_4048_6[1], addr_4048_6, addr_positional[64775:64772], addr_16193_7);

wire[31:0] addr_16194_7;

Selector_2 s16194_7(wires_4048_6[2], addr_4048_6, addr_positional[64779:64776], addr_16194_7);

wire[31:0] addr_16195_7;

Selector_2 s16195_7(wires_4048_6[3], addr_4048_6, addr_positional[64783:64780], addr_16195_7);

wire[31:0] addr_16196_7;

Selector_2 s16196_7(wires_4049_6[0], addr_4049_6, addr_positional[64787:64784], addr_16196_7);

wire[31:0] addr_16197_7;

Selector_2 s16197_7(wires_4049_6[1], addr_4049_6, addr_positional[64791:64788], addr_16197_7);

wire[31:0] addr_16198_7;

Selector_2 s16198_7(wires_4049_6[2], addr_4049_6, addr_positional[64795:64792], addr_16198_7);

wire[31:0] addr_16199_7;

Selector_2 s16199_7(wires_4049_6[3], addr_4049_6, addr_positional[64799:64796], addr_16199_7);

wire[31:0] addr_16200_7;

Selector_2 s16200_7(wires_4050_6[0], addr_4050_6, addr_positional[64803:64800], addr_16200_7);

wire[31:0] addr_16201_7;

Selector_2 s16201_7(wires_4050_6[1], addr_4050_6, addr_positional[64807:64804], addr_16201_7);

wire[31:0] addr_16202_7;

Selector_2 s16202_7(wires_4050_6[2], addr_4050_6, addr_positional[64811:64808], addr_16202_7);

wire[31:0] addr_16203_7;

Selector_2 s16203_7(wires_4050_6[3], addr_4050_6, addr_positional[64815:64812], addr_16203_7);

wire[31:0] addr_16204_7;

Selector_2 s16204_7(wires_4051_6[0], addr_4051_6, addr_positional[64819:64816], addr_16204_7);

wire[31:0] addr_16205_7;

Selector_2 s16205_7(wires_4051_6[1], addr_4051_6, addr_positional[64823:64820], addr_16205_7);

wire[31:0] addr_16206_7;

Selector_2 s16206_7(wires_4051_6[2], addr_4051_6, addr_positional[64827:64824], addr_16206_7);

wire[31:0] addr_16207_7;

Selector_2 s16207_7(wires_4051_6[3], addr_4051_6, addr_positional[64831:64828], addr_16207_7);

wire[31:0] addr_16208_7;

Selector_2 s16208_7(wires_4052_6[0], addr_4052_6, addr_positional[64835:64832], addr_16208_7);

wire[31:0] addr_16209_7;

Selector_2 s16209_7(wires_4052_6[1], addr_4052_6, addr_positional[64839:64836], addr_16209_7);

wire[31:0] addr_16210_7;

Selector_2 s16210_7(wires_4052_6[2], addr_4052_6, addr_positional[64843:64840], addr_16210_7);

wire[31:0] addr_16211_7;

Selector_2 s16211_7(wires_4052_6[3], addr_4052_6, addr_positional[64847:64844], addr_16211_7);

wire[31:0] addr_16212_7;

Selector_2 s16212_7(wires_4053_6[0], addr_4053_6, addr_positional[64851:64848], addr_16212_7);

wire[31:0] addr_16213_7;

Selector_2 s16213_7(wires_4053_6[1], addr_4053_6, addr_positional[64855:64852], addr_16213_7);

wire[31:0] addr_16214_7;

Selector_2 s16214_7(wires_4053_6[2], addr_4053_6, addr_positional[64859:64856], addr_16214_7);

wire[31:0] addr_16215_7;

Selector_2 s16215_7(wires_4053_6[3], addr_4053_6, addr_positional[64863:64860], addr_16215_7);

wire[31:0] addr_16216_7;

Selector_2 s16216_7(wires_4054_6[0], addr_4054_6, addr_positional[64867:64864], addr_16216_7);

wire[31:0] addr_16217_7;

Selector_2 s16217_7(wires_4054_6[1], addr_4054_6, addr_positional[64871:64868], addr_16217_7);

wire[31:0] addr_16218_7;

Selector_2 s16218_7(wires_4054_6[2], addr_4054_6, addr_positional[64875:64872], addr_16218_7);

wire[31:0] addr_16219_7;

Selector_2 s16219_7(wires_4054_6[3], addr_4054_6, addr_positional[64879:64876], addr_16219_7);

wire[31:0] addr_16220_7;

Selector_2 s16220_7(wires_4055_6[0], addr_4055_6, addr_positional[64883:64880], addr_16220_7);

wire[31:0] addr_16221_7;

Selector_2 s16221_7(wires_4055_6[1], addr_4055_6, addr_positional[64887:64884], addr_16221_7);

wire[31:0] addr_16222_7;

Selector_2 s16222_7(wires_4055_6[2], addr_4055_6, addr_positional[64891:64888], addr_16222_7);

wire[31:0] addr_16223_7;

Selector_2 s16223_7(wires_4055_6[3], addr_4055_6, addr_positional[64895:64892], addr_16223_7);

wire[31:0] addr_16224_7;

Selector_2 s16224_7(wires_4056_6[0], addr_4056_6, addr_positional[64899:64896], addr_16224_7);

wire[31:0] addr_16225_7;

Selector_2 s16225_7(wires_4056_6[1], addr_4056_6, addr_positional[64903:64900], addr_16225_7);

wire[31:0] addr_16226_7;

Selector_2 s16226_7(wires_4056_6[2], addr_4056_6, addr_positional[64907:64904], addr_16226_7);

wire[31:0] addr_16227_7;

Selector_2 s16227_7(wires_4056_6[3], addr_4056_6, addr_positional[64911:64908], addr_16227_7);

wire[31:0] addr_16228_7;

Selector_2 s16228_7(wires_4057_6[0], addr_4057_6, addr_positional[64915:64912], addr_16228_7);

wire[31:0] addr_16229_7;

Selector_2 s16229_7(wires_4057_6[1], addr_4057_6, addr_positional[64919:64916], addr_16229_7);

wire[31:0] addr_16230_7;

Selector_2 s16230_7(wires_4057_6[2], addr_4057_6, addr_positional[64923:64920], addr_16230_7);

wire[31:0] addr_16231_7;

Selector_2 s16231_7(wires_4057_6[3], addr_4057_6, addr_positional[64927:64924], addr_16231_7);

wire[31:0] addr_16232_7;

Selector_2 s16232_7(wires_4058_6[0], addr_4058_6, addr_positional[64931:64928], addr_16232_7);

wire[31:0] addr_16233_7;

Selector_2 s16233_7(wires_4058_6[1], addr_4058_6, addr_positional[64935:64932], addr_16233_7);

wire[31:0] addr_16234_7;

Selector_2 s16234_7(wires_4058_6[2], addr_4058_6, addr_positional[64939:64936], addr_16234_7);

wire[31:0] addr_16235_7;

Selector_2 s16235_7(wires_4058_6[3], addr_4058_6, addr_positional[64943:64940], addr_16235_7);

wire[31:0] addr_16236_7;

Selector_2 s16236_7(wires_4059_6[0], addr_4059_6, addr_positional[64947:64944], addr_16236_7);

wire[31:0] addr_16237_7;

Selector_2 s16237_7(wires_4059_6[1], addr_4059_6, addr_positional[64951:64948], addr_16237_7);

wire[31:0] addr_16238_7;

Selector_2 s16238_7(wires_4059_6[2], addr_4059_6, addr_positional[64955:64952], addr_16238_7);

wire[31:0] addr_16239_7;

Selector_2 s16239_7(wires_4059_6[3], addr_4059_6, addr_positional[64959:64956], addr_16239_7);

wire[31:0] addr_16240_7;

Selector_2 s16240_7(wires_4060_6[0], addr_4060_6, addr_positional[64963:64960], addr_16240_7);

wire[31:0] addr_16241_7;

Selector_2 s16241_7(wires_4060_6[1], addr_4060_6, addr_positional[64967:64964], addr_16241_7);

wire[31:0] addr_16242_7;

Selector_2 s16242_7(wires_4060_6[2], addr_4060_6, addr_positional[64971:64968], addr_16242_7);

wire[31:0] addr_16243_7;

Selector_2 s16243_7(wires_4060_6[3], addr_4060_6, addr_positional[64975:64972], addr_16243_7);

wire[31:0] addr_16244_7;

Selector_2 s16244_7(wires_4061_6[0], addr_4061_6, addr_positional[64979:64976], addr_16244_7);

wire[31:0] addr_16245_7;

Selector_2 s16245_7(wires_4061_6[1], addr_4061_6, addr_positional[64983:64980], addr_16245_7);

wire[31:0] addr_16246_7;

Selector_2 s16246_7(wires_4061_6[2], addr_4061_6, addr_positional[64987:64984], addr_16246_7);

wire[31:0] addr_16247_7;

Selector_2 s16247_7(wires_4061_6[3], addr_4061_6, addr_positional[64991:64988], addr_16247_7);

wire[31:0] addr_16248_7;

Selector_2 s16248_7(wires_4062_6[0], addr_4062_6, addr_positional[64995:64992], addr_16248_7);

wire[31:0] addr_16249_7;

Selector_2 s16249_7(wires_4062_6[1], addr_4062_6, addr_positional[64999:64996], addr_16249_7);

wire[31:0] addr_16250_7;

Selector_2 s16250_7(wires_4062_6[2], addr_4062_6, addr_positional[65003:65000], addr_16250_7);

wire[31:0] addr_16251_7;

Selector_2 s16251_7(wires_4062_6[3], addr_4062_6, addr_positional[65007:65004], addr_16251_7);

wire[31:0] addr_16252_7;

Selector_2 s16252_7(wires_4063_6[0], addr_4063_6, addr_positional[65011:65008], addr_16252_7);

wire[31:0] addr_16253_7;

Selector_2 s16253_7(wires_4063_6[1], addr_4063_6, addr_positional[65015:65012], addr_16253_7);

wire[31:0] addr_16254_7;

Selector_2 s16254_7(wires_4063_6[2], addr_4063_6, addr_positional[65019:65016], addr_16254_7);

wire[31:0] addr_16255_7;

Selector_2 s16255_7(wires_4063_6[3], addr_4063_6, addr_positional[65023:65020], addr_16255_7);

wire[31:0] addr_16256_7;

Selector_2 s16256_7(wires_4064_6[0], addr_4064_6, addr_positional[65027:65024], addr_16256_7);

wire[31:0] addr_16257_7;

Selector_2 s16257_7(wires_4064_6[1], addr_4064_6, addr_positional[65031:65028], addr_16257_7);

wire[31:0] addr_16258_7;

Selector_2 s16258_7(wires_4064_6[2], addr_4064_6, addr_positional[65035:65032], addr_16258_7);

wire[31:0] addr_16259_7;

Selector_2 s16259_7(wires_4064_6[3], addr_4064_6, addr_positional[65039:65036], addr_16259_7);

wire[31:0] addr_16260_7;

Selector_2 s16260_7(wires_4065_6[0], addr_4065_6, addr_positional[65043:65040], addr_16260_7);

wire[31:0] addr_16261_7;

Selector_2 s16261_7(wires_4065_6[1], addr_4065_6, addr_positional[65047:65044], addr_16261_7);

wire[31:0] addr_16262_7;

Selector_2 s16262_7(wires_4065_6[2], addr_4065_6, addr_positional[65051:65048], addr_16262_7);

wire[31:0] addr_16263_7;

Selector_2 s16263_7(wires_4065_6[3], addr_4065_6, addr_positional[65055:65052], addr_16263_7);

wire[31:0] addr_16264_7;

Selector_2 s16264_7(wires_4066_6[0], addr_4066_6, addr_positional[65059:65056], addr_16264_7);

wire[31:0] addr_16265_7;

Selector_2 s16265_7(wires_4066_6[1], addr_4066_6, addr_positional[65063:65060], addr_16265_7);

wire[31:0] addr_16266_7;

Selector_2 s16266_7(wires_4066_6[2], addr_4066_6, addr_positional[65067:65064], addr_16266_7);

wire[31:0] addr_16267_7;

Selector_2 s16267_7(wires_4066_6[3], addr_4066_6, addr_positional[65071:65068], addr_16267_7);

wire[31:0] addr_16268_7;

Selector_2 s16268_7(wires_4067_6[0], addr_4067_6, addr_positional[65075:65072], addr_16268_7);

wire[31:0] addr_16269_7;

Selector_2 s16269_7(wires_4067_6[1], addr_4067_6, addr_positional[65079:65076], addr_16269_7);

wire[31:0] addr_16270_7;

Selector_2 s16270_7(wires_4067_6[2], addr_4067_6, addr_positional[65083:65080], addr_16270_7);

wire[31:0] addr_16271_7;

Selector_2 s16271_7(wires_4067_6[3], addr_4067_6, addr_positional[65087:65084], addr_16271_7);

wire[31:0] addr_16272_7;

Selector_2 s16272_7(wires_4068_6[0], addr_4068_6, addr_positional[65091:65088], addr_16272_7);

wire[31:0] addr_16273_7;

Selector_2 s16273_7(wires_4068_6[1], addr_4068_6, addr_positional[65095:65092], addr_16273_7);

wire[31:0] addr_16274_7;

Selector_2 s16274_7(wires_4068_6[2], addr_4068_6, addr_positional[65099:65096], addr_16274_7);

wire[31:0] addr_16275_7;

Selector_2 s16275_7(wires_4068_6[3], addr_4068_6, addr_positional[65103:65100], addr_16275_7);

wire[31:0] addr_16276_7;

Selector_2 s16276_7(wires_4069_6[0], addr_4069_6, addr_positional[65107:65104], addr_16276_7);

wire[31:0] addr_16277_7;

Selector_2 s16277_7(wires_4069_6[1], addr_4069_6, addr_positional[65111:65108], addr_16277_7);

wire[31:0] addr_16278_7;

Selector_2 s16278_7(wires_4069_6[2], addr_4069_6, addr_positional[65115:65112], addr_16278_7);

wire[31:0] addr_16279_7;

Selector_2 s16279_7(wires_4069_6[3], addr_4069_6, addr_positional[65119:65116], addr_16279_7);

wire[31:0] addr_16280_7;

Selector_2 s16280_7(wires_4070_6[0], addr_4070_6, addr_positional[65123:65120], addr_16280_7);

wire[31:0] addr_16281_7;

Selector_2 s16281_7(wires_4070_6[1], addr_4070_6, addr_positional[65127:65124], addr_16281_7);

wire[31:0] addr_16282_7;

Selector_2 s16282_7(wires_4070_6[2], addr_4070_6, addr_positional[65131:65128], addr_16282_7);

wire[31:0] addr_16283_7;

Selector_2 s16283_7(wires_4070_6[3], addr_4070_6, addr_positional[65135:65132], addr_16283_7);

wire[31:0] addr_16284_7;

Selector_2 s16284_7(wires_4071_6[0], addr_4071_6, addr_positional[65139:65136], addr_16284_7);

wire[31:0] addr_16285_7;

Selector_2 s16285_7(wires_4071_6[1], addr_4071_6, addr_positional[65143:65140], addr_16285_7);

wire[31:0] addr_16286_7;

Selector_2 s16286_7(wires_4071_6[2], addr_4071_6, addr_positional[65147:65144], addr_16286_7);

wire[31:0] addr_16287_7;

Selector_2 s16287_7(wires_4071_6[3], addr_4071_6, addr_positional[65151:65148], addr_16287_7);

wire[31:0] addr_16288_7;

Selector_2 s16288_7(wires_4072_6[0], addr_4072_6, addr_positional[65155:65152], addr_16288_7);

wire[31:0] addr_16289_7;

Selector_2 s16289_7(wires_4072_6[1], addr_4072_6, addr_positional[65159:65156], addr_16289_7);

wire[31:0] addr_16290_7;

Selector_2 s16290_7(wires_4072_6[2], addr_4072_6, addr_positional[65163:65160], addr_16290_7);

wire[31:0] addr_16291_7;

Selector_2 s16291_7(wires_4072_6[3], addr_4072_6, addr_positional[65167:65164], addr_16291_7);

wire[31:0] addr_16292_7;

Selector_2 s16292_7(wires_4073_6[0], addr_4073_6, addr_positional[65171:65168], addr_16292_7);

wire[31:0] addr_16293_7;

Selector_2 s16293_7(wires_4073_6[1], addr_4073_6, addr_positional[65175:65172], addr_16293_7);

wire[31:0] addr_16294_7;

Selector_2 s16294_7(wires_4073_6[2], addr_4073_6, addr_positional[65179:65176], addr_16294_7);

wire[31:0] addr_16295_7;

Selector_2 s16295_7(wires_4073_6[3], addr_4073_6, addr_positional[65183:65180], addr_16295_7);

wire[31:0] addr_16296_7;

Selector_2 s16296_7(wires_4074_6[0], addr_4074_6, addr_positional[65187:65184], addr_16296_7);

wire[31:0] addr_16297_7;

Selector_2 s16297_7(wires_4074_6[1], addr_4074_6, addr_positional[65191:65188], addr_16297_7);

wire[31:0] addr_16298_7;

Selector_2 s16298_7(wires_4074_6[2], addr_4074_6, addr_positional[65195:65192], addr_16298_7);

wire[31:0] addr_16299_7;

Selector_2 s16299_7(wires_4074_6[3], addr_4074_6, addr_positional[65199:65196], addr_16299_7);

wire[31:0] addr_16300_7;

Selector_2 s16300_7(wires_4075_6[0], addr_4075_6, addr_positional[65203:65200], addr_16300_7);

wire[31:0] addr_16301_7;

Selector_2 s16301_7(wires_4075_6[1], addr_4075_6, addr_positional[65207:65204], addr_16301_7);

wire[31:0] addr_16302_7;

Selector_2 s16302_7(wires_4075_6[2], addr_4075_6, addr_positional[65211:65208], addr_16302_7);

wire[31:0] addr_16303_7;

Selector_2 s16303_7(wires_4075_6[3], addr_4075_6, addr_positional[65215:65212], addr_16303_7);

wire[31:0] addr_16304_7;

Selector_2 s16304_7(wires_4076_6[0], addr_4076_6, addr_positional[65219:65216], addr_16304_7);

wire[31:0] addr_16305_7;

Selector_2 s16305_7(wires_4076_6[1], addr_4076_6, addr_positional[65223:65220], addr_16305_7);

wire[31:0] addr_16306_7;

Selector_2 s16306_7(wires_4076_6[2], addr_4076_6, addr_positional[65227:65224], addr_16306_7);

wire[31:0] addr_16307_7;

Selector_2 s16307_7(wires_4076_6[3], addr_4076_6, addr_positional[65231:65228], addr_16307_7);

wire[31:0] addr_16308_7;

Selector_2 s16308_7(wires_4077_6[0], addr_4077_6, addr_positional[65235:65232], addr_16308_7);

wire[31:0] addr_16309_7;

Selector_2 s16309_7(wires_4077_6[1], addr_4077_6, addr_positional[65239:65236], addr_16309_7);

wire[31:0] addr_16310_7;

Selector_2 s16310_7(wires_4077_6[2], addr_4077_6, addr_positional[65243:65240], addr_16310_7);

wire[31:0] addr_16311_7;

Selector_2 s16311_7(wires_4077_6[3], addr_4077_6, addr_positional[65247:65244], addr_16311_7);

wire[31:0] addr_16312_7;

Selector_2 s16312_7(wires_4078_6[0], addr_4078_6, addr_positional[65251:65248], addr_16312_7);

wire[31:0] addr_16313_7;

Selector_2 s16313_7(wires_4078_6[1], addr_4078_6, addr_positional[65255:65252], addr_16313_7);

wire[31:0] addr_16314_7;

Selector_2 s16314_7(wires_4078_6[2], addr_4078_6, addr_positional[65259:65256], addr_16314_7);

wire[31:0] addr_16315_7;

Selector_2 s16315_7(wires_4078_6[3], addr_4078_6, addr_positional[65263:65260], addr_16315_7);

wire[31:0] addr_16316_7;

Selector_2 s16316_7(wires_4079_6[0], addr_4079_6, addr_positional[65267:65264], addr_16316_7);

wire[31:0] addr_16317_7;

Selector_2 s16317_7(wires_4079_6[1], addr_4079_6, addr_positional[65271:65268], addr_16317_7);

wire[31:0] addr_16318_7;

Selector_2 s16318_7(wires_4079_6[2], addr_4079_6, addr_positional[65275:65272], addr_16318_7);

wire[31:0] addr_16319_7;

Selector_2 s16319_7(wires_4079_6[3], addr_4079_6, addr_positional[65279:65276], addr_16319_7);

wire[31:0] addr_16320_7;

Selector_2 s16320_7(wires_4080_6[0], addr_4080_6, addr_positional[65283:65280], addr_16320_7);

wire[31:0] addr_16321_7;

Selector_2 s16321_7(wires_4080_6[1], addr_4080_6, addr_positional[65287:65284], addr_16321_7);

wire[31:0] addr_16322_7;

Selector_2 s16322_7(wires_4080_6[2], addr_4080_6, addr_positional[65291:65288], addr_16322_7);

wire[31:0] addr_16323_7;

Selector_2 s16323_7(wires_4080_6[3], addr_4080_6, addr_positional[65295:65292], addr_16323_7);

wire[31:0] addr_16324_7;

Selector_2 s16324_7(wires_4081_6[0], addr_4081_6, addr_positional[65299:65296], addr_16324_7);

wire[31:0] addr_16325_7;

Selector_2 s16325_7(wires_4081_6[1], addr_4081_6, addr_positional[65303:65300], addr_16325_7);

wire[31:0] addr_16326_7;

Selector_2 s16326_7(wires_4081_6[2], addr_4081_6, addr_positional[65307:65304], addr_16326_7);

wire[31:0] addr_16327_7;

Selector_2 s16327_7(wires_4081_6[3], addr_4081_6, addr_positional[65311:65308], addr_16327_7);

wire[31:0] addr_16328_7;

Selector_2 s16328_7(wires_4082_6[0], addr_4082_6, addr_positional[65315:65312], addr_16328_7);

wire[31:0] addr_16329_7;

Selector_2 s16329_7(wires_4082_6[1], addr_4082_6, addr_positional[65319:65316], addr_16329_7);

wire[31:0] addr_16330_7;

Selector_2 s16330_7(wires_4082_6[2], addr_4082_6, addr_positional[65323:65320], addr_16330_7);

wire[31:0] addr_16331_7;

Selector_2 s16331_7(wires_4082_6[3], addr_4082_6, addr_positional[65327:65324], addr_16331_7);

wire[31:0] addr_16332_7;

Selector_2 s16332_7(wires_4083_6[0], addr_4083_6, addr_positional[65331:65328], addr_16332_7);

wire[31:0] addr_16333_7;

Selector_2 s16333_7(wires_4083_6[1], addr_4083_6, addr_positional[65335:65332], addr_16333_7);

wire[31:0] addr_16334_7;

Selector_2 s16334_7(wires_4083_6[2], addr_4083_6, addr_positional[65339:65336], addr_16334_7);

wire[31:0] addr_16335_7;

Selector_2 s16335_7(wires_4083_6[3], addr_4083_6, addr_positional[65343:65340], addr_16335_7);

wire[31:0] addr_16336_7;

Selector_2 s16336_7(wires_4084_6[0], addr_4084_6, addr_positional[65347:65344], addr_16336_7);

wire[31:0] addr_16337_7;

Selector_2 s16337_7(wires_4084_6[1], addr_4084_6, addr_positional[65351:65348], addr_16337_7);

wire[31:0] addr_16338_7;

Selector_2 s16338_7(wires_4084_6[2], addr_4084_6, addr_positional[65355:65352], addr_16338_7);

wire[31:0] addr_16339_7;

Selector_2 s16339_7(wires_4084_6[3], addr_4084_6, addr_positional[65359:65356], addr_16339_7);

wire[31:0] addr_16340_7;

Selector_2 s16340_7(wires_4085_6[0], addr_4085_6, addr_positional[65363:65360], addr_16340_7);

wire[31:0] addr_16341_7;

Selector_2 s16341_7(wires_4085_6[1], addr_4085_6, addr_positional[65367:65364], addr_16341_7);

wire[31:0] addr_16342_7;

Selector_2 s16342_7(wires_4085_6[2], addr_4085_6, addr_positional[65371:65368], addr_16342_7);

wire[31:0] addr_16343_7;

Selector_2 s16343_7(wires_4085_6[3], addr_4085_6, addr_positional[65375:65372], addr_16343_7);

wire[31:0] addr_16344_7;

Selector_2 s16344_7(wires_4086_6[0], addr_4086_6, addr_positional[65379:65376], addr_16344_7);

wire[31:0] addr_16345_7;

Selector_2 s16345_7(wires_4086_6[1], addr_4086_6, addr_positional[65383:65380], addr_16345_7);

wire[31:0] addr_16346_7;

Selector_2 s16346_7(wires_4086_6[2], addr_4086_6, addr_positional[65387:65384], addr_16346_7);

wire[31:0] addr_16347_7;

Selector_2 s16347_7(wires_4086_6[3], addr_4086_6, addr_positional[65391:65388], addr_16347_7);

wire[31:0] addr_16348_7;

Selector_2 s16348_7(wires_4087_6[0], addr_4087_6, addr_positional[65395:65392], addr_16348_7);

wire[31:0] addr_16349_7;

Selector_2 s16349_7(wires_4087_6[1], addr_4087_6, addr_positional[65399:65396], addr_16349_7);

wire[31:0] addr_16350_7;

Selector_2 s16350_7(wires_4087_6[2], addr_4087_6, addr_positional[65403:65400], addr_16350_7);

wire[31:0] addr_16351_7;

Selector_2 s16351_7(wires_4087_6[3], addr_4087_6, addr_positional[65407:65404], addr_16351_7);

wire[31:0] addr_16352_7;

Selector_2 s16352_7(wires_4088_6[0], addr_4088_6, addr_positional[65411:65408], addr_16352_7);

wire[31:0] addr_16353_7;

Selector_2 s16353_7(wires_4088_6[1], addr_4088_6, addr_positional[65415:65412], addr_16353_7);

wire[31:0] addr_16354_7;

Selector_2 s16354_7(wires_4088_6[2], addr_4088_6, addr_positional[65419:65416], addr_16354_7);

wire[31:0] addr_16355_7;

Selector_2 s16355_7(wires_4088_6[3], addr_4088_6, addr_positional[65423:65420], addr_16355_7);

wire[31:0] addr_16356_7;

Selector_2 s16356_7(wires_4089_6[0], addr_4089_6, addr_positional[65427:65424], addr_16356_7);

wire[31:0] addr_16357_7;

Selector_2 s16357_7(wires_4089_6[1], addr_4089_6, addr_positional[65431:65428], addr_16357_7);

wire[31:0] addr_16358_7;

Selector_2 s16358_7(wires_4089_6[2], addr_4089_6, addr_positional[65435:65432], addr_16358_7);

wire[31:0] addr_16359_7;

Selector_2 s16359_7(wires_4089_6[3], addr_4089_6, addr_positional[65439:65436], addr_16359_7);

wire[31:0] addr_16360_7;

Selector_2 s16360_7(wires_4090_6[0], addr_4090_6, addr_positional[65443:65440], addr_16360_7);

wire[31:0] addr_16361_7;

Selector_2 s16361_7(wires_4090_6[1], addr_4090_6, addr_positional[65447:65444], addr_16361_7);

wire[31:0] addr_16362_7;

Selector_2 s16362_7(wires_4090_6[2], addr_4090_6, addr_positional[65451:65448], addr_16362_7);

wire[31:0] addr_16363_7;

Selector_2 s16363_7(wires_4090_6[3], addr_4090_6, addr_positional[65455:65452], addr_16363_7);

wire[31:0] addr_16364_7;

Selector_2 s16364_7(wires_4091_6[0], addr_4091_6, addr_positional[65459:65456], addr_16364_7);

wire[31:0] addr_16365_7;

Selector_2 s16365_7(wires_4091_6[1], addr_4091_6, addr_positional[65463:65460], addr_16365_7);

wire[31:0] addr_16366_7;

Selector_2 s16366_7(wires_4091_6[2], addr_4091_6, addr_positional[65467:65464], addr_16366_7);

wire[31:0] addr_16367_7;

Selector_2 s16367_7(wires_4091_6[3], addr_4091_6, addr_positional[65471:65468], addr_16367_7);

wire[31:0] addr_16368_7;

Selector_2 s16368_7(wires_4092_6[0], addr_4092_6, addr_positional[65475:65472], addr_16368_7);

wire[31:0] addr_16369_7;

Selector_2 s16369_7(wires_4092_6[1], addr_4092_6, addr_positional[65479:65476], addr_16369_7);

wire[31:0] addr_16370_7;

Selector_2 s16370_7(wires_4092_6[2], addr_4092_6, addr_positional[65483:65480], addr_16370_7);

wire[31:0] addr_16371_7;

Selector_2 s16371_7(wires_4092_6[3], addr_4092_6, addr_positional[65487:65484], addr_16371_7);

wire[31:0] addr_16372_7;

Selector_2 s16372_7(wires_4093_6[0], addr_4093_6, addr_positional[65491:65488], addr_16372_7);

wire[31:0] addr_16373_7;

Selector_2 s16373_7(wires_4093_6[1], addr_4093_6, addr_positional[65495:65492], addr_16373_7);

wire[31:0] addr_16374_7;

Selector_2 s16374_7(wires_4093_6[2], addr_4093_6, addr_positional[65499:65496], addr_16374_7);

wire[31:0] addr_16375_7;

Selector_2 s16375_7(wires_4093_6[3], addr_4093_6, addr_positional[65503:65500], addr_16375_7);

wire[31:0] addr_16376_7;

Selector_2 s16376_7(wires_4094_6[0], addr_4094_6, addr_positional[65507:65504], addr_16376_7);

wire[31:0] addr_16377_7;

Selector_2 s16377_7(wires_4094_6[1], addr_4094_6, addr_positional[65511:65508], addr_16377_7);

wire[31:0] addr_16378_7;

Selector_2 s16378_7(wires_4094_6[2], addr_4094_6, addr_positional[65515:65512], addr_16378_7);

wire[31:0] addr_16379_7;

Selector_2 s16379_7(wires_4094_6[3], addr_4094_6, addr_positional[65519:65516], addr_16379_7);

wire[31:0] addr_16380_7;

Selector_2 s16380_7(wires_4095_6[0], addr_4095_6, addr_positional[65523:65520], addr_16380_7);

wire[31:0] addr_16381_7;

Selector_2 s16381_7(wires_4095_6[1], addr_4095_6, addr_positional[65527:65524], addr_16381_7);

wire[31:0] addr_16382_7;

Selector_2 s16382_7(wires_4095_6[2], addr_4095_6, addr_positional[65531:65528], addr_16382_7);

wire[31:0] addr_16383_7;

Selector_2 s16383_7(wires_4095_6[3], addr_4095_6, addr_positional[65535:65532], addr_16383_7);



endmodule

